.include "/home/taf27/hspice/libs/CMOS_180nm_L49.lib"
.include "sram_cell.sp"

Vdd vdd gnd dc 1.8
Vword word gnd pulse 0 1.8 20n 1n 1n 100n 200n

.param W1 = 11
.param W5 = 18

X1 q qb bit bitb word vdd gnd SRAM_Cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2
Cb bit gnd 2p
Cbb bitb gnd 2p

.ic q=0 qb=1.8 bit=1.8 bitb = 1.8
.options post probe 

.tran 0.5p 120n uic sweep data=myData
.probe tran V(bit) V(bitb) V(word) V(q) V(qb)
.measure tran q_max MAX V(q) FROM 0n TO 120n
.measure tran bitline_min MIN V(bit) FROM 0n TO 120n

.data myData W1 W5
2 2
2 3
3 2
2 4
3 3
4 2
2 5
3 4
4 3
5 2
2 6
3 5
4 4
5 3
6 2
2 7
3 6
4 5
5 4
6 3
7 2
2 8
3 7
4 6
5 5
6 4
7 3
8 2
2 9
3 8
4 7
5 6
6 5
7 4
8 3
9 2
2 10
3 9
4 8
5 7
6 6
7 5
8 4
9 3
10 2
2 11
3 10
4 9
5 8
6 7
7 6
8 5
9 4
10 3
11 2
2 12
3 11
4 10
5 9
6 8
7 7
8 6
9 5
10 4
11 3
12 2
2 13
3 12
4 11
5 10
6 9
7 8
8 7
9 6
10 5
11 4
12 3
13 2
2 14
3 13
4 12
5 11
6 10
7 9
8 8
9 7
10 6
11 5
12 4
13 3
14 2
2 15
3 14
4 13
5 12
6 11
7 10
8 9
9 8
10 7
11 6
12 5
13 4
14 3
15 2
2 16
3 15
4 14
5 13
6 12
7 11
8 10
9 9
10 8
11 7
12 6
13 5
14 4
15 3
16 2
2 17
3 16
4 15
5 14
6 13
7 12
8 11
9 10
10 9
11 8
12 7
13 6
14 5
15 4
16 3
17 2
2 18
3 17
4 16
5 15
6 14
7 13
8 12
9 11
10 10
11 9
12 8
13 7
14 6
15 5
16 4
17 3
18 2
2 19
3 18
4 17
5 16
6 15
7 14
8 13
9 12
10 11
11 10
12 9
13 8
14 7
15 6
16 5
17 4
18 3
19 2
2 20
3 19
4 18
5 17
6 16
7 15
8 14
9 13
10 12
11 11
12 10
13 9
14 8
15 7
16 6
17 5
18 4
19 3
20 2
3 20
4 19
5 18
6 17
7 16
8 15
9 14
10 13
11 12
12 11
13 10
14 9
15 8
16 7
17 6
18 5
19 4
20 3
4 20
5 19
6 18
7 17
8 16
9 15
10 14
11 13
12 12
13 11
14 10
15 9
16 8
17 7
18 6
19 5
20 4
5 20
6 19
7 18
8 17
9 16
10 15
11 14
12 13
13 12
14 11
15 10
16 9
17 8
18 7
19 6
20 5
6 20
7 19
8 18
9 17
10 16
11 15
12 14
13 13
14 12
15 11
16 10
17 9
18 8
19 7
20 6
7 20
8 19
9 18
10 17
11 16
12 15
13 14
14 13
15 12
16 11
17 10
18 9
19 8
20 7
8 20
9 19
10 18
11 17
12 16
13 15
14 14
15 13
16 12
17 11
18 10
19 9
20 8
9 20
10 19
11 18
12 17
13 16
14 15
15 14
16 13
17 12
18 11
19 10
20 9
10 20
11 19
12 18
13 17
14 16
15 15
16 14
17 13
18 12
19 11
20 10
11 20
12 19
13 18
14 17
15 16
16 15
17 14
18 13
19 12
20 11
12 20
13 19
14 18
15 17
16 16
17 15
18 14
19 13
20 12
13 20
14 19
15 18
16 17
17 16
18 15
19 14
20 13
14 20
15 19
16 18
17 17
18 16
19 15
20 14
15 20
16 19
17 18
18 17
19 16
20 15
16 20
17 19
18 18
19 17
20 16
17 20
18 19
19 18
20 17
18 20
19 19
20 18
19 20
20 19
20 20
.enddata

.end
