* 100x100 SRAM Array Netlist
.include "/home/taf27/hspice/libs/CMOS_180nm_L49.lib"
.include "sram_cell.sp"
.include "write_driver.sp"
.include "read_driver.sp"
.include "column_pull_up.sp"


*+++++++++++++++++++++++++++++++++
*++++++++++++SOURCES++++++++++++++
*+++++++++++++++++++++++++++++++++
Vdd vdd 0 1.8
Vss gnd 0 0
.param R_wl=0.5
.param C_wl=5.75f
Vwl_0 word_0 0 0
Rw0_0 word_0 word0_0 R_wl
Cwl_0_0 word0_0 gnd C_wl
Rw1_0 word1_0 word0_0 R_wl
Cwl_1_0 word1_0 gnd C_wl
Rw2_0 word2_0 word1_0 R_wl
Cwl_2_0 word2_0 gnd C_wl
Rw3_0 word3_0 word2_0 R_wl
Cwl_3_0 word3_0 gnd C_wl
Rw4_0 word4_0 word3_0 R_wl
Cwl_4_0 word4_0 gnd C_wl
Rw5_0 word5_0 word4_0 R_wl
Cwl_5_0 word5_0 gnd C_wl
Rw6_0 word6_0 word5_0 R_wl
Cwl_6_0 word6_0 gnd C_wl
Rw7_0 word7_0 word6_0 R_wl
Cwl_7_0 word7_0 gnd C_wl
Rw8_0 word8_0 word7_0 R_wl
Cwl_8_0 word8_0 gnd C_wl
Rw9_0 word9_0 word8_0 R_wl
Cwl_9_0 word9_0 gnd C_wl
Rw10_0 word10_0 word9_0 R_wl
Cwl_10_0 word10_0 gnd C_wl
Rw11_0 word11_0 word10_0 R_wl
Cwl_11_0 word11_0 gnd C_wl
Rw12_0 word12_0 word11_0 R_wl
Cwl_12_0 word12_0 gnd C_wl
Rw13_0 word13_0 word12_0 R_wl
Cwl_13_0 word13_0 gnd C_wl
Rw14_0 word14_0 word13_0 R_wl
Cwl_14_0 word14_0 gnd C_wl
Rw15_0 word15_0 word14_0 R_wl
Cwl_15_0 word15_0 gnd C_wl
Rw16_0 word16_0 word15_0 R_wl
Cwl_16_0 word16_0 gnd C_wl
Rw17_0 word17_0 word16_0 R_wl
Cwl_17_0 word17_0 gnd C_wl
Rw18_0 word18_0 word17_0 R_wl
Cwl_18_0 word18_0 gnd C_wl
Rw19_0 word19_0 word18_0 R_wl
Cwl_19_0 word19_0 gnd C_wl
Rw20_0 word20_0 word19_0 R_wl
Cwl_20_0 word20_0 gnd C_wl
Rw21_0 word21_0 word20_0 R_wl
Cwl_21_0 word21_0 gnd C_wl
Rw22_0 word22_0 word21_0 R_wl
Cwl_22_0 word22_0 gnd C_wl
Rw23_0 word23_0 word22_0 R_wl
Cwl_23_0 word23_0 gnd C_wl
Rw24_0 word24_0 word23_0 R_wl
Cwl_24_0 word24_0 gnd C_wl
Rw25_0 word25_0 word24_0 R_wl
Cwl_25_0 word25_0 gnd C_wl
Rw26_0 word26_0 word25_0 R_wl
Cwl_26_0 word26_0 gnd C_wl
Rw27_0 word27_0 word26_0 R_wl
Cwl_27_0 word27_0 gnd C_wl
Rw28_0 word28_0 word27_0 R_wl
Cwl_28_0 word28_0 gnd C_wl
Rw29_0 word29_0 word28_0 R_wl
Cwl_29_0 word29_0 gnd C_wl
Rw30_0 word30_0 word29_0 R_wl
Cwl_30_0 word30_0 gnd C_wl
Rw31_0 word31_0 word30_0 R_wl
Cwl_31_0 word31_0 gnd C_wl
Rw32_0 word32_0 word31_0 R_wl
Cwl_32_0 word32_0 gnd C_wl
Rw33_0 word33_0 word32_0 R_wl
Cwl_33_0 word33_0 gnd C_wl
Rw34_0 word34_0 word33_0 R_wl
Cwl_34_0 word34_0 gnd C_wl
Rw35_0 word35_0 word34_0 R_wl
Cwl_35_0 word35_0 gnd C_wl
Rw36_0 word36_0 word35_0 R_wl
Cwl_36_0 word36_0 gnd C_wl
Rw37_0 word37_0 word36_0 R_wl
Cwl_37_0 word37_0 gnd C_wl
Rw38_0 word38_0 word37_0 R_wl
Cwl_38_0 word38_0 gnd C_wl
Rw39_0 word39_0 word38_0 R_wl
Cwl_39_0 word39_0 gnd C_wl
Rw40_0 word40_0 word39_0 R_wl
Cwl_40_0 word40_0 gnd C_wl
Rw41_0 word41_0 word40_0 R_wl
Cwl_41_0 word41_0 gnd C_wl
Rw42_0 word42_0 word41_0 R_wl
Cwl_42_0 word42_0 gnd C_wl
Rw43_0 word43_0 word42_0 R_wl
Cwl_43_0 word43_0 gnd C_wl
Rw44_0 word44_0 word43_0 R_wl
Cwl_44_0 word44_0 gnd C_wl
Rw45_0 word45_0 word44_0 R_wl
Cwl_45_0 word45_0 gnd C_wl
Rw46_0 word46_0 word45_0 R_wl
Cwl_46_0 word46_0 gnd C_wl
Rw47_0 word47_0 word46_0 R_wl
Cwl_47_0 word47_0 gnd C_wl
Rw48_0 word48_0 word47_0 R_wl
Cwl_48_0 word48_0 gnd C_wl
Rw49_0 word49_0 word48_0 R_wl
Cwl_49_0 word49_0 gnd C_wl
Rw50_0 word50_0 word49_0 R_wl
Cwl_50_0 word50_0 gnd C_wl
Rw51_0 word51_0 word50_0 R_wl
Cwl_51_0 word51_0 gnd C_wl
Rw52_0 word52_0 word51_0 R_wl
Cwl_52_0 word52_0 gnd C_wl
Rw53_0 word53_0 word52_0 R_wl
Cwl_53_0 word53_0 gnd C_wl
Rw54_0 word54_0 word53_0 R_wl
Cwl_54_0 word54_0 gnd C_wl
Rw55_0 word55_0 word54_0 R_wl
Cwl_55_0 word55_0 gnd C_wl
Rw56_0 word56_0 word55_0 R_wl
Cwl_56_0 word56_0 gnd C_wl
Rw57_0 word57_0 word56_0 R_wl
Cwl_57_0 word57_0 gnd C_wl
Rw58_0 word58_0 word57_0 R_wl
Cwl_58_0 word58_0 gnd C_wl
Rw59_0 word59_0 word58_0 R_wl
Cwl_59_0 word59_0 gnd C_wl
Rw60_0 word60_0 word59_0 R_wl
Cwl_60_0 word60_0 gnd C_wl
Rw61_0 word61_0 word60_0 R_wl
Cwl_61_0 word61_0 gnd C_wl
Rw62_0 word62_0 word61_0 R_wl
Cwl_62_0 word62_0 gnd C_wl
Rw63_0 word63_0 word62_0 R_wl
Cwl_63_0 word63_0 gnd C_wl
Rw64_0 word64_0 word63_0 R_wl
Cwl_64_0 word64_0 gnd C_wl
Rw65_0 word65_0 word64_0 R_wl
Cwl_65_0 word65_0 gnd C_wl
Rw66_0 word66_0 word65_0 R_wl
Cwl_66_0 word66_0 gnd C_wl
Rw67_0 word67_0 word66_0 R_wl
Cwl_67_0 word67_0 gnd C_wl
Rw68_0 word68_0 word67_0 R_wl
Cwl_68_0 word68_0 gnd C_wl
Rw69_0 word69_0 word68_0 R_wl
Cwl_69_0 word69_0 gnd C_wl
Rw70_0 word70_0 word69_0 R_wl
Cwl_70_0 word70_0 gnd C_wl
Rw71_0 word71_0 word70_0 R_wl
Cwl_71_0 word71_0 gnd C_wl
Rw72_0 word72_0 word71_0 R_wl
Cwl_72_0 word72_0 gnd C_wl
Rw73_0 word73_0 word72_0 R_wl
Cwl_73_0 word73_0 gnd C_wl
Rw74_0 word74_0 word73_0 R_wl
Cwl_74_0 word74_0 gnd C_wl
Rw75_0 word75_0 word74_0 R_wl
Cwl_75_0 word75_0 gnd C_wl
Rw76_0 word76_0 word75_0 R_wl
Cwl_76_0 word76_0 gnd C_wl
Rw77_0 word77_0 word76_0 R_wl
Cwl_77_0 word77_0 gnd C_wl
Rw78_0 word78_0 word77_0 R_wl
Cwl_78_0 word78_0 gnd C_wl
Rw79_0 word79_0 word78_0 R_wl
Cwl_79_0 word79_0 gnd C_wl
Rw80_0 word80_0 word79_0 R_wl
Cwl_80_0 word80_0 gnd C_wl
Rw81_0 word81_0 word80_0 R_wl
Cwl_81_0 word81_0 gnd C_wl
Rw82_0 word82_0 word81_0 R_wl
Cwl_82_0 word82_0 gnd C_wl
Rw83_0 word83_0 word82_0 R_wl
Cwl_83_0 word83_0 gnd C_wl
Rw84_0 word84_0 word83_0 R_wl
Cwl_84_0 word84_0 gnd C_wl
Rw85_0 word85_0 word84_0 R_wl
Cwl_85_0 word85_0 gnd C_wl
Rw86_0 word86_0 word85_0 R_wl
Cwl_86_0 word86_0 gnd C_wl
Rw87_0 word87_0 word86_0 R_wl
Cwl_87_0 word87_0 gnd C_wl
Rw88_0 word88_0 word87_0 R_wl
Cwl_88_0 word88_0 gnd C_wl
Rw89_0 word89_0 word88_0 R_wl
Cwl_89_0 word89_0 gnd C_wl
Rw90_0 word90_0 word89_0 R_wl
Cwl_90_0 word90_0 gnd C_wl
Rw91_0 word91_0 word90_0 R_wl
Cwl_91_0 word91_0 gnd C_wl
Rw92_0 word92_0 word91_0 R_wl
Cwl_92_0 word92_0 gnd C_wl
Rw93_0 word93_0 word92_0 R_wl
Cwl_93_0 word93_0 gnd C_wl
Rw94_0 word94_0 word93_0 R_wl
Cwl_94_0 word94_0 gnd C_wl
Rw95_0 word95_0 word94_0 R_wl
Cwl_95_0 word95_0 gnd C_wl
Rw96_0 word96_0 word95_0 R_wl
Cwl_96_0 word96_0 gnd C_wl
Rw97_0 word97_0 word96_0 R_wl
Cwl_97_0 word97_0 gnd C_wl
Rw98_0 word98_0 word97_0 R_wl
Cwl_98_0 word98_0 gnd C_wl
Rw99_0 word99_0 word98_0 R_wl
Cwl_99_0 word99_0 gnd C_wl
Vwl_1 word_1 0 0
Rw0_1 word_1 word0_1 R_wl
Cwl_0_1 word0_1 gnd C_wl
Rw1_1 word1_1 word0_1 R_wl
Cwl_1_1 word1_1 gnd C_wl
Rw2_1 word2_1 word1_1 R_wl
Cwl_2_1 word2_1 gnd C_wl
Rw3_1 word3_1 word2_1 R_wl
Cwl_3_1 word3_1 gnd C_wl
Rw4_1 word4_1 word3_1 R_wl
Cwl_4_1 word4_1 gnd C_wl
Rw5_1 word5_1 word4_1 R_wl
Cwl_5_1 word5_1 gnd C_wl
Rw6_1 word6_1 word5_1 R_wl
Cwl_6_1 word6_1 gnd C_wl
Rw7_1 word7_1 word6_1 R_wl
Cwl_7_1 word7_1 gnd C_wl
Rw8_1 word8_1 word7_1 R_wl
Cwl_8_1 word8_1 gnd C_wl
Rw9_1 word9_1 word8_1 R_wl
Cwl_9_1 word9_1 gnd C_wl
Rw10_1 word10_1 word9_1 R_wl
Cwl_10_1 word10_1 gnd C_wl
Rw11_1 word11_1 word10_1 R_wl
Cwl_11_1 word11_1 gnd C_wl
Rw12_1 word12_1 word11_1 R_wl
Cwl_12_1 word12_1 gnd C_wl
Rw13_1 word13_1 word12_1 R_wl
Cwl_13_1 word13_1 gnd C_wl
Rw14_1 word14_1 word13_1 R_wl
Cwl_14_1 word14_1 gnd C_wl
Rw15_1 word15_1 word14_1 R_wl
Cwl_15_1 word15_1 gnd C_wl
Rw16_1 word16_1 word15_1 R_wl
Cwl_16_1 word16_1 gnd C_wl
Rw17_1 word17_1 word16_1 R_wl
Cwl_17_1 word17_1 gnd C_wl
Rw18_1 word18_1 word17_1 R_wl
Cwl_18_1 word18_1 gnd C_wl
Rw19_1 word19_1 word18_1 R_wl
Cwl_19_1 word19_1 gnd C_wl
Rw20_1 word20_1 word19_1 R_wl
Cwl_20_1 word20_1 gnd C_wl
Rw21_1 word21_1 word20_1 R_wl
Cwl_21_1 word21_1 gnd C_wl
Rw22_1 word22_1 word21_1 R_wl
Cwl_22_1 word22_1 gnd C_wl
Rw23_1 word23_1 word22_1 R_wl
Cwl_23_1 word23_1 gnd C_wl
Rw24_1 word24_1 word23_1 R_wl
Cwl_24_1 word24_1 gnd C_wl
Rw25_1 word25_1 word24_1 R_wl
Cwl_25_1 word25_1 gnd C_wl
Rw26_1 word26_1 word25_1 R_wl
Cwl_26_1 word26_1 gnd C_wl
Rw27_1 word27_1 word26_1 R_wl
Cwl_27_1 word27_1 gnd C_wl
Rw28_1 word28_1 word27_1 R_wl
Cwl_28_1 word28_1 gnd C_wl
Rw29_1 word29_1 word28_1 R_wl
Cwl_29_1 word29_1 gnd C_wl
Rw30_1 word30_1 word29_1 R_wl
Cwl_30_1 word30_1 gnd C_wl
Rw31_1 word31_1 word30_1 R_wl
Cwl_31_1 word31_1 gnd C_wl
Rw32_1 word32_1 word31_1 R_wl
Cwl_32_1 word32_1 gnd C_wl
Rw33_1 word33_1 word32_1 R_wl
Cwl_33_1 word33_1 gnd C_wl
Rw34_1 word34_1 word33_1 R_wl
Cwl_34_1 word34_1 gnd C_wl
Rw35_1 word35_1 word34_1 R_wl
Cwl_35_1 word35_1 gnd C_wl
Rw36_1 word36_1 word35_1 R_wl
Cwl_36_1 word36_1 gnd C_wl
Rw37_1 word37_1 word36_1 R_wl
Cwl_37_1 word37_1 gnd C_wl
Rw38_1 word38_1 word37_1 R_wl
Cwl_38_1 word38_1 gnd C_wl
Rw39_1 word39_1 word38_1 R_wl
Cwl_39_1 word39_1 gnd C_wl
Rw40_1 word40_1 word39_1 R_wl
Cwl_40_1 word40_1 gnd C_wl
Rw41_1 word41_1 word40_1 R_wl
Cwl_41_1 word41_1 gnd C_wl
Rw42_1 word42_1 word41_1 R_wl
Cwl_42_1 word42_1 gnd C_wl
Rw43_1 word43_1 word42_1 R_wl
Cwl_43_1 word43_1 gnd C_wl
Rw44_1 word44_1 word43_1 R_wl
Cwl_44_1 word44_1 gnd C_wl
Rw45_1 word45_1 word44_1 R_wl
Cwl_45_1 word45_1 gnd C_wl
Rw46_1 word46_1 word45_1 R_wl
Cwl_46_1 word46_1 gnd C_wl
Rw47_1 word47_1 word46_1 R_wl
Cwl_47_1 word47_1 gnd C_wl
Rw48_1 word48_1 word47_1 R_wl
Cwl_48_1 word48_1 gnd C_wl
Rw49_1 word49_1 word48_1 R_wl
Cwl_49_1 word49_1 gnd C_wl
Rw50_1 word50_1 word49_1 R_wl
Cwl_50_1 word50_1 gnd C_wl
Rw51_1 word51_1 word50_1 R_wl
Cwl_51_1 word51_1 gnd C_wl
Rw52_1 word52_1 word51_1 R_wl
Cwl_52_1 word52_1 gnd C_wl
Rw53_1 word53_1 word52_1 R_wl
Cwl_53_1 word53_1 gnd C_wl
Rw54_1 word54_1 word53_1 R_wl
Cwl_54_1 word54_1 gnd C_wl
Rw55_1 word55_1 word54_1 R_wl
Cwl_55_1 word55_1 gnd C_wl
Rw56_1 word56_1 word55_1 R_wl
Cwl_56_1 word56_1 gnd C_wl
Rw57_1 word57_1 word56_1 R_wl
Cwl_57_1 word57_1 gnd C_wl
Rw58_1 word58_1 word57_1 R_wl
Cwl_58_1 word58_1 gnd C_wl
Rw59_1 word59_1 word58_1 R_wl
Cwl_59_1 word59_1 gnd C_wl
Rw60_1 word60_1 word59_1 R_wl
Cwl_60_1 word60_1 gnd C_wl
Rw61_1 word61_1 word60_1 R_wl
Cwl_61_1 word61_1 gnd C_wl
Rw62_1 word62_1 word61_1 R_wl
Cwl_62_1 word62_1 gnd C_wl
Rw63_1 word63_1 word62_1 R_wl
Cwl_63_1 word63_1 gnd C_wl
Rw64_1 word64_1 word63_1 R_wl
Cwl_64_1 word64_1 gnd C_wl
Rw65_1 word65_1 word64_1 R_wl
Cwl_65_1 word65_1 gnd C_wl
Rw66_1 word66_1 word65_1 R_wl
Cwl_66_1 word66_1 gnd C_wl
Rw67_1 word67_1 word66_1 R_wl
Cwl_67_1 word67_1 gnd C_wl
Rw68_1 word68_1 word67_1 R_wl
Cwl_68_1 word68_1 gnd C_wl
Rw69_1 word69_1 word68_1 R_wl
Cwl_69_1 word69_1 gnd C_wl
Rw70_1 word70_1 word69_1 R_wl
Cwl_70_1 word70_1 gnd C_wl
Rw71_1 word71_1 word70_1 R_wl
Cwl_71_1 word71_1 gnd C_wl
Rw72_1 word72_1 word71_1 R_wl
Cwl_72_1 word72_1 gnd C_wl
Rw73_1 word73_1 word72_1 R_wl
Cwl_73_1 word73_1 gnd C_wl
Rw74_1 word74_1 word73_1 R_wl
Cwl_74_1 word74_1 gnd C_wl
Rw75_1 word75_1 word74_1 R_wl
Cwl_75_1 word75_1 gnd C_wl
Rw76_1 word76_1 word75_1 R_wl
Cwl_76_1 word76_1 gnd C_wl
Rw77_1 word77_1 word76_1 R_wl
Cwl_77_1 word77_1 gnd C_wl
Rw78_1 word78_1 word77_1 R_wl
Cwl_78_1 word78_1 gnd C_wl
Rw79_1 word79_1 word78_1 R_wl
Cwl_79_1 word79_1 gnd C_wl
Rw80_1 word80_1 word79_1 R_wl
Cwl_80_1 word80_1 gnd C_wl
Rw81_1 word81_1 word80_1 R_wl
Cwl_81_1 word81_1 gnd C_wl
Rw82_1 word82_1 word81_1 R_wl
Cwl_82_1 word82_1 gnd C_wl
Rw83_1 word83_1 word82_1 R_wl
Cwl_83_1 word83_1 gnd C_wl
Rw84_1 word84_1 word83_1 R_wl
Cwl_84_1 word84_1 gnd C_wl
Rw85_1 word85_1 word84_1 R_wl
Cwl_85_1 word85_1 gnd C_wl
Rw86_1 word86_1 word85_1 R_wl
Cwl_86_1 word86_1 gnd C_wl
Rw87_1 word87_1 word86_1 R_wl
Cwl_87_1 word87_1 gnd C_wl
Rw88_1 word88_1 word87_1 R_wl
Cwl_88_1 word88_1 gnd C_wl
Rw89_1 word89_1 word88_1 R_wl
Cwl_89_1 word89_1 gnd C_wl
Rw90_1 word90_1 word89_1 R_wl
Cwl_90_1 word90_1 gnd C_wl
Rw91_1 word91_1 word90_1 R_wl
Cwl_91_1 word91_1 gnd C_wl
Rw92_1 word92_1 word91_1 R_wl
Cwl_92_1 word92_1 gnd C_wl
Rw93_1 word93_1 word92_1 R_wl
Cwl_93_1 word93_1 gnd C_wl
Rw94_1 word94_1 word93_1 R_wl
Cwl_94_1 word94_1 gnd C_wl
Rw95_1 word95_1 word94_1 R_wl
Cwl_95_1 word95_1 gnd C_wl
Rw96_1 word96_1 word95_1 R_wl
Cwl_96_1 word96_1 gnd C_wl
Rw97_1 word97_1 word96_1 R_wl
Cwl_97_1 word97_1 gnd C_wl
Rw98_1 word98_1 word97_1 R_wl
Cwl_98_1 word98_1 gnd C_wl
Rw99_1 word99_1 word98_1 R_wl
Cwl_99_1 word99_1 gnd C_wl
Vwl_2 word_2 0 0
Rw0_2 word_2 word0_2 R_wl
Cwl_0_2 word0_2 gnd C_wl
Rw1_2 word1_2 word0_2 R_wl
Cwl_1_2 word1_2 gnd C_wl
Rw2_2 word2_2 word1_2 R_wl
Cwl_2_2 word2_2 gnd C_wl
Rw3_2 word3_2 word2_2 R_wl
Cwl_3_2 word3_2 gnd C_wl
Rw4_2 word4_2 word3_2 R_wl
Cwl_4_2 word4_2 gnd C_wl
Rw5_2 word5_2 word4_2 R_wl
Cwl_5_2 word5_2 gnd C_wl
Rw6_2 word6_2 word5_2 R_wl
Cwl_6_2 word6_2 gnd C_wl
Rw7_2 word7_2 word6_2 R_wl
Cwl_7_2 word7_2 gnd C_wl
Rw8_2 word8_2 word7_2 R_wl
Cwl_8_2 word8_2 gnd C_wl
Rw9_2 word9_2 word8_2 R_wl
Cwl_9_2 word9_2 gnd C_wl
Rw10_2 word10_2 word9_2 R_wl
Cwl_10_2 word10_2 gnd C_wl
Rw11_2 word11_2 word10_2 R_wl
Cwl_11_2 word11_2 gnd C_wl
Rw12_2 word12_2 word11_2 R_wl
Cwl_12_2 word12_2 gnd C_wl
Rw13_2 word13_2 word12_2 R_wl
Cwl_13_2 word13_2 gnd C_wl
Rw14_2 word14_2 word13_2 R_wl
Cwl_14_2 word14_2 gnd C_wl
Rw15_2 word15_2 word14_2 R_wl
Cwl_15_2 word15_2 gnd C_wl
Rw16_2 word16_2 word15_2 R_wl
Cwl_16_2 word16_2 gnd C_wl
Rw17_2 word17_2 word16_2 R_wl
Cwl_17_2 word17_2 gnd C_wl
Rw18_2 word18_2 word17_2 R_wl
Cwl_18_2 word18_2 gnd C_wl
Rw19_2 word19_2 word18_2 R_wl
Cwl_19_2 word19_2 gnd C_wl
Rw20_2 word20_2 word19_2 R_wl
Cwl_20_2 word20_2 gnd C_wl
Rw21_2 word21_2 word20_2 R_wl
Cwl_21_2 word21_2 gnd C_wl
Rw22_2 word22_2 word21_2 R_wl
Cwl_22_2 word22_2 gnd C_wl
Rw23_2 word23_2 word22_2 R_wl
Cwl_23_2 word23_2 gnd C_wl
Rw24_2 word24_2 word23_2 R_wl
Cwl_24_2 word24_2 gnd C_wl
Rw25_2 word25_2 word24_2 R_wl
Cwl_25_2 word25_2 gnd C_wl
Rw26_2 word26_2 word25_2 R_wl
Cwl_26_2 word26_2 gnd C_wl
Rw27_2 word27_2 word26_2 R_wl
Cwl_27_2 word27_2 gnd C_wl
Rw28_2 word28_2 word27_2 R_wl
Cwl_28_2 word28_2 gnd C_wl
Rw29_2 word29_2 word28_2 R_wl
Cwl_29_2 word29_2 gnd C_wl
Rw30_2 word30_2 word29_2 R_wl
Cwl_30_2 word30_2 gnd C_wl
Rw31_2 word31_2 word30_2 R_wl
Cwl_31_2 word31_2 gnd C_wl
Rw32_2 word32_2 word31_2 R_wl
Cwl_32_2 word32_2 gnd C_wl
Rw33_2 word33_2 word32_2 R_wl
Cwl_33_2 word33_2 gnd C_wl
Rw34_2 word34_2 word33_2 R_wl
Cwl_34_2 word34_2 gnd C_wl
Rw35_2 word35_2 word34_2 R_wl
Cwl_35_2 word35_2 gnd C_wl
Rw36_2 word36_2 word35_2 R_wl
Cwl_36_2 word36_2 gnd C_wl
Rw37_2 word37_2 word36_2 R_wl
Cwl_37_2 word37_2 gnd C_wl
Rw38_2 word38_2 word37_2 R_wl
Cwl_38_2 word38_2 gnd C_wl
Rw39_2 word39_2 word38_2 R_wl
Cwl_39_2 word39_2 gnd C_wl
Rw40_2 word40_2 word39_2 R_wl
Cwl_40_2 word40_2 gnd C_wl
Rw41_2 word41_2 word40_2 R_wl
Cwl_41_2 word41_2 gnd C_wl
Rw42_2 word42_2 word41_2 R_wl
Cwl_42_2 word42_2 gnd C_wl
Rw43_2 word43_2 word42_2 R_wl
Cwl_43_2 word43_2 gnd C_wl
Rw44_2 word44_2 word43_2 R_wl
Cwl_44_2 word44_2 gnd C_wl
Rw45_2 word45_2 word44_2 R_wl
Cwl_45_2 word45_2 gnd C_wl
Rw46_2 word46_2 word45_2 R_wl
Cwl_46_2 word46_2 gnd C_wl
Rw47_2 word47_2 word46_2 R_wl
Cwl_47_2 word47_2 gnd C_wl
Rw48_2 word48_2 word47_2 R_wl
Cwl_48_2 word48_2 gnd C_wl
Rw49_2 word49_2 word48_2 R_wl
Cwl_49_2 word49_2 gnd C_wl
Rw50_2 word50_2 word49_2 R_wl
Cwl_50_2 word50_2 gnd C_wl
Rw51_2 word51_2 word50_2 R_wl
Cwl_51_2 word51_2 gnd C_wl
Rw52_2 word52_2 word51_2 R_wl
Cwl_52_2 word52_2 gnd C_wl
Rw53_2 word53_2 word52_2 R_wl
Cwl_53_2 word53_2 gnd C_wl
Rw54_2 word54_2 word53_2 R_wl
Cwl_54_2 word54_2 gnd C_wl
Rw55_2 word55_2 word54_2 R_wl
Cwl_55_2 word55_2 gnd C_wl
Rw56_2 word56_2 word55_2 R_wl
Cwl_56_2 word56_2 gnd C_wl
Rw57_2 word57_2 word56_2 R_wl
Cwl_57_2 word57_2 gnd C_wl
Rw58_2 word58_2 word57_2 R_wl
Cwl_58_2 word58_2 gnd C_wl
Rw59_2 word59_2 word58_2 R_wl
Cwl_59_2 word59_2 gnd C_wl
Rw60_2 word60_2 word59_2 R_wl
Cwl_60_2 word60_2 gnd C_wl
Rw61_2 word61_2 word60_2 R_wl
Cwl_61_2 word61_2 gnd C_wl
Rw62_2 word62_2 word61_2 R_wl
Cwl_62_2 word62_2 gnd C_wl
Rw63_2 word63_2 word62_2 R_wl
Cwl_63_2 word63_2 gnd C_wl
Rw64_2 word64_2 word63_2 R_wl
Cwl_64_2 word64_2 gnd C_wl
Rw65_2 word65_2 word64_2 R_wl
Cwl_65_2 word65_2 gnd C_wl
Rw66_2 word66_2 word65_2 R_wl
Cwl_66_2 word66_2 gnd C_wl
Rw67_2 word67_2 word66_2 R_wl
Cwl_67_2 word67_2 gnd C_wl
Rw68_2 word68_2 word67_2 R_wl
Cwl_68_2 word68_2 gnd C_wl
Rw69_2 word69_2 word68_2 R_wl
Cwl_69_2 word69_2 gnd C_wl
Rw70_2 word70_2 word69_2 R_wl
Cwl_70_2 word70_2 gnd C_wl
Rw71_2 word71_2 word70_2 R_wl
Cwl_71_2 word71_2 gnd C_wl
Rw72_2 word72_2 word71_2 R_wl
Cwl_72_2 word72_2 gnd C_wl
Rw73_2 word73_2 word72_2 R_wl
Cwl_73_2 word73_2 gnd C_wl
Rw74_2 word74_2 word73_2 R_wl
Cwl_74_2 word74_2 gnd C_wl
Rw75_2 word75_2 word74_2 R_wl
Cwl_75_2 word75_2 gnd C_wl
Rw76_2 word76_2 word75_2 R_wl
Cwl_76_2 word76_2 gnd C_wl
Rw77_2 word77_2 word76_2 R_wl
Cwl_77_2 word77_2 gnd C_wl
Rw78_2 word78_2 word77_2 R_wl
Cwl_78_2 word78_2 gnd C_wl
Rw79_2 word79_2 word78_2 R_wl
Cwl_79_2 word79_2 gnd C_wl
Rw80_2 word80_2 word79_2 R_wl
Cwl_80_2 word80_2 gnd C_wl
Rw81_2 word81_2 word80_2 R_wl
Cwl_81_2 word81_2 gnd C_wl
Rw82_2 word82_2 word81_2 R_wl
Cwl_82_2 word82_2 gnd C_wl
Rw83_2 word83_2 word82_2 R_wl
Cwl_83_2 word83_2 gnd C_wl
Rw84_2 word84_2 word83_2 R_wl
Cwl_84_2 word84_2 gnd C_wl
Rw85_2 word85_2 word84_2 R_wl
Cwl_85_2 word85_2 gnd C_wl
Rw86_2 word86_2 word85_2 R_wl
Cwl_86_2 word86_2 gnd C_wl
Rw87_2 word87_2 word86_2 R_wl
Cwl_87_2 word87_2 gnd C_wl
Rw88_2 word88_2 word87_2 R_wl
Cwl_88_2 word88_2 gnd C_wl
Rw89_2 word89_2 word88_2 R_wl
Cwl_89_2 word89_2 gnd C_wl
Rw90_2 word90_2 word89_2 R_wl
Cwl_90_2 word90_2 gnd C_wl
Rw91_2 word91_2 word90_2 R_wl
Cwl_91_2 word91_2 gnd C_wl
Rw92_2 word92_2 word91_2 R_wl
Cwl_92_2 word92_2 gnd C_wl
Rw93_2 word93_2 word92_2 R_wl
Cwl_93_2 word93_2 gnd C_wl
Rw94_2 word94_2 word93_2 R_wl
Cwl_94_2 word94_2 gnd C_wl
Rw95_2 word95_2 word94_2 R_wl
Cwl_95_2 word95_2 gnd C_wl
Rw96_2 word96_2 word95_2 R_wl
Cwl_96_2 word96_2 gnd C_wl
Rw97_2 word97_2 word96_2 R_wl
Cwl_97_2 word97_2 gnd C_wl
Rw98_2 word98_2 word97_2 R_wl
Cwl_98_2 word98_2 gnd C_wl
Rw99_2 word99_2 word98_2 R_wl
Cwl_99_2 word99_2 gnd C_wl
Vwl_3 word_3 0 0
Rw0_3 word_3 word0_3 R_wl
Cwl_0_3 word0_3 gnd C_wl
Rw1_3 word1_3 word0_3 R_wl
Cwl_1_3 word1_3 gnd C_wl
Rw2_3 word2_3 word1_3 R_wl
Cwl_2_3 word2_3 gnd C_wl
Rw3_3 word3_3 word2_3 R_wl
Cwl_3_3 word3_3 gnd C_wl
Rw4_3 word4_3 word3_3 R_wl
Cwl_4_3 word4_3 gnd C_wl
Rw5_3 word5_3 word4_3 R_wl
Cwl_5_3 word5_3 gnd C_wl
Rw6_3 word6_3 word5_3 R_wl
Cwl_6_3 word6_3 gnd C_wl
Rw7_3 word7_3 word6_3 R_wl
Cwl_7_3 word7_3 gnd C_wl
Rw8_3 word8_3 word7_3 R_wl
Cwl_8_3 word8_3 gnd C_wl
Rw9_3 word9_3 word8_3 R_wl
Cwl_9_3 word9_3 gnd C_wl
Rw10_3 word10_3 word9_3 R_wl
Cwl_10_3 word10_3 gnd C_wl
Rw11_3 word11_3 word10_3 R_wl
Cwl_11_3 word11_3 gnd C_wl
Rw12_3 word12_3 word11_3 R_wl
Cwl_12_3 word12_3 gnd C_wl
Rw13_3 word13_3 word12_3 R_wl
Cwl_13_3 word13_3 gnd C_wl
Rw14_3 word14_3 word13_3 R_wl
Cwl_14_3 word14_3 gnd C_wl
Rw15_3 word15_3 word14_3 R_wl
Cwl_15_3 word15_3 gnd C_wl
Rw16_3 word16_3 word15_3 R_wl
Cwl_16_3 word16_3 gnd C_wl
Rw17_3 word17_3 word16_3 R_wl
Cwl_17_3 word17_3 gnd C_wl
Rw18_3 word18_3 word17_3 R_wl
Cwl_18_3 word18_3 gnd C_wl
Rw19_3 word19_3 word18_3 R_wl
Cwl_19_3 word19_3 gnd C_wl
Rw20_3 word20_3 word19_3 R_wl
Cwl_20_3 word20_3 gnd C_wl
Rw21_3 word21_3 word20_3 R_wl
Cwl_21_3 word21_3 gnd C_wl
Rw22_3 word22_3 word21_3 R_wl
Cwl_22_3 word22_3 gnd C_wl
Rw23_3 word23_3 word22_3 R_wl
Cwl_23_3 word23_3 gnd C_wl
Rw24_3 word24_3 word23_3 R_wl
Cwl_24_3 word24_3 gnd C_wl
Rw25_3 word25_3 word24_3 R_wl
Cwl_25_3 word25_3 gnd C_wl
Rw26_3 word26_3 word25_3 R_wl
Cwl_26_3 word26_3 gnd C_wl
Rw27_3 word27_3 word26_3 R_wl
Cwl_27_3 word27_3 gnd C_wl
Rw28_3 word28_3 word27_3 R_wl
Cwl_28_3 word28_3 gnd C_wl
Rw29_3 word29_3 word28_3 R_wl
Cwl_29_3 word29_3 gnd C_wl
Rw30_3 word30_3 word29_3 R_wl
Cwl_30_3 word30_3 gnd C_wl
Rw31_3 word31_3 word30_3 R_wl
Cwl_31_3 word31_3 gnd C_wl
Rw32_3 word32_3 word31_3 R_wl
Cwl_32_3 word32_3 gnd C_wl
Rw33_3 word33_3 word32_3 R_wl
Cwl_33_3 word33_3 gnd C_wl
Rw34_3 word34_3 word33_3 R_wl
Cwl_34_3 word34_3 gnd C_wl
Rw35_3 word35_3 word34_3 R_wl
Cwl_35_3 word35_3 gnd C_wl
Rw36_3 word36_3 word35_3 R_wl
Cwl_36_3 word36_3 gnd C_wl
Rw37_3 word37_3 word36_3 R_wl
Cwl_37_3 word37_3 gnd C_wl
Rw38_3 word38_3 word37_3 R_wl
Cwl_38_3 word38_3 gnd C_wl
Rw39_3 word39_3 word38_3 R_wl
Cwl_39_3 word39_3 gnd C_wl
Rw40_3 word40_3 word39_3 R_wl
Cwl_40_3 word40_3 gnd C_wl
Rw41_3 word41_3 word40_3 R_wl
Cwl_41_3 word41_3 gnd C_wl
Rw42_3 word42_3 word41_3 R_wl
Cwl_42_3 word42_3 gnd C_wl
Rw43_3 word43_3 word42_3 R_wl
Cwl_43_3 word43_3 gnd C_wl
Rw44_3 word44_3 word43_3 R_wl
Cwl_44_3 word44_3 gnd C_wl
Rw45_3 word45_3 word44_3 R_wl
Cwl_45_3 word45_3 gnd C_wl
Rw46_3 word46_3 word45_3 R_wl
Cwl_46_3 word46_3 gnd C_wl
Rw47_3 word47_3 word46_3 R_wl
Cwl_47_3 word47_3 gnd C_wl
Rw48_3 word48_3 word47_3 R_wl
Cwl_48_3 word48_3 gnd C_wl
Rw49_3 word49_3 word48_3 R_wl
Cwl_49_3 word49_3 gnd C_wl
Rw50_3 word50_3 word49_3 R_wl
Cwl_50_3 word50_3 gnd C_wl
Rw51_3 word51_3 word50_3 R_wl
Cwl_51_3 word51_3 gnd C_wl
Rw52_3 word52_3 word51_3 R_wl
Cwl_52_3 word52_3 gnd C_wl
Rw53_3 word53_3 word52_3 R_wl
Cwl_53_3 word53_3 gnd C_wl
Rw54_3 word54_3 word53_3 R_wl
Cwl_54_3 word54_3 gnd C_wl
Rw55_3 word55_3 word54_3 R_wl
Cwl_55_3 word55_3 gnd C_wl
Rw56_3 word56_3 word55_3 R_wl
Cwl_56_3 word56_3 gnd C_wl
Rw57_3 word57_3 word56_3 R_wl
Cwl_57_3 word57_3 gnd C_wl
Rw58_3 word58_3 word57_3 R_wl
Cwl_58_3 word58_3 gnd C_wl
Rw59_3 word59_3 word58_3 R_wl
Cwl_59_3 word59_3 gnd C_wl
Rw60_3 word60_3 word59_3 R_wl
Cwl_60_3 word60_3 gnd C_wl
Rw61_3 word61_3 word60_3 R_wl
Cwl_61_3 word61_3 gnd C_wl
Rw62_3 word62_3 word61_3 R_wl
Cwl_62_3 word62_3 gnd C_wl
Rw63_3 word63_3 word62_3 R_wl
Cwl_63_3 word63_3 gnd C_wl
Rw64_3 word64_3 word63_3 R_wl
Cwl_64_3 word64_3 gnd C_wl
Rw65_3 word65_3 word64_3 R_wl
Cwl_65_3 word65_3 gnd C_wl
Rw66_3 word66_3 word65_3 R_wl
Cwl_66_3 word66_3 gnd C_wl
Rw67_3 word67_3 word66_3 R_wl
Cwl_67_3 word67_3 gnd C_wl
Rw68_3 word68_3 word67_3 R_wl
Cwl_68_3 word68_3 gnd C_wl
Rw69_3 word69_3 word68_3 R_wl
Cwl_69_3 word69_3 gnd C_wl
Rw70_3 word70_3 word69_3 R_wl
Cwl_70_3 word70_3 gnd C_wl
Rw71_3 word71_3 word70_3 R_wl
Cwl_71_3 word71_3 gnd C_wl
Rw72_3 word72_3 word71_3 R_wl
Cwl_72_3 word72_3 gnd C_wl
Rw73_3 word73_3 word72_3 R_wl
Cwl_73_3 word73_3 gnd C_wl
Rw74_3 word74_3 word73_3 R_wl
Cwl_74_3 word74_3 gnd C_wl
Rw75_3 word75_3 word74_3 R_wl
Cwl_75_3 word75_3 gnd C_wl
Rw76_3 word76_3 word75_3 R_wl
Cwl_76_3 word76_3 gnd C_wl
Rw77_3 word77_3 word76_3 R_wl
Cwl_77_3 word77_3 gnd C_wl
Rw78_3 word78_3 word77_3 R_wl
Cwl_78_3 word78_3 gnd C_wl
Rw79_3 word79_3 word78_3 R_wl
Cwl_79_3 word79_3 gnd C_wl
Rw80_3 word80_3 word79_3 R_wl
Cwl_80_3 word80_3 gnd C_wl
Rw81_3 word81_3 word80_3 R_wl
Cwl_81_3 word81_3 gnd C_wl
Rw82_3 word82_3 word81_3 R_wl
Cwl_82_3 word82_3 gnd C_wl
Rw83_3 word83_3 word82_3 R_wl
Cwl_83_3 word83_3 gnd C_wl
Rw84_3 word84_3 word83_3 R_wl
Cwl_84_3 word84_3 gnd C_wl
Rw85_3 word85_3 word84_3 R_wl
Cwl_85_3 word85_3 gnd C_wl
Rw86_3 word86_3 word85_3 R_wl
Cwl_86_3 word86_3 gnd C_wl
Rw87_3 word87_3 word86_3 R_wl
Cwl_87_3 word87_3 gnd C_wl
Rw88_3 word88_3 word87_3 R_wl
Cwl_88_3 word88_3 gnd C_wl
Rw89_3 word89_3 word88_3 R_wl
Cwl_89_3 word89_3 gnd C_wl
Rw90_3 word90_3 word89_3 R_wl
Cwl_90_3 word90_3 gnd C_wl
Rw91_3 word91_3 word90_3 R_wl
Cwl_91_3 word91_3 gnd C_wl
Rw92_3 word92_3 word91_3 R_wl
Cwl_92_3 word92_3 gnd C_wl
Rw93_3 word93_3 word92_3 R_wl
Cwl_93_3 word93_3 gnd C_wl
Rw94_3 word94_3 word93_3 R_wl
Cwl_94_3 word94_3 gnd C_wl
Rw95_3 word95_3 word94_3 R_wl
Cwl_95_3 word95_3 gnd C_wl
Rw96_3 word96_3 word95_3 R_wl
Cwl_96_3 word96_3 gnd C_wl
Rw97_3 word97_3 word96_3 R_wl
Cwl_97_3 word97_3 gnd C_wl
Rw98_3 word98_3 word97_3 R_wl
Cwl_98_3 word98_3 gnd C_wl
Rw99_3 word99_3 word98_3 R_wl
Cwl_99_3 word99_3 gnd C_wl
Vwl_4 word_4 0 0
Rw0_4 word_4 word0_4 R_wl
Cwl_0_4 word0_4 gnd C_wl
Rw1_4 word1_4 word0_4 R_wl
Cwl_1_4 word1_4 gnd C_wl
Rw2_4 word2_4 word1_4 R_wl
Cwl_2_4 word2_4 gnd C_wl
Rw3_4 word3_4 word2_4 R_wl
Cwl_3_4 word3_4 gnd C_wl
Rw4_4 word4_4 word3_4 R_wl
Cwl_4_4 word4_4 gnd C_wl
Rw5_4 word5_4 word4_4 R_wl
Cwl_5_4 word5_4 gnd C_wl
Rw6_4 word6_4 word5_4 R_wl
Cwl_6_4 word6_4 gnd C_wl
Rw7_4 word7_4 word6_4 R_wl
Cwl_7_4 word7_4 gnd C_wl
Rw8_4 word8_4 word7_4 R_wl
Cwl_8_4 word8_4 gnd C_wl
Rw9_4 word9_4 word8_4 R_wl
Cwl_9_4 word9_4 gnd C_wl
Rw10_4 word10_4 word9_4 R_wl
Cwl_10_4 word10_4 gnd C_wl
Rw11_4 word11_4 word10_4 R_wl
Cwl_11_4 word11_4 gnd C_wl
Rw12_4 word12_4 word11_4 R_wl
Cwl_12_4 word12_4 gnd C_wl
Rw13_4 word13_4 word12_4 R_wl
Cwl_13_4 word13_4 gnd C_wl
Rw14_4 word14_4 word13_4 R_wl
Cwl_14_4 word14_4 gnd C_wl
Rw15_4 word15_4 word14_4 R_wl
Cwl_15_4 word15_4 gnd C_wl
Rw16_4 word16_4 word15_4 R_wl
Cwl_16_4 word16_4 gnd C_wl
Rw17_4 word17_4 word16_4 R_wl
Cwl_17_4 word17_4 gnd C_wl
Rw18_4 word18_4 word17_4 R_wl
Cwl_18_4 word18_4 gnd C_wl
Rw19_4 word19_4 word18_4 R_wl
Cwl_19_4 word19_4 gnd C_wl
Rw20_4 word20_4 word19_4 R_wl
Cwl_20_4 word20_4 gnd C_wl
Rw21_4 word21_4 word20_4 R_wl
Cwl_21_4 word21_4 gnd C_wl
Rw22_4 word22_4 word21_4 R_wl
Cwl_22_4 word22_4 gnd C_wl
Rw23_4 word23_4 word22_4 R_wl
Cwl_23_4 word23_4 gnd C_wl
Rw24_4 word24_4 word23_4 R_wl
Cwl_24_4 word24_4 gnd C_wl
Rw25_4 word25_4 word24_4 R_wl
Cwl_25_4 word25_4 gnd C_wl
Rw26_4 word26_4 word25_4 R_wl
Cwl_26_4 word26_4 gnd C_wl
Rw27_4 word27_4 word26_4 R_wl
Cwl_27_4 word27_4 gnd C_wl
Rw28_4 word28_4 word27_4 R_wl
Cwl_28_4 word28_4 gnd C_wl
Rw29_4 word29_4 word28_4 R_wl
Cwl_29_4 word29_4 gnd C_wl
Rw30_4 word30_4 word29_4 R_wl
Cwl_30_4 word30_4 gnd C_wl
Rw31_4 word31_4 word30_4 R_wl
Cwl_31_4 word31_4 gnd C_wl
Rw32_4 word32_4 word31_4 R_wl
Cwl_32_4 word32_4 gnd C_wl
Rw33_4 word33_4 word32_4 R_wl
Cwl_33_4 word33_4 gnd C_wl
Rw34_4 word34_4 word33_4 R_wl
Cwl_34_4 word34_4 gnd C_wl
Rw35_4 word35_4 word34_4 R_wl
Cwl_35_4 word35_4 gnd C_wl
Rw36_4 word36_4 word35_4 R_wl
Cwl_36_4 word36_4 gnd C_wl
Rw37_4 word37_4 word36_4 R_wl
Cwl_37_4 word37_4 gnd C_wl
Rw38_4 word38_4 word37_4 R_wl
Cwl_38_4 word38_4 gnd C_wl
Rw39_4 word39_4 word38_4 R_wl
Cwl_39_4 word39_4 gnd C_wl
Rw40_4 word40_4 word39_4 R_wl
Cwl_40_4 word40_4 gnd C_wl
Rw41_4 word41_4 word40_4 R_wl
Cwl_41_4 word41_4 gnd C_wl
Rw42_4 word42_4 word41_4 R_wl
Cwl_42_4 word42_4 gnd C_wl
Rw43_4 word43_4 word42_4 R_wl
Cwl_43_4 word43_4 gnd C_wl
Rw44_4 word44_4 word43_4 R_wl
Cwl_44_4 word44_4 gnd C_wl
Rw45_4 word45_4 word44_4 R_wl
Cwl_45_4 word45_4 gnd C_wl
Rw46_4 word46_4 word45_4 R_wl
Cwl_46_4 word46_4 gnd C_wl
Rw47_4 word47_4 word46_4 R_wl
Cwl_47_4 word47_4 gnd C_wl
Rw48_4 word48_4 word47_4 R_wl
Cwl_48_4 word48_4 gnd C_wl
Rw49_4 word49_4 word48_4 R_wl
Cwl_49_4 word49_4 gnd C_wl
Rw50_4 word50_4 word49_4 R_wl
Cwl_50_4 word50_4 gnd C_wl
Rw51_4 word51_4 word50_4 R_wl
Cwl_51_4 word51_4 gnd C_wl
Rw52_4 word52_4 word51_4 R_wl
Cwl_52_4 word52_4 gnd C_wl
Rw53_4 word53_4 word52_4 R_wl
Cwl_53_4 word53_4 gnd C_wl
Rw54_4 word54_4 word53_4 R_wl
Cwl_54_4 word54_4 gnd C_wl
Rw55_4 word55_4 word54_4 R_wl
Cwl_55_4 word55_4 gnd C_wl
Rw56_4 word56_4 word55_4 R_wl
Cwl_56_4 word56_4 gnd C_wl
Rw57_4 word57_4 word56_4 R_wl
Cwl_57_4 word57_4 gnd C_wl
Rw58_4 word58_4 word57_4 R_wl
Cwl_58_4 word58_4 gnd C_wl
Rw59_4 word59_4 word58_4 R_wl
Cwl_59_4 word59_4 gnd C_wl
Rw60_4 word60_4 word59_4 R_wl
Cwl_60_4 word60_4 gnd C_wl
Rw61_4 word61_4 word60_4 R_wl
Cwl_61_4 word61_4 gnd C_wl
Rw62_4 word62_4 word61_4 R_wl
Cwl_62_4 word62_4 gnd C_wl
Rw63_4 word63_4 word62_4 R_wl
Cwl_63_4 word63_4 gnd C_wl
Rw64_4 word64_4 word63_4 R_wl
Cwl_64_4 word64_4 gnd C_wl
Rw65_4 word65_4 word64_4 R_wl
Cwl_65_4 word65_4 gnd C_wl
Rw66_4 word66_4 word65_4 R_wl
Cwl_66_4 word66_4 gnd C_wl
Rw67_4 word67_4 word66_4 R_wl
Cwl_67_4 word67_4 gnd C_wl
Rw68_4 word68_4 word67_4 R_wl
Cwl_68_4 word68_4 gnd C_wl
Rw69_4 word69_4 word68_4 R_wl
Cwl_69_4 word69_4 gnd C_wl
Rw70_4 word70_4 word69_4 R_wl
Cwl_70_4 word70_4 gnd C_wl
Rw71_4 word71_4 word70_4 R_wl
Cwl_71_4 word71_4 gnd C_wl
Rw72_4 word72_4 word71_4 R_wl
Cwl_72_4 word72_4 gnd C_wl
Rw73_4 word73_4 word72_4 R_wl
Cwl_73_4 word73_4 gnd C_wl
Rw74_4 word74_4 word73_4 R_wl
Cwl_74_4 word74_4 gnd C_wl
Rw75_4 word75_4 word74_4 R_wl
Cwl_75_4 word75_4 gnd C_wl
Rw76_4 word76_4 word75_4 R_wl
Cwl_76_4 word76_4 gnd C_wl
Rw77_4 word77_4 word76_4 R_wl
Cwl_77_4 word77_4 gnd C_wl
Rw78_4 word78_4 word77_4 R_wl
Cwl_78_4 word78_4 gnd C_wl
Rw79_4 word79_4 word78_4 R_wl
Cwl_79_4 word79_4 gnd C_wl
Rw80_4 word80_4 word79_4 R_wl
Cwl_80_4 word80_4 gnd C_wl
Rw81_4 word81_4 word80_4 R_wl
Cwl_81_4 word81_4 gnd C_wl
Rw82_4 word82_4 word81_4 R_wl
Cwl_82_4 word82_4 gnd C_wl
Rw83_4 word83_4 word82_4 R_wl
Cwl_83_4 word83_4 gnd C_wl
Rw84_4 word84_4 word83_4 R_wl
Cwl_84_4 word84_4 gnd C_wl
Rw85_4 word85_4 word84_4 R_wl
Cwl_85_4 word85_4 gnd C_wl
Rw86_4 word86_4 word85_4 R_wl
Cwl_86_4 word86_4 gnd C_wl
Rw87_4 word87_4 word86_4 R_wl
Cwl_87_4 word87_4 gnd C_wl
Rw88_4 word88_4 word87_4 R_wl
Cwl_88_4 word88_4 gnd C_wl
Rw89_4 word89_4 word88_4 R_wl
Cwl_89_4 word89_4 gnd C_wl
Rw90_4 word90_4 word89_4 R_wl
Cwl_90_4 word90_4 gnd C_wl
Rw91_4 word91_4 word90_4 R_wl
Cwl_91_4 word91_4 gnd C_wl
Rw92_4 word92_4 word91_4 R_wl
Cwl_92_4 word92_4 gnd C_wl
Rw93_4 word93_4 word92_4 R_wl
Cwl_93_4 word93_4 gnd C_wl
Rw94_4 word94_4 word93_4 R_wl
Cwl_94_4 word94_4 gnd C_wl
Rw95_4 word95_4 word94_4 R_wl
Cwl_95_4 word95_4 gnd C_wl
Rw96_4 word96_4 word95_4 R_wl
Cwl_96_4 word96_4 gnd C_wl
Rw97_4 word97_4 word96_4 R_wl
Cwl_97_4 word97_4 gnd C_wl
Rw98_4 word98_4 word97_4 R_wl
Cwl_98_4 word98_4 gnd C_wl
Rw99_4 word99_4 word98_4 R_wl
Cwl_99_4 word99_4 gnd C_wl
Vwl_5 word_5 0 0
Rw0_5 word_5 word0_5 R_wl
Cwl_0_5 word0_5 gnd C_wl
Rw1_5 word1_5 word0_5 R_wl
Cwl_1_5 word1_5 gnd C_wl
Rw2_5 word2_5 word1_5 R_wl
Cwl_2_5 word2_5 gnd C_wl
Rw3_5 word3_5 word2_5 R_wl
Cwl_3_5 word3_5 gnd C_wl
Rw4_5 word4_5 word3_5 R_wl
Cwl_4_5 word4_5 gnd C_wl
Rw5_5 word5_5 word4_5 R_wl
Cwl_5_5 word5_5 gnd C_wl
Rw6_5 word6_5 word5_5 R_wl
Cwl_6_5 word6_5 gnd C_wl
Rw7_5 word7_5 word6_5 R_wl
Cwl_7_5 word7_5 gnd C_wl
Rw8_5 word8_5 word7_5 R_wl
Cwl_8_5 word8_5 gnd C_wl
Rw9_5 word9_5 word8_5 R_wl
Cwl_9_5 word9_5 gnd C_wl
Rw10_5 word10_5 word9_5 R_wl
Cwl_10_5 word10_5 gnd C_wl
Rw11_5 word11_5 word10_5 R_wl
Cwl_11_5 word11_5 gnd C_wl
Rw12_5 word12_5 word11_5 R_wl
Cwl_12_5 word12_5 gnd C_wl
Rw13_5 word13_5 word12_5 R_wl
Cwl_13_5 word13_5 gnd C_wl
Rw14_5 word14_5 word13_5 R_wl
Cwl_14_5 word14_5 gnd C_wl
Rw15_5 word15_5 word14_5 R_wl
Cwl_15_5 word15_5 gnd C_wl
Rw16_5 word16_5 word15_5 R_wl
Cwl_16_5 word16_5 gnd C_wl
Rw17_5 word17_5 word16_5 R_wl
Cwl_17_5 word17_5 gnd C_wl
Rw18_5 word18_5 word17_5 R_wl
Cwl_18_5 word18_5 gnd C_wl
Rw19_5 word19_5 word18_5 R_wl
Cwl_19_5 word19_5 gnd C_wl
Rw20_5 word20_5 word19_5 R_wl
Cwl_20_5 word20_5 gnd C_wl
Rw21_5 word21_5 word20_5 R_wl
Cwl_21_5 word21_5 gnd C_wl
Rw22_5 word22_5 word21_5 R_wl
Cwl_22_5 word22_5 gnd C_wl
Rw23_5 word23_5 word22_5 R_wl
Cwl_23_5 word23_5 gnd C_wl
Rw24_5 word24_5 word23_5 R_wl
Cwl_24_5 word24_5 gnd C_wl
Rw25_5 word25_5 word24_5 R_wl
Cwl_25_5 word25_5 gnd C_wl
Rw26_5 word26_5 word25_5 R_wl
Cwl_26_5 word26_5 gnd C_wl
Rw27_5 word27_5 word26_5 R_wl
Cwl_27_5 word27_5 gnd C_wl
Rw28_5 word28_5 word27_5 R_wl
Cwl_28_5 word28_5 gnd C_wl
Rw29_5 word29_5 word28_5 R_wl
Cwl_29_5 word29_5 gnd C_wl
Rw30_5 word30_5 word29_5 R_wl
Cwl_30_5 word30_5 gnd C_wl
Rw31_5 word31_5 word30_5 R_wl
Cwl_31_5 word31_5 gnd C_wl
Rw32_5 word32_5 word31_5 R_wl
Cwl_32_5 word32_5 gnd C_wl
Rw33_5 word33_5 word32_5 R_wl
Cwl_33_5 word33_5 gnd C_wl
Rw34_5 word34_5 word33_5 R_wl
Cwl_34_5 word34_5 gnd C_wl
Rw35_5 word35_5 word34_5 R_wl
Cwl_35_5 word35_5 gnd C_wl
Rw36_5 word36_5 word35_5 R_wl
Cwl_36_5 word36_5 gnd C_wl
Rw37_5 word37_5 word36_5 R_wl
Cwl_37_5 word37_5 gnd C_wl
Rw38_5 word38_5 word37_5 R_wl
Cwl_38_5 word38_5 gnd C_wl
Rw39_5 word39_5 word38_5 R_wl
Cwl_39_5 word39_5 gnd C_wl
Rw40_5 word40_5 word39_5 R_wl
Cwl_40_5 word40_5 gnd C_wl
Rw41_5 word41_5 word40_5 R_wl
Cwl_41_5 word41_5 gnd C_wl
Rw42_5 word42_5 word41_5 R_wl
Cwl_42_5 word42_5 gnd C_wl
Rw43_5 word43_5 word42_5 R_wl
Cwl_43_5 word43_5 gnd C_wl
Rw44_5 word44_5 word43_5 R_wl
Cwl_44_5 word44_5 gnd C_wl
Rw45_5 word45_5 word44_5 R_wl
Cwl_45_5 word45_5 gnd C_wl
Rw46_5 word46_5 word45_5 R_wl
Cwl_46_5 word46_5 gnd C_wl
Rw47_5 word47_5 word46_5 R_wl
Cwl_47_5 word47_5 gnd C_wl
Rw48_5 word48_5 word47_5 R_wl
Cwl_48_5 word48_5 gnd C_wl
Rw49_5 word49_5 word48_5 R_wl
Cwl_49_5 word49_5 gnd C_wl
Rw50_5 word50_5 word49_5 R_wl
Cwl_50_5 word50_5 gnd C_wl
Rw51_5 word51_5 word50_5 R_wl
Cwl_51_5 word51_5 gnd C_wl
Rw52_5 word52_5 word51_5 R_wl
Cwl_52_5 word52_5 gnd C_wl
Rw53_5 word53_5 word52_5 R_wl
Cwl_53_5 word53_5 gnd C_wl
Rw54_5 word54_5 word53_5 R_wl
Cwl_54_5 word54_5 gnd C_wl
Rw55_5 word55_5 word54_5 R_wl
Cwl_55_5 word55_5 gnd C_wl
Rw56_5 word56_5 word55_5 R_wl
Cwl_56_5 word56_5 gnd C_wl
Rw57_5 word57_5 word56_5 R_wl
Cwl_57_5 word57_5 gnd C_wl
Rw58_5 word58_5 word57_5 R_wl
Cwl_58_5 word58_5 gnd C_wl
Rw59_5 word59_5 word58_5 R_wl
Cwl_59_5 word59_5 gnd C_wl
Rw60_5 word60_5 word59_5 R_wl
Cwl_60_5 word60_5 gnd C_wl
Rw61_5 word61_5 word60_5 R_wl
Cwl_61_5 word61_5 gnd C_wl
Rw62_5 word62_5 word61_5 R_wl
Cwl_62_5 word62_5 gnd C_wl
Rw63_5 word63_5 word62_5 R_wl
Cwl_63_5 word63_5 gnd C_wl
Rw64_5 word64_5 word63_5 R_wl
Cwl_64_5 word64_5 gnd C_wl
Rw65_5 word65_5 word64_5 R_wl
Cwl_65_5 word65_5 gnd C_wl
Rw66_5 word66_5 word65_5 R_wl
Cwl_66_5 word66_5 gnd C_wl
Rw67_5 word67_5 word66_5 R_wl
Cwl_67_5 word67_5 gnd C_wl
Rw68_5 word68_5 word67_5 R_wl
Cwl_68_5 word68_5 gnd C_wl
Rw69_5 word69_5 word68_5 R_wl
Cwl_69_5 word69_5 gnd C_wl
Rw70_5 word70_5 word69_5 R_wl
Cwl_70_5 word70_5 gnd C_wl
Rw71_5 word71_5 word70_5 R_wl
Cwl_71_5 word71_5 gnd C_wl
Rw72_5 word72_5 word71_5 R_wl
Cwl_72_5 word72_5 gnd C_wl
Rw73_5 word73_5 word72_5 R_wl
Cwl_73_5 word73_5 gnd C_wl
Rw74_5 word74_5 word73_5 R_wl
Cwl_74_5 word74_5 gnd C_wl
Rw75_5 word75_5 word74_5 R_wl
Cwl_75_5 word75_5 gnd C_wl
Rw76_5 word76_5 word75_5 R_wl
Cwl_76_5 word76_5 gnd C_wl
Rw77_5 word77_5 word76_5 R_wl
Cwl_77_5 word77_5 gnd C_wl
Rw78_5 word78_5 word77_5 R_wl
Cwl_78_5 word78_5 gnd C_wl
Rw79_5 word79_5 word78_5 R_wl
Cwl_79_5 word79_5 gnd C_wl
Rw80_5 word80_5 word79_5 R_wl
Cwl_80_5 word80_5 gnd C_wl
Rw81_5 word81_5 word80_5 R_wl
Cwl_81_5 word81_5 gnd C_wl
Rw82_5 word82_5 word81_5 R_wl
Cwl_82_5 word82_5 gnd C_wl
Rw83_5 word83_5 word82_5 R_wl
Cwl_83_5 word83_5 gnd C_wl
Rw84_5 word84_5 word83_5 R_wl
Cwl_84_5 word84_5 gnd C_wl
Rw85_5 word85_5 word84_5 R_wl
Cwl_85_5 word85_5 gnd C_wl
Rw86_5 word86_5 word85_5 R_wl
Cwl_86_5 word86_5 gnd C_wl
Rw87_5 word87_5 word86_5 R_wl
Cwl_87_5 word87_5 gnd C_wl
Rw88_5 word88_5 word87_5 R_wl
Cwl_88_5 word88_5 gnd C_wl
Rw89_5 word89_5 word88_5 R_wl
Cwl_89_5 word89_5 gnd C_wl
Rw90_5 word90_5 word89_5 R_wl
Cwl_90_5 word90_5 gnd C_wl
Rw91_5 word91_5 word90_5 R_wl
Cwl_91_5 word91_5 gnd C_wl
Rw92_5 word92_5 word91_5 R_wl
Cwl_92_5 word92_5 gnd C_wl
Rw93_5 word93_5 word92_5 R_wl
Cwl_93_5 word93_5 gnd C_wl
Rw94_5 word94_5 word93_5 R_wl
Cwl_94_5 word94_5 gnd C_wl
Rw95_5 word95_5 word94_5 R_wl
Cwl_95_5 word95_5 gnd C_wl
Rw96_5 word96_5 word95_5 R_wl
Cwl_96_5 word96_5 gnd C_wl
Rw97_5 word97_5 word96_5 R_wl
Cwl_97_5 word97_5 gnd C_wl
Rw98_5 word98_5 word97_5 R_wl
Cwl_98_5 word98_5 gnd C_wl
Rw99_5 word99_5 word98_5 R_wl
Cwl_99_5 word99_5 gnd C_wl
Vwl_6 word_6 0 0
Rw0_6 word_6 word0_6 R_wl
Cwl_0_6 word0_6 gnd C_wl
Rw1_6 word1_6 word0_6 R_wl
Cwl_1_6 word1_6 gnd C_wl
Rw2_6 word2_6 word1_6 R_wl
Cwl_2_6 word2_6 gnd C_wl
Rw3_6 word3_6 word2_6 R_wl
Cwl_3_6 word3_6 gnd C_wl
Rw4_6 word4_6 word3_6 R_wl
Cwl_4_6 word4_6 gnd C_wl
Rw5_6 word5_6 word4_6 R_wl
Cwl_5_6 word5_6 gnd C_wl
Rw6_6 word6_6 word5_6 R_wl
Cwl_6_6 word6_6 gnd C_wl
Rw7_6 word7_6 word6_6 R_wl
Cwl_7_6 word7_6 gnd C_wl
Rw8_6 word8_6 word7_6 R_wl
Cwl_8_6 word8_6 gnd C_wl
Rw9_6 word9_6 word8_6 R_wl
Cwl_9_6 word9_6 gnd C_wl
Rw10_6 word10_6 word9_6 R_wl
Cwl_10_6 word10_6 gnd C_wl
Rw11_6 word11_6 word10_6 R_wl
Cwl_11_6 word11_6 gnd C_wl
Rw12_6 word12_6 word11_6 R_wl
Cwl_12_6 word12_6 gnd C_wl
Rw13_6 word13_6 word12_6 R_wl
Cwl_13_6 word13_6 gnd C_wl
Rw14_6 word14_6 word13_6 R_wl
Cwl_14_6 word14_6 gnd C_wl
Rw15_6 word15_6 word14_6 R_wl
Cwl_15_6 word15_6 gnd C_wl
Rw16_6 word16_6 word15_6 R_wl
Cwl_16_6 word16_6 gnd C_wl
Rw17_6 word17_6 word16_6 R_wl
Cwl_17_6 word17_6 gnd C_wl
Rw18_6 word18_6 word17_6 R_wl
Cwl_18_6 word18_6 gnd C_wl
Rw19_6 word19_6 word18_6 R_wl
Cwl_19_6 word19_6 gnd C_wl
Rw20_6 word20_6 word19_6 R_wl
Cwl_20_6 word20_6 gnd C_wl
Rw21_6 word21_6 word20_6 R_wl
Cwl_21_6 word21_6 gnd C_wl
Rw22_6 word22_6 word21_6 R_wl
Cwl_22_6 word22_6 gnd C_wl
Rw23_6 word23_6 word22_6 R_wl
Cwl_23_6 word23_6 gnd C_wl
Rw24_6 word24_6 word23_6 R_wl
Cwl_24_6 word24_6 gnd C_wl
Rw25_6 word25_6 word24_6 R_wl
Cwl_25_6 word25_6 gnd C_wl
Rw26_6 word26_6 word25_6 R_wl
Cwl_26_6 word26_6 gnd C_wl
Rw27_6 word27_6 word26_6 R_wl
Cwl_27_6 word27_6 gnd C_wl
Rw28_6 word28_6 word27_6 R_wl
Cwl_28_6 word28_6 gnd C_wl
Rw29_6 word29_6 word28_6 R_wl
Cwl_29_6 word29_6 gnd C_wl
Rw30_6 word30_6 word29_6 R_wl
Cwl_30_6 word30_6 gnd C_wl
Rw31_6 word31_6 word30_6 R_wl
Cwl_31_6 word31_6 gnd C_wl
Rw32_6 word32_6 word31_6 R_wl
Cwl_32_6 word32_6 gnd C_wl
Rw33_6 word33_6 word32_6 R_wl
Cwl_33_6 word33_6 gnd C_wl
Rw34_6 word34_6 word33_6 R_wl
Cwl_34_6 word34_6 gnd C_wl
Rw35_6 word35_6 word34_6 R_wl
Cwl_35_6 word35_6 gnd C_wl
Rw36_6 word36_6 word35_6 R_wl
Cwl_36_6 word36_6 gnd C_wl
Rw37_6 word37_6 word36_6 R_wl
Cwl_37_6 word37_6 gnd C_wl
Rw38_6 word38_6 word37_6 R_wl
Cwl_38_6 word38_6 gnd C_wl
Rw39_6 word39_6 word38_6 R_wl
Cwl_39_6 word39_6 gnd C_wl
Rw40_6 word40_6 word39_6 R_wl
Cwl_40_6 word40_6 gnd C_wl
Rw41_6 word41_6 word40_6 R_wl
Cwl_41_6 word41_6 gnd C_wl
Rw42_6 word42_6 word41_6 R_wl
Cwl_42_6 word42_6 gnd C_wl
Rw43_6 word43_6 word42_6 R_wl
Cwl_43_6 word43_6 gnd C_wl
Rw44_6 word44_6 word43_6 R_wl
Cwl_44_6 word44_6 gnd C_wl
Rw45_6 word45_6 word44_6 R_wl
Cwl_45_6 word45_6 gnd C_wl
Rw46_6 word46_6 word45_6 R_wl
Cwl_46_6 word46_6 gnd C_wl
Rw47_6 word47_6 word46_6 R_wl
Cwl_47_6 word47_6 gnd C_wl
Rw48_6 word48_6 word47_6 R_wl
Cwl_48_6 word48_6 gnd C_wl
Rw49_6 word49_6 word48_6 R_wl
Cwl_49_6 word49_6 gnd C_wl
Rw50_6 word50_6 word49_6 R_wl
Cwl_50_6 word50_6 gnd C_wl
Rw51_6 word51_6 word50_6 R_wl
Cwl_51_6 word51_6 gnd C_wl
Rw52_6 word52_6 word51_6 R_wl
Cwl_52_6 word52_6 gnd C_wl
Rw53_6 word53_6 word52_6 R_wl
Cwl_53_6 word53_6 gnd C_wl
Rw54_6 word54_6 word53_6 R_wl
Cwl_54_6 word54_6 gnd C_wl
Rw55_6 word55_6 word54_6 R_wl
Cwl_55_6 word55_6 gnd C_wl
Rw56_6 word56_6 word55_6 R_wl
Cwl_56_6 word56_6 gnd C_wl
Rw57_6 word57_6 word56_6 R_wl
Cwl_57_6 word57_6 gnd C_wl
Rw58_6 word58_6 word57_6 R_wl
Cwl_58_6 word58_6 gnd C_wl
Rw59_6 word59_6 word58_6 R_wl
Cwl_59_6 word59_6 gnd C_wl
Rw60_6 word60_6 word59_6 R_wl
Cwl_60_6 word60_6 gnd C_wl
Rw61_6 word61_6 word60_6 R_wl
Cwl_61_6 word61_6 gnd C_wl
Rw62_6 word62_6 word61_6 R_wl
Cwl_62_6 word62_6 gnd C_wl
Rw63_6 word63_6 word62_6 R_wl
Cwl_63_6 word63_6 gnd C_wl
Rw64_6 word64_6 word63_6 R_wl
Cwl_64_6 word64_6 gnd C_wl
Rw65_6 word65_6 word64_6 R_wl
Cwl_65_6 word65_6 gnd C_wl
Rw66_6 word66_6 word65_6 R_wl
Cwl_66_6 word66_6 gnd C_wl
Rw67_6 word67_6 word66_6 R_wl
Cwl_67_6 word67_6 gnd C_wl
Rw68_6 word68_6 word67_6 R_wl
Cwl_68_6 word68_6 gnd C_wl
Rw69_6 word69_6 word68_6 R_wl
Cwl_69_6 word69_6 gnd C_wl
Rw70_6 word70_6 word69_6 R_wl
Cwl_70_6 word70_6 gnd C_wl
Rw71_6 word71_6 word70_6 R_wl
Cwl_71_6 word71_6 gnd C_wl
Rw72_6 word72_6 word71_6 R_wl
Cwl_72_6 word72_6 gnd C_wl
Rw73_6 word73_6 word72_6 R_wl
Cwl_73_6 word73_6 gnd C_wl
Rw74_6 word74_6 word73_6 R_wl
Cwl_74_6 word74_6 gnd C_wl
Rw75_6 word75_6 word74_6 R_wl
Cwl_75_6 word75_6 gnd C_wl
Rw76_6 word76_6 word75_6 R_wl
Cwl_76_6 word76_6 gnd C_wl
Rw77_6 word77_6 word76_6 R_wl
Cwl_77_6 word77_6 gnd C_wl
Rw78_6 word78_6 word77_6 R_wl
Cwl_78_6 word78_6 gnd C_wl
Rw79_6 word79_6 word78_6 R_wl
Cwl_79_6 word79_6 gnd C_wl
Rw80_6 word80_6 word79_6 R_wl
Cwl_80_6 word80_6 gnd C_wl
Rw81_6 word81_6 word80_6 R_wl
Cwl_81_6 word81_6 gnd C_wl
Rw82_6 word82_6 word81_6 R_wl
Cwl_82_6 word82_6 gnd C_wl
Rw83_6 word83_6 word82_6 R_wl
Cwl_83_6 word83_6 gnd C_wl
Rw84_6 word84_6 word83_6 R_wl
Cwl_84_6 word84_6 gnd C_wl
Rw85_6 word85_6 word84_6 R_wl
Cwl_85_6 word85_6 gnd C_wl
Rw86_6 word86_6 word85_6 R_wl
Cwl_86_6 word86_6 gnd C_wl
Rw87_6 word87_6 word86_6 R_wl
Cwl_87_6 word87_6 gnd C_wl
Rw88_6 word88_6 word87_6 R_wl
Cwl_88_6 word88_6 gnd C_wl
Rw89_6 word89_6 word88_6 R_wl
Cwl_89_6 word89_6 gnd C_wl
Rw90_6 word90_6 word89_6 R_wl
Cwl_90_6 word90_6 gnd C_wl
Rw91_6 word91_6 word90_6 R_wl
Cwl_91_6 word91_6 gnd C_wl
Rw92_6 word92_6 word91_6 R_wl
Cwl_92_6 word92_6 gnd C_wl
Rw93_6 word93_6 word92_6 R_wl
Cwl_93_6 word93_6 gnd C_wl
Rw94_6 word94_6 word93_6 R_wl
Cwl_94_6 word94_6 gnd C_wl
Rw95_6 word95_6 word94_6 R_wl
Cwl_95_6 word95_6 gnd C_wl
Rw96_6 word96_6 word95_6 R_wl
Cwl_96_6 word96_6 gnd C_wl
Rw97_6 word97_6 word96_6 R_wl
Cwl_97_6 word97_6 gnd C_wl
Rw98_6 word98_6 word97_6 R_wl
Cwl_98_6 word98_6 gnd C_wl
Rw99_6 word99_6 word98_6 R_wl
Cwl_99_6 word99_6 gnd C_wl
Vwl_7 word_7 0 0
Rw0_7 word_7 word0_7 R_wl
Cwl_0_7 word0_7 gnd C_wl
Rw1_7 word1_7 word0_7 R_wl
Cwl_1_7 word1_7 gnd C_wl
Rw2_7 word2_7 word1_7 R_wl
Cwl_2_7 word2_7 gnd C_wl
Rw3_7 word3_7 word2_7 R_wl
Cwl_3_7 word3_7 gnd C_wl
Rw4_7 word4_7 word3_7 R_wl
Cwl_4_7 word4_7 gnd C_wl
Rw5_7 word5_7 word4_7 R_wl
Cwl_5_7 word5_7 gnd C_wl
Rw6_7 word6_7 word5_7 R_wl
Cwl_6_7 word6_7 gnd C_wl
Rw7_7 word7_7 word6_7 R_wl
Cwl_7_7 word7_7 gnd C_wl
Rw8_7 word8_7 word7_7 R_wl
Cwl_8_7 word8_7 gnd C_wl
Rw9_7 word9_7 word8_7 R_wl
Cwl_9_7 word9_7 gnd C_wl
Rw10_7 word10_7 word9_7 R_wl
Cwl_10_7 word10_7 gnd C_wl
Rw11_7 word11_7 word10_7 R_wl
Cwl_11_7 word11_7 gnd C_wl
Rw12_7 word12_7 word11_7 R_wl
Cwl_12_7 word12_7 gnd C_wl
Rw13_7 word13_7 word12_7 R_wl
Cwl_13_7 word13_7 gnd C_wl
Rw14_7 word14_7 word13_7 R_wl
Cwl_14_7 word14_7 gnd C_wl
Rw15_7 word15_7 word14_7 R_wl
Cwl_15_7 word15_7 gnd C_wl
Rw16_7 word16_7 word15_7 R_wl
Cwl_16_7 word16_7 gnd C_wl
Rw17_7 word17_7 word16_7 R_wl
Cwl_17_7 word17_7 gnd C_wl
Rw18_7 word18_7 word17_7 R_wl
Cwl_18_7 word18_7 gnd C_wl
Rw19_7 word19_7 word18_7 R_wl
Cwl_19_7 word19_7 gnd C_wl
Rw20_7 word20_7 word19_7 R_wl
Cwl_20_7 word20_7 gnd C_wl
Rw21_7 word21_7 word20_7 R_wl
Cwl_21_7 word21_7 gnd C_wl
Rw22_7 word22_7 word21_7 R_wl
Cwl_22_7 word22_7 gnd C_wl
Rw23_7 word23_7 word22_7 R_wl
Cwl_23_7 word23_7 gnd C_wl
Rw24_7 word24_7 word23_7 R_wl
Cwl_24_7 word24_7 gnd C_wl
Rw25_7 word25_7 word24_7 R_wl
Cwl_25_7 word25_7 gnd C_wl
Rw26_7 word26_7 word25_7 R_wl
Cwl_26_7 word26_7 gnd C_wl
Rw27_7 word27_7 word26_7 R_wl
Cwl_27_7 word27_7 gnd C_wl
Rw28_7 word28_7 word27_7 R_wl
Cwl_28_7 word28_7 gnd C_wl
Rw29_7 word29_7 word28_7 R_wl
Cwl_29_7 word29_7 gnd C_wl
Rw30_7 word30_7 word29_7 R_wl
Cwl_30_7 word30_7 gnd C_wl
Rw31_7 word31_7 word30_7 R_wl
Cwl_31_7 word31_7 gnd C_wl
Rw32_7 word32_7 word31_7 R_wl
Cwl_32_7 word32_7 gnd C_wl
Rw33_7 word33_7 word32_7 R_wl
Cwl_33_7 word33_7 gnd C_wl
Rw34_7 word34_7 word33_7 R_wl
Cwl_34_7 word34_7 gnd C_wl
Rw35_7 word35_7 word34_7 R_wl
Cwl_35_7 word35_7 gnd C_wl
Rw36_7 word36_7 word35_7 R_wl
Cwl_36_7 word36_7 gnd C_wl
Rw37_7 word37_7 word36_7 R_wl
Cwl_37_7 word37_7 gnd C_wl
Rw38_7 word38_7 word37_7 R_wl
Cwl_38_7 word38_7 gnd C_wl
Rw39_7 word39_7 word38_7 R_wl
Cwl_39_7 word39_7 gnd C_wl
Rw40_7 word40_7 word39_7 R_wl
Cwl_40_7 word40_7 gnd C_wl
Rw41_7 word41_7 word40_7 R_wl
Cwl_41_7 word41_7 gnd C_wl
Rw42_7 word42_7 word41_7 R_wl
Cwl_42_7 word42_7 gnd C_wl
Rw43_7 word43_7 word42_7 R_wl
Cwl_43_7 word43_7 gnd C_wl
Rw44_7 word44_7 word43_7 R_wl
Cwl_44_7 word44_7 gnd C_wl
Rw45_7 word45_7 word44_7 R_wl
Cwl_45_7 word45_7 gnd C_wl
Rw46_7 word46_7 word45_7 R_wl
Cwl_46_7 word46_7 gnd C_wl
Rw47_7 word47_7 word46_7 R_wl
Cwl_47_7 word47_7 gnd C_wl
Rw48_7 word48_7 word47_7 R_wl
Cwl_48_7 word48_7 gnd C_wl
Rw49_7 word49_7 word48_7 R_wl
Cwl_49_7 word49_7 gnd C_wl
Rw50_7 word50_7 word49_7 R_wl
Cwl_50_7 word50_7 gnd C_wl
Rw51_7 word51_7 word50_7 R_wl
Cwl_51_7 word51_7 gnd C_wl
Rw52_7 word52_7 word51_7 R_wl
Cwl_52_7 word52_7 gnd C_wl
Rw53_7 word53_7 word52_7 R_wl
Cwl_53_7 word53_7 gnd C_wl
Rw54_7 word54_7 word53_7 R_wl
Cwl_54_7 word54_7 gnd C_wl
Rw55_7 word55_7 word54_7 R_wl
Cwl_55_7 word55_7 gnd C_wl
Rw56_7 word56_7 word55_7 R_wl
Cwl_56_7 word56_7 gnd C_wl
Rw57_7 word57_7 word56_7 R_wl
Cwl_57_7 word57_7 gnd C_wl
Rw58_7 word58_7 word57_7 R_wl
Cwl_58_7 word58_7 gnd C_wl
Rw59_7 word59_7 word58_7 R_wl
Cwl_59_7 word59_7 gnd C_wl
Rw60_7 word60_7 word59_7 R_wl
Cwl_60_7 word60_7 gnd C_wl
Rw61_7 word61_7 word60_7 R_wl
Cwl_61_7 word61_7 gnd C_wl
Rw62_7 word62_7 word61_7 R_wl
Cwl_62_7 word62_7 gnd C_wl
Rw63_7 word63_7 word62_7 R_wl
Cwl_63_7 word63_7 gnd C_wl
Rw64_7 word64_7 word63_7 R_wl
Cwl_64_7 word64_7 gnd C_wl
Rw65_7 word65_7 word64_7 R_wl
Cwl_65_7 word65_7 gnd C_wl
Rw66_7 word66_7 word65_7 R_wl
Cwl_66_7 word66_7 gnd C_wl
Rw67_7 word67_7 word66_7 R_wl
Cwl_67_7 word67_7 gnd C_wl
Rw68_7 word68_7 word67_7 R_wl
Cwl_68_7 word68_7 gnd C_wl
Rw69_7 word69_7 word68_7 R_wl
Cwl_69_7 word69_7 gnd C_wl
Rw70_7 word70_7 word69_7 R_wl
Cwl_70_7 word70_7 gnd C_wl
Rw71_7 word71_7 word70_7 R_wl
Cwl_71_7 word71_7 gnd C_wl
Rw72_7 word72_7 word71_7 R_wl
Cwl_72_7 word72_7 gnd C_wl
Rw73_7 word73_7 word72_7 R_wl
Cwl_73_7 word73_7 gnd C_wl
Rw74_7 word74_7 word73_7 R_wl
Cwl_74_7 word74_7 gnd C_wl
Rw75_7 word75_7 word74_7 R_wl
Cwl_75_7 word75_7 gnd C_wl
Rw76_7 word76_7 word75_7 R_wl
Cwl_76_7 word76_7 gnd C_wl
Rw77_7 word77_7 word76_7 R_wl
Cwl_77_7 word77_7 gnd C_wl
Rw78_7 word78_7 word77_7 R_wl
Cwl_78_7 word78_7 gnd C_wl
Rw79_7 word79_7 word78_7 R_wl
Cwl_79_7 word79_7 gnd C_wl
Rw80_7 word80_7 word79_7 R_wl
Cwl_80_7 word80_7 gnd C_wl
Rw81_7 word81_7 word80_7 R_wl
Cwl_81_7 word81_7 gnd C_wl
Rw82_7 word82_7 word81_7 R_wl
Cwl_82_7 word82_7 gnd C_wl
Rw83_7 word83_7 word82_7 R_wl
Cwl_83_7 word83_7 gnd C_wl
Rw84_7 word84_7 word83_7 R_wl
Cwl_84_7 word84_7 gnd C_wl
Rw85_7 word85_7 word84_7 R_wl
Cwl_85_7 word85_7 gnd C_wl
Rw86_7 word86_7 word85_7 R_wl
Cwl_86_7 word86_7 gnd C_wl
Rw87_7 word87_7 word86_7 R_wl
Cwl_87_7 word87_7 gnd C_wl
Rw88_7 word88_7 word87_7 R_wl
Cwl_88_7 word88_7 gnd C_wl
Rw89_7 word89_7 word88_7 R_wl
Cwl_89_7 word89_7 gnd C_wl
Rw90_7 word90_7 word89_7 R_wl
Cwl_90_7 word90_7 gnd C_wl
Rw91_7 word91_7 word90_7 R_wl
Cwl_91_7 word91_7 gnd C_wl
Rw92_7 word92_7 word91_7 R_wl
Cwl_92_7 word92_7 gnd C_wl
Rw93_7 word93_7 word92_7 R_wl
Cwl_93_7 word93_7 gnd C_wl
Rw94_7 word94_7 word93_7 R_wl
Cwl_94_7 word94_7 gnd C_wl
Rw95_7 word95_7 word94_7 R_wl
Cwl_95_7 word95_7 gnd C_wl
Rw96_7 word96_7 word95_7 R_wl
Cwl_96_7 word96_7 gnd C_wl
Rw97_7 word97_7 word96_7 R_wl
Cwl_97_7 word97_7 gnd C_wl
Rw98_7 word98_7 word97_7 R_wl
Cwl_98_7 word98_7 gnd C_wl
Rw99_7 word99_7 word98_7 R_wl
Cwl_99_7 word99_7 gnd C_wl
Vwl_8 word_8 0 0
Rw0_8 word_8 word0_8 R_wl
Cwl_0_8 word0_8 gnd C_wl
Rw1_8 word1_8 word0_8 R_wl
Cwl_1_8 word1_8 gnd C_wl
Rw2_8 word2_8 word1_8 R_wl
Cwl_2_8 word2_8 gnd C_wl
Rw3_8 word3_8 word2_8 R_wl
Cwl_3_8 word3_8 gnd C_wl
Rw4_8 word4_8 word3_8 R_wl
Cwl_4_8 word4_8 gnd C_wl
Rw5_8 word5_8 word4_8 R_wl
Cwl_5_8 word5_8 gnd C_wl
Rw6_8 word6_8 word5_8 R_wl
Cwl_6_8 word6_8 gnd C_wl
Rw7_8 word7_8 word6_8 R_wl
Cwl_7_8 word7_8 gnd C_wl
Rw8_8 word8_8 word7_8 R_wl
Cwl_8_8 word8_8 gnd C_wl
Rw9_8 word9_8 word8_8 R_wl
Cwl_9_8 word9_8 gnd C_wl
Rw10_8 word10_8 word9_8 R_wl
Cwl_10_8 word10_8 gnd C_wl
Rw11_8 word11_8 word10_8 R_wl
Cwl_11_8 word11_8 gnd C_wl
Rw12_8 word12_8 word11_8 R_wl
Cwl_12_8 word12_8 gnd C_wl
Rw13_8 word13_8 word12_8 R_wl
Cwl_13_8 word13_8 gnd C_wl
Rw14_8 word14_8 word13_8 R_wl
Cwl_14_8 word14_8 gnd C_wl
Rw15_8 word15_8 word14_8 R_wl
Cwl_15_8 word15_8 gnd C_wl
Rw16_8 word16_8 word15_8 R_wl
Cwl_16_8 word16_8 gnd C_wl
Rw17_8 word17_8 word16_8 R_wl
Cwl_17_8 word17_8 gnd C_wl
Rw18_8 word18_8 word17_8 R_wl
Cwl_18_8 word18_8 gnd C_wl
Rw19_8 word19_8 word18_8 R_wl
Cwl_19_8 word19_8 gnd C_wl
Rw20_8 word20_8 word19_8 R_wl
Cwl_20_8 word20_8 gnd C_wl
Rw21_8 word21_8 word20_8 R_wl
Cwl_21_8 word21_8 gnd C_wl
Rw22_8 word22_8 word21_8 R_wl
Cwl_22_8 word22_8 gnd C_wl
Rw23_8 word23_8 word22_8 R_wl
Cwl_23_8 word23_8 gnd C_wl
Rw24_8 word24_8 word23_8 R_wl
Cwl_24_8 word24_8 gnd C_wl
Rw25_8 word25_8 word24_8 R_wl
Cwl_25_8 word25_8 gnd C_wl
Rw26_8 word26_8 word25_8 R_wl
Cwl_26_8 word26_8 gnd C_wl
Rw27_8 word27_8 word26_8 R_wl
Cwl_27_8 word27_8 gnd C_wl
Rw28_8 word28_8 word27_8 R_wl
Cwl_28_8 word28_8 gnd C_wl
Rw29_8 word29_8 word28_8 R_wl
Cwl_29_8 word29_8 gnd C_wl
Rw30_8 word30_8 word29_8 R_wl
Cwl_30_8 word30_8 gnd C_wl
Rw31_8 word31_8 word30_8 R_wl
Cwl_31_8 word31_8 gnd C_wl
Rw32_8 word32_8 word31_8 R_wl
Cwl_32_8 word32_8 gnd C_wl
Rw33_8 word33_8 word32_8 R_wl
Cwl_33_8 word33_8 gnd C_wl
Rw34_8 word34_8 word33_8 R_wl
Cwl_34_8 word34_8 gnd C_wl
Rw35_8 word35_8 word34_8 R_wl
Cwl_35_8 word35_8 gnd C_wl
Rw36_8 word36_8 word35_8 R_wl
Cwl_36_8 word36_8 gnd C_wl
Rw37_8 word37_8 word36_8 R_wl
Cwl_37_8 word37_8 gnd C_wl
Rw38_8 word38_8 word37_8 R_wl
Cwl_38_8 word38_8 gnd C_wl
Rw39_8 word39_8 word38_8 R_wl
Cwl_39_8 word39_8 gnd C_wl
Rw40_8 word40_8 word39_8 R_wl
Cwl_40_8 word40_8 gnd C_wl
Rw41_8 word41_8 word40_8 R_wl
Cwl_41_8 word41_8 gnd C_wl
Rw42_8 word42_8 word41_8 R_wl
Cwl_42_8 word42_8 gnd C_wl
Rw43_8 word43_8 word42_8 R_wl
Cwl_43_8 word43_8 gnd C_wl
Rw44_8 word44_8 word43_8 R_wl
Cwl_44_8 word44_8 gnd C_wl
Rw45_8 word45_8 word44_8 R_wl
Cwl_45_8 word45_8 gnd C_wl
Rw46_8 word46_8 word45_8 R_wl
Cwl_46_8 word46_8 gnd C_wl
Rw47_8 word47_8 word46_8 R_wl
Cwl_47_8 word47_8 gnd C_wl
Rw48_8 word48_8 word47_8 R_wl
Cwl_48_8 word48_8 gnd C_wl
Rw49_8 word49_8 word48_8 R_wl
Cwl_49_8 word49_8 gnd C_wl
Rw50_8 word50_8 word49_8 R_wl
Cwl_50_8 word50_8 gnd C_wl
Rw51_8 word51_8 word50_8 R_wl
Cwl_51_8 word51_8 gnd C_wl
Rw52_8 word52_8 word51_8 R_wl
Cwl_52_8 word52_8 gnd C_wl
Rw53_8 word53_8 word52_8 R_wl
Cwl_53_8 word53_8 gnd C_wl
Rw54_8 word54_8 word53_8 R_wl
Cwl_54_8 word54_8 gnd C_wl
Rw55_8 word55_8 word54_8 R_wl
Cwl_55_8 word55_8 gnd C_wl
Rw56_8 word56_8 word55_8 R_wl
Cwl_56_8 word56_8 gnd C_wl
Rw57_8 word57_8 word56_8 R_wl
Cwl_57_8 word57_8 gnd C_wl
Rw58_8 word58_8 word57_8 R_wl
Cwl_58_8 word58_8 gnd C_wl
Rw59_8 word59_8 word58_8 R_wl
Cwl_59_8 word59_8 gnd C_wl
Rw60_8 word60_8 word59_8 R_wl
Cwl_60_8 word60_8 gnd C_wl
Rw61_8 word61_8 word60_8 R_wl
Cwl_61_8 word61_8 gnd C_wl
Rw62_8 word62_8 word61_8 R_wl
Cwl_62_8 word62_8 gnd C_wl
Rw63_8 word63_8 word62_8 R_wl
Cwl_63_8 word63_8 gnd C_wl
Rw64_8 word64_8 word63_8 R_wl
Cwl_64_8 word64_8 gnd C_wl
Rw65_8 word65_8 word64_8 R_wl
Cwl_65_8 word65_8 gnd C_wl
Rw66_8 word66_8 word65_8 R_wl
Cwl_66_8 word66_8 gnd C_wl
Rw67_8 word67_8 word66_8 R_wl
Cwl_67_8 word67_8 gnd C_wl
Rw68_8 word68_8 word67_8 R_wl
Cwl_68_8 word68_8 gnd C_wl
Rw69_8 word69_8 word68_8 R_wl
Cwl_69_8 word69_8 gnd C_wl
Rw70_8 word70_8 word69_8 R_wl
Cwl_70_8 word70_8 gnd C_wl
Rw71_8 word71_8 word70_8 R_wl
Cwl_71_8 word71_8 gnd C_wl
Rw72_8 word72_8 word71_8 R_wl
Cwl_72_8 word72_8 gnd C_wl
Rw73_8 word73_8 word72_8 R_wl
Cwl_73_8 word73_8 gnd C_wl
Rw74_8 word74_8 word73_8 R_wl
Cwl_74_8 word74_8 gnd C_wl
Rw75_8 word75_8 word74_8 R_wl
Cwl_75_8 word75_8 gnd C_wl
Rw76_8 word76_8 word75_8 R_wl
Cwl_76_8 word76_8 gnd C_wl
Rw77_8 word77_8 word76_8 R_wl
Cwl_77_8 word77_8 gnd C_wl
Rw78_8 word78_8 word77_8 R_wl
Cwl_78_8 word78_8 gnd C_wl
Rw79_8 word79_8 word78_8 R_wl
Cwl_79_8 word79_8 gnd C_wl
Rw80_8 word80_8 word79_8 R_wl
Cwl_80_8 word80_8 gnd C_wl
Rw81_8 word81_8 word80_8 R_wl
Cwl_81_8 word81_8 gnd C_wl
Rw82_8 word82_8 word81_8 R_wl
Cwl_82_8 word82_8 gnd C_wl
Rw83_8 word83_8 word82_8 R_wl
Cwl_83_8 word83_8 gnd C_wl
Rw84_8 word84_8 word83_8 R_wl
Cwl_84_8 word84_8 gnd C_wl
Rw85_8 word85_8 word84_8 R_wl
Cwl_85_8 word85_8 gnd C_wl
Rw86_8 word86_8 word85_8 R_wl
Cwl_86_8 word86_8 gnd C_wl
Rw87_8 word87_8 word86_8 R_wl
Cwl_87_8 word87_8 gnd C_wl
Rw88_8 word88_8 word87_8 R_wl
Cwl_88_8 word88_8 gnd C_wl
Rw89_8 word89_8 word88_8 R_wl
Cwl_89_8 word89_8 gnd C_wl
Rw90_8 word90_8 word89_8 R_wl
Cwl_90_8 word90_8 gnd C_wl
Rw91_8 word91_8 word90_8 R_wl
Cwl_91_8 word91_8 gnd C_wl
Rw92_8 word92_8 word91_8 R_wl
Cwl_92_8 word92_8 gnd C_wl
Rw93_8 word93_8 word92_8 R_wl
Cwl_93_8 word93_8 gnd C_wl
Rw94_8 word94_8 word93_8 R_wl
Cwl_94_8 word94_8 gnd C_wl
Rw95_8 word95_8 word94_8 R_wl
Cwl_95_8 word95_8 gnd C_wl
Rw96_8 word96_8 word95_8 R_wl
Cwl_96_8 word96_8 gnd C_wl
Rw97_8 word97_8 word96_8 R_wl
Cwl_97_8 word97_8 gnd C_wl
Rw98_8 word98_8 word97_8 R_wl
Cwl_98_8 word98_8 gnd C_wl
Rw99_8 word99_8 word98_8 R_wl
Cwl_99_8 word99_8 gnd C_wl
Vwl_9 word_9 0 0
Rw0_9 word_9 word0_9 R_wl
Cwl_0_9 word0_9 gnd C_wl
Rw1_9 word1_9 word0_9 R_wl
Cwl_1_9 word1_9 gnd C_wl
Rw2_9 word2_9 word1_9 R_wl
Cwl_2_9 word2_9 gnd C_wl
Rw3_9 word3_9 word2_9 R_wl
Cwl_3_9 word3_9 gnd C_wl
Rw4_9 word4_9 word3_9 R_wl
Cwl_4_9 word4_9 gnd C_wl
Rw5_9 word5_9 word4_9 R_wl
Cwl_5_9 word5_9 gnd C_wl
Rw6_9 word6_9 word5_9 R_wl
Cwl_6_9 word6_9 gnd C_wl
Rw7_9 word7_9 word6_9 R_wl
Cwl_7_9 word7_9 gnd C_wl
Rw8_9 word8_9 word7_9 R_wl
Cwl_8_9 word8_9 gnd C_wl
Rw9_9 word9_9 word8_9 R_wl
Cwl_9_9 word9_9 gnd C_wl
Rw10_9 word10_9 word9_9 R_wl
Cwl_10_9 word10_9 gnd C_wl
Rw11_9 word11_9 word10_9 R_wl
Cwl_11_9 word11_9 gnd C_wl
Rw12_9 word12_9 word11_9 R_wl
Cwl_12_9 word12_9 gnd C_wl
Rw13_9 word13_9 word12_9 R_wl
Cwl_13_9 word13_9 gnd C_wl
Rw14_9 word14_9 word13_9 R_wl
Cwl_14_9 word14_9 gnd C_wl
Rw15_9 word15_9 word14_9 R_wl
Cwl_15_9 word15_9 gnd C_wl
Rw16_9 word16_9 word15_9 R_wl
Cwl_16_9 word16_9 gnd C_wl
Rw17_9 word17_9 word16_9 R_wl
Cwl_17_9 word17_9 gnd C_wl
Rw18_9 word18_9 word17_9 R_wl
Cwl_18_9 word18_9 gnd C_wl
Rw19_9 word19_9 word18_9 R_wl
Cwl_19_9 word19_9 gnd C_wl
Rw20_9 word20_9 word19_9 R_wl
Cwl_20_9 word20_9 gnd C_wl
Rw21_9 word21_9 word20_9 R_wl
Cwl_21_9 word21_9 gnd C_wl
Rw22_9 word22_9 word21_9 R_wl
Cwl_22_9 word22_9 gnd C_wl
Rw23_9 word23_9 word22_9 R_wl
Cwl_23_9 word23_9 gnd C_wl
Rw24_9 word24_9 word23_9 R_wl
Cwl_24_9 word24_9 gnd C_wl
Rw25_9 word25_9 word24_9 R_wl
Cwl_25_9 word25_9 gnd C_wl
Rw26_9 word26_9 word25_9 R_wl
Cwl_26_9 word26_9 gnd C_wl
Rw27_9 word27_9 word26_9 R_wl
Cwl_27_9 word27_9 gnd C_wl
Rw28_9 word28_9 word27_9 R_wl
Cwl_28_9 word28_9 gnd C_wl
Rw29_9 word29_9 word28_9 R_wl
Cwl_29_9 word29_9 gnd C_wl
Rw30_9 word30_9 word29_9 R_wl
Cwl_30_9 word30_9 gnd C_wl
Rw31_9 word31_9 word30_9 R_wl
Cwl_31_9 word31_9 gnd C_wl
Rw32_9 word32_9 word31_9 R_wl
Cwl_32_9 word32_9 gnd C_wl
Rw33_9 word33_9 word32_9 R_wl
Cwl_33_9 word33_9 gnd C_wl
Rw34_9 word34_9 word33_9 R_wl
Cwl_34_9 word34_9 gnd C_wl
Rw35_9 word35_9 word34_9 R_wl
Cwl_35_9 word35_9 gnd C_wl
Rw36_9 word36_9 word35_9 R_wl
Cwl_36_9 word36_9 gnd C_wl
Rw37_9 word37_9 word36_9 R_wl
Cwl_37_9 word37_9 gnd C_wl
Rw38_9 word38_9 word37_9 R_wl
Cwl_38_9 word38_9 gnd C_wl
Rw39_9 word39_9 word38_9 R_wl
Cwl_39_9 word39_9 gnd C_wl
Rw40_9 word40_9 word39_9 R_wl
Cwl_40_9 word40_9 gnd C_wl
Rw41_9 word41_9 word40_9 R_wl
Cwl_41_9 word41_9 gnd C_wl
Rw42_9 word42_9 word41_9 R_wl
Cwl_42_9 word42_9 gnd C_wl
Rw43_9 word43_9 word42_9 R_wl
Cwl_43_9 word43_9 gnd C_wl
Rw44_9 word44_9 word43_9 R_wl
Cwl_44_9 word44_9 gnd C_wl
Rw45_9 word45_9 word44_9 R_wl
Cwl_45_9 word45_9 gnd C_wl
Rw46_9 word46_9 word45_9 R_wl
Cwl_46_9 word46_9 gnd C_wl
Rw47_9 word47_9 word46_9 R_wl
Cwl_47_9 word47_9 gnd C_wl
Rw48_9 word48_9 word47_9 R_wl
Cwl_48_9 word48_9 gnd C_wl
Rw49_9 word49_9 word48_9 R_wl
Cwl_49_9 word49_9 gnd C_wl
Rw50_9 word50_9 word49_9 R_wl
Cwl_50_9 word50_9 gnd C_wl
Rw51_9 word51_9 word50_9 R_wl
Cwl_51_9 word51_9 gnd C_wl
Rw52_9 word52_9 word51_9 R_wl
Cwl_52_9 word52_9 gnd C_wl
Rw53_9 word53_9 word52_9 R_wl
Cwl_53_9 word53_9 gnd C_wl
Rw54_9 word54_9 word53_9 R_wl
Cwl_54_9 word54_9 gnd C_wl
Rw55_9 word55_9 word54_9 R_wl
Cwl_55_9 word55_9 gnd C_wl
Rw56_9 word56_9 word55_9 R_wl
Cwl_56_9 word56_9 gnd C_wl
Rw57_9 word57_9 word56_9 R_wl
Cwl_57_9 word57_9 gnd C_wl
Rw58_9 word58_9 word57_9 R_wl
Cwl_58_9 word58_9 gnd C_wl
Rw59_9 word59_9 word58_9 R_wl
Cwl_59_9 word59_9 gnd C_wl
Rw60_9 word60_9 word59_9 R_wl
Cwl_60_9 word60_9 gnd C_wl
Rw61_9 word61_9 word60_9 R_wl
Cwl_61_9 word61_9 gnd C_wl
Rw62_9 word62_9 word61_9 R_wl
Cwl_62_9 word62_9 gnd C_wl
Rw63_9 word63_9 word62_9 R_wl
Cwl_63_9 word63_9 gnd C_wl
Rw64_9 word64_9 word63_9 R_wl
Cwl_64_9 word64_9 gnd C_wl
Rw65_9 word65_9 word64_9 R_wl
Cwl_65_9 word65_9 gnd C_wl
Rw66_9 word66_9 word65_9 R_wl
Cwl_66_9 word66_9 gnd C_wl
Rw67_9 word67_9 word66_9 R_wl
Cwl_67_9 word67_9 gnd C_wl
Rw68_9 word68_9 word67_9 R_wl
Cwl_68_9 word68_9 gnd C_wl
Rw69_9 word69_9 word68_9 R_wl
Cwl_69_9 word69_9 gnd C_wl
Rw70_9 word70_9 word69_9 R_wl
Cwl_70_9 word70_9 gnd C_wl
Rw71_9 word71_9 word70_9 R_wl
Cwl_71_9 word71_9 gnd C_wl
Rw72_9 word72_9 word71_9 R_wl
Cwl_72_9 word72_9 gnd C_wl
Rw73_9 word73_9 word72_9 R_wl
Cwl_73_9 word73_9 gnd C_wl
Rw74_9 word74_9 word73_9 R_wl
Cwl_74_9 word74_9 gnd C_wl
Rw75_9 word75_9 word74_9 R_wl
Cwl_75_9 word75_9 gnd C_wl
Rw76_9 word76_9 word75_9 R_wl
Cwl_76_9 word76_9 gnd C_wl
Rw77_9 word77_9 word76_9 R_wl
Cwl_77_9 word77_9 gnd C_wl
Rw78_9 word78_9 word77_9 R_wl
Cwl_78_9 word78_9 gnd C_wl
Rw79_9 word79_9 word78_9 R_wl
Cwl_79_9 word79_9 gnd C_wl
Rw80_9 word80_9 word79_9 R_wl
Cwl_80_9 word80_9 gnd C_wl
Rw81_9 word81_9 word80_9 R_wl
Cwl_81_9 word81_9 gnd C_wl
Rw82_9 word82_9 word81_9 R_wl
Cwl_82_9 word82_9 gnd C_wl
Rw83_9 word83_9 word82_9 R_wl
Cwl_83_9 word83_9 gnd C_wl
Rw84_9 word84_9 word83_9 R_wl
Cwl_84_9 word84_9 gnd C_wl
Rw85_9 word85_9 word84_9 R_wl
Cwl_85_9 word85_9 gnd C_wl
Rw86_9 word86_9 word85_9 R_wl
Cwl_86_9 word86_9 gnd C_wl
Rw87_9 word87_9 word86_9 R_wl
Cwl_87_9 word87_9 gnd C_wl
Rw88_9 word88_9 word87_9 R_wl
Cwl_88_9 word88_9 gnd C_wl
Rw89_9 word89_9 word88_9 R_wl
Cwl_89_9 word89_9 gnd C_wl
Rw90_9 word90_9 word89_9 R_wl
Cwl_90_9 word90_9 gnd C_wl
Rw91_9 word91_9 word90_9 R_wl
Cwl_91_9 word91_9 gnd C_wl
Rw92_9 word92_9 word91_9 R_wl
Cwl_92_9 word92_9 gnd C_wl
Rw93_9 word93_9 word92_9 R_wl
Cwl_93_9 word93_9 gnd C_wl
Rw94_9 word94_9 word93_9 R_wl
Cwl_94_9 word94_9 gnd C_wl
Rw95_9 word95_9 word94_9 R_wl
Cwl_95_9 word95_9 gnd C_wl
Rw96_9 word96_9 word95_9 R_wl
Cwl_96_9 word96_9 gnd C_wl
Rw97_9 word97_9 word96_9 R_wl
Cwl_97_9 word97_9 gnd C_wl
Rw98_9 word98_9 word97_9 R_wl
Cwl_98_9 word98_9 gnd C_wl
Rw99_9 word99_9 word98_9 R_wl
Cwl_99_9 word99_9 gnd C_wl
Vwl_10 word_10 0 0
Rw0_10 word_10 word0_10 R_wl
Cwl_0_10 word0_10 gnd C_wl
Rw1_10 word1_10 word0_10 R_wl
Cwl_1_10 word1_10 gnd C_wl
Rw2_10 word2_10 word1_10 R_wl
Cwl_2_10 word2_10 gnd C_wl
Rw3_10 word3_10 word2_10 R_wl
Cwl_3_10 word3_10 gnd C_wl
Rw4_10 word4_10 word3_10 R_wl
Cwl_4_10 word4_10 gnd C_wl
Rw5_10 word5_10 word4_10 R_wl
Cwl_5_10 word5_10 gnd C_wl
Rw6_10 word6_10 word5_10 R_wl
Cwl_6_10 word6_10 gnd C_wl
Rw7_10 word7_10 word6_10 R_wl
Cwl_7_10 word7_10 gnd C_wl
Rw8_10 word8_10 word7_10 R_wl
Cwl_8_10 word8_10 gnd C_wl
Rw9_10 word9_10 word8_10 R_wl
Cwl_9_10 word9_10 gnd C_wl
Rw10_10 word10_10 word9_10 R_wl
Cwl_10_10 word10_10 gnd C_wl
Rw11_10 word11_10 word10_10 R_wl
Cwl_11_10 word11_10 gnd C_wl
Rw12_10 word12_10 word11_10 R_wl
Cwl_12_10 word12_10 gnd C_wl
Rw13_10 word13_10 word12_10 R_wl
Cwl_13_10 word13_10 gnd C_wl
Rw14_10 word14_10 word13_10 R_wl
Cwl_14_10 word14_10 gnd C_wl
Rw15_10 word15_10 word14_10 R_wl
Cwl_15_10 word15_10 gnd C_wl
Rw16_10 word16_10 word15_10 R_wl
Cwl_16_10 word16_10 gnd C_wl
Rw17_10 word17_10 word16_10 R_wl
Cwl_17_10 word17_10 gnd C_wl
Rw18_10 word18_10 word17_10 R_wl
Cwl_18_10 word18_10 gnd C_wl
Rw19_10 word19_10 word18_10 R_wl
Cwl_19_10 word19_10 gnd C_wl
Rw20_10 word20_10 word19_10 R_wl
Cwl_20_10 word20_10 gnd C_wl
Rw21_10 word21_10 word20_10 R_wl
Cwl_21_10 word21_10 gnd C_wl
Rw22_10 word22_10 word21_10 R_wl
Cwl_22_10 word22_10 gnd C_wl
Rw23_10 word23_10 word22_10 R_wl
Cwl_23_10 word23_10 gnd C_wl
Rw24_10 word24_10 word23_10 R_wl
Cwl_24_10 word24_10 gnd C_wl
Rw25_10 word25_10 word24_10 R_wl
Cwl_25_10 word25_10 gnd C_wl
Rw26_10 word26_10 word25_10 R_wl
Cwl_26_10 word26_10 gnd C_wl
Rw27_10 word27_10 word26_10 R_wl
Cwl_27_10 word27_10 gnd C_wl
Rw28_10 word28_10 word27_10 R_wl
Cwl_28_10 word28_10 gnd C_wl
Rw29_10 word29_10 word28_10 R_wl
Cwl_29_10 word29_10 gnd C_wl
Rw30_10 word30_10 word29_10 R_wl
Cwl_30_10 word30_10 gnd C_wl
Rw31_10 word31_10 word30_10 R_wl
Cwl_31_10 word31_10 gnd C_wl
Rw32_10 word32_10 word31_10 R_wl
Cwl_32_10 word32_10 gnd C_wl
Rw33_10 word33_10 word32_10 R_wl
Cwl_33_10 word33_10 gnd C_wl
Rw34_10 word34_10 word33_10 R_wl
Cwl_34_10 word34_10 gnd C_wl
Rw35_10 word35_10 word34_10 R_wl
Cwl_35_10 word35_10 gnd C_wl
Rw36_10 word36_10 word35_10 R_wl
Cwl_36_10 word36_10 gnd C_wl
Rw37_10 word37_10 word36_10 R_wl
Cwl_37_10 word37_10 gnd C_wl
Rw38_10 word38_10 word37_10 R_wl
Cwl_38_10 word38_10 gnd C_wl
Rw39_10 word39_10 word38_10 R_wl
Cwl_39_10 word39_10 gnd C_wl
Rw40_10 word40_10 word39_10 R_wl
Cwl_40_10 word40_10 gnd C_wl
Rw41_10 word41_10 word40_10 R_wl
Cwl_41_10 word41_10 gnd C_wl
Rw42_10 word42_10 word41_10 R_wl
Cwl_42_10 word42_10 gnd C_wl
Rw43_10 word43_10 word42_10 R_wl
Cwl_43_10 word43_10 gnd C_wl
Rw44_10 word44_10 word43_10 R_wl
Cwl_44_10 word44_10 gnd C_wl
Rw45_10 word45_10 word44_10 R_wl
Cwl_45_10 word45_10 gnd C_wl
Rw46_10 word46_10 word45_10 R_wl
Cwl_46_10 word46_10 gnd C_wl
Rw47_10 word47_10 word46_10 R_wl
Cwl_47_10 word47_10 gnd C_wl
Rw48_10 word48_10 word47_10 R_wl
Cwl_48_10 word48_10 gnd C_wl
Rw49_10 word49_10 word48_10 R_wl
Cwl_49_10 word49_10 gnd C_wl
Rw50_10 word50_10 word49_10 R_wl
Cwl_50_10 word50_10 gnd C_wl
Rw51_10 word51_10 word50_10 R_wl
Cwl_51_10 word51_10 gnd C_wl
Rw52_10 word52_10 word51_10 R_wl
Cwl_52_10 word52_10 gnd C_wl
Rw53_10 word53_10 word52_10 R_wl
Cwl_53_10 word53_10 gnd C_wl
Rw54_10 word54_10 word53_10 R_wl
Cwl_54_10 word54_10 gnd C_wl
Rw55_10 word55_10 word54_10 R_wl
Cwl_55_10 word55_10 gnd C_wl
Rw56_10 word56_10 word55_10 R_wl
Cwl_56_10 word56_10 gnd C_wl
Rw57_10 word57_10 word56_10 R_wl
Cwl_57_10 word57_10 gnd C_wl
Rw58_10 word58_10 word57_10 R_wl
Cwl_58_10 word58_10 gnd C_wl
Rw59_10 word59_10 word58_10 R_wl
Cwl_59_10 word59_10 gnd C_wl
Rw60_10 word60_10 word59_10 R_wl
Cwl_60_10 word60_10 gnd C_wl
Rw61_10 word61_10 word60_10 R_wl
Cwl_61_10 word61_10 gnd C_wl
Rw62_10 word62_10 word61_10 R_wl
Cwl_62_10 word62_10 gnd C_wl
Rw63_10 word63_10 word62_10 R_wl
Cwl_63_10 word63_10 gnd C_wl
Rw64_10 word64_10 word63_10 R_wl
Cwl_64_10 word64_10 gnd C_wl
Rw65_10 word65_10 word64_10 R_wl
Cwl_65_10 word65_10 gnd C_wl
Rw66_10 word66_10 word65_10 R_wl
Cwl_66_10 word66_10 gnd C_wl
Rw67_10 word67_10 word66_10 R_wl
Cwl_67_10 word67_10 gnd C_wl
Rw68_10 word68_10 word67_10 R_wl
Cwl_68_10 word68_10 gnd C_wl
Rw69_10 word69_10 word68_10 R_wl
Cwl_69_10 word69_10 gnd C_wl
Rw70_10 word70_10 word69_10 R_wl
Cwl_70_10 word70_10 gnd C_wl
Rw71_10 word71_10 word70_10 R_wl
Cwl_71_10 word71_10 gnd C_wl
Rw72_10 word72_10 word71_10 R_wl
Cwl_72_10 word72_10 gnd C_wl
Rw73_10 word73_10 word72_10 R_wl
Cwl_73_10 word73_10 gnd C_wl
Rw74_10 word74_10 word73_10 R_wl
Cwl_74_10 word74_10 gnd C_wl
Rw75_10 word75_10 word74_10 R_wl
Cwl_75_10 word75_10 gnd C_wl
Rw76_10 word76_10 word75_10 R_wl
Cwl_76_10 word76_10 gnd C_wl
Rw77_10 word77_10 word76_10 R_wl
Cwl_77_10 word77_10 gnd C_wl
Rw78_10 word78_10 word77_10 R_wl
Cwl_78_10 word78_10 gnd C_wl
Rw79_10 word79_10 word78_10 R_wl
Cwl_79_10 word79_10 gnd C_wl
Rw80_10 word80_10 word79_10 R_wl
Cwl_80_10 word80_10 gnd C_wl
Rw81_10 word81_10 word80_10 R_wl
Cwl_81_10 word81_10 gnd C_wl
Rw82_10 word82_10 word81_10 R_wl
Cwl_82_10 word82_10 gnd C_wl
Rw83_10 word83_10 word82_10 R_wl
Cwl_83_10 word83_10 gnd C_wl
Rw84_10 word84_10 word83_10 R_wl
Cwl_84_10 word84_10 gnd C_wl
Rw85_10 word85_10 word84_10 R_wl
Cwl_85_10 word85_10 gnd C_wl
Rw86_10 word86_10 word85_10 R_wl
Cwl_86_10 word86_10 gnd C_wl
Rw87_10 word87_10 word86_10 R_wl
Cwl_87_10 word87_10 gnd C_wl
Rw88_10 word88_10 word87_10 R_wl
Cwl_88_10 word88_10 gnd C_wl
Rw89_10 word89_10 word88_10 R_wl
Cwl_89_10 word89_10 gnd C_wl
Rw90_10 word90_10 word89_10 R_wl
Cwl_90_10 word90_10 gnd C_wl
Rw91_10 word91_10 word90_10 R_wl
Cwl_91_10 word91_10 gnd C_wl
Rw92_10 word92_10 word91_10 R_wl
Cwl_92_10 word92_10 gnd C_wl
Rw93_10 word93_10 word92_10 R_wl
Cwl_93_10 word93_10 gnd C_wl
Rw94_10 word94_10 word93_10 R_wl
Cwl_94_10 word94_10 gnd C_wl
Rw95_10 word95_10 word94_10 R_wl
Cwl_95_10 word95_10 gnd C_wl
Rw96_10 word96_10 word95_10 R_wl
Cwl_96_10 word96_10 gnd C_wl
Rw97_10 word97_10 word96_10 R_wl
Cwl_97_10 word97_10 gnd C_wl
Rw98_10 word98_10 word97_10 R_wl
Cwl_98_10 word98_10 gnd C_wl
Rw99_10 word99_10 word98_10 R_wl
Cwl_99_10 word99_10 gnd C_wl
Vwl_11 word_11 0 0
Rw0_11 word_11 word0_11 R_wl
Cwl_0_11 word0_11 gnd C_wl
Rw1_11 word1_11 word0_11 R_wl
Cwl_1_11 word1_11 gnd C_wl
Rw2_11 word2_11 word1_11 R_wl
Cwl_2_11 word2_11 gnd C_wl
Rw3_11 word3_11 word2_11 R_wl
Cwl_3_11 word3_11 gnd C_wl
Rw4_11 word4_11 word3_11 R_wl
Cwl_4_11 word4_11 gnd C_wl
Rw5_11 word5_11 word4_11 R_wl
Cwl_5_11 word5_11 gnd C_wl
Rw6_11 word6_11 word5_11 R_wl
Cwl_6_11 word6_11 gnd C_wl
Rw7_11 word7_11 word6_11 R_wl
Cwl_7_11 word7_11 gnd C_wl
Rw8_11 word8_11 word7_11 R_wl
Cwl_8_11 word8_11 gnd C_wl
Rw9_11 word9_11 word8_11 R_wl
Cwl_9_11 word9_11 gnd C_wl
Rw10_11 word10_11 word9_11 R_wl
Cwl_10_11 word10_11 gnd C_wl
Rw11_11 word11_11 word10_11 R_wl
Cwl_11_11 word11_11 gnd C_wl
Rw12_11 word12_11 word11_11 R_wl
Cwl_12_11 word12_11 gnd C_wl
Rw13_11 word13_11 word12_11 R_wl
Cwl_13_11 word13_11 gnd C_wl
Rw14_11 word14_11 word13_11 R_wl
Cwl_14_11 word14_11 gnd C_wl
Rw15_11 word15_11 word14_11 R_wl
Cwl_15_11 word15_11 gnd C_wl
Rw16_11 word16_11 word15_11 R_wl
Cwl_16_11 word16_11 gnd C_wl
Rw17_11 word17_11 word16_11 R_wl
Cwl_17_11 word17_11 gnd C_wl
Rw18_11 word18_11 word17_11 R_wl
Cwl_18_11 word18_11 gnd C_wl
Rw19_11 word19_11 word18_11 R_wl
Cwl_19_11 word19_11 gnd C_wl
Rw20_11 word20_11 word19_11 R_wl
Cwl_20_11 word20_11 gnd C_wl
Rw21_11 word21_11 word20_11 R_wl
Cwl_21_11 word21_11 gnd C_wl
Rw22_11 word22_11 word21_11 R_wl
Cwl_22_11 word22_11 gnd C_wl
Rw23_11 word23_11 word22_11 R_wl
Cwl_23_11 word23_11 gnd C_wl
Rw24_11 word24_11 word23_11 R_wl
Cwl_24_11 word24_11 gnd C_wl
Rw25_11 word25_11 word24_11 R_wl
Cwl_25_11 word25_11 gnd C_wl
Rw26_11 word26_11 word25_11 R_wl
Cwl_26_11 word26_11 gnd C_wl
Rw27_11 word27_11 word26_11 R_wl
Cwl_27_11 word27_11 gnd C_wl
Rw28_11 word28_11 word27_11 R_wl
Cwl_28_11 word28_11 gnd C_wl
Rw29_11 word29_11 word28_11 R_wl
Cwl_29_11 word29_11 gnd C_wl
Rw30_11 word30_11 word29_11 R_wl
Cwl_30_11 word30_11 gnd C_wl
Rw31_11 word31_11 word30_11 R_wl
Cwl_31_11 word31_11 gnd C_wl
Rw32_11 word32_11 word31_11 R_wl
Cwl_32_11 word32_11 gnd C_wl
Rw33_11 word33_11 word32_11 R_wl
Cwl_33_11 word33_11 gnd C_wl
Rw34_11 word34_11 word33_11 R_wl
Cwl_34_11 word34_11 gnd C_wl
Rw35_11 word35_11 word34_11 R_wl
Cwl_35_11 word35_11 gnd C_wl
Rw36_11 word36_11 word35_11 R_wl
Cwl_36_11 word36_11 gnd C_wl
Rw37_11 word37_11 word36_11 R_wl
Cwl_37_11 word37_11 gnd C_wl
Rw38_11 word38_11 word37_11 R_wl
Cwl_38_11 word38_11 gnd C_wl
Rw39_11 word39_11 word38_11 R_wl
Cwl_39_11 word39_11 gnd C_wl
Rw40_11 word40_11 word39_11 R_wl
Cwl_40_11 word40_11 gnd C_wl
Rw41_11 word41_11 word40_11 R_wl
Cwl_41_11 word41_11 gnd C_wl
Rw42_11 word42_11 word41_11 R_wl
Cwl_42_11 word42_11 gnd C_wl
Rw43_11 word43_11 word42_11 R_wl
Cwl_43_11 word43_11 gnd C_wl
Rw44_11 word44_11 word43_11 R_wl
Cwl_44_11 word44_11 gnd C_wl
Rw45_11 word45_11 word44_11 R_wl
Cwl_45_11 word45_11 gnd C_wl
Rw46_11 word46_11 word45_11 R_wl
Cwl_46_11 word46_11 gnd C_wl
Rw47_11 word47_11 word46_11 R_wl
Cwl_47_11 word47_11 gnd C_wl
Rw48_11 word48_11 word47_11 R_wl
Cwl_48_11 word48_11 gnd C_wl
Rw49_11 word49_11 word48_11 R_wl
Cwl_49_11 word49_11 gnd C_wl
Rw50_11 word50_11 word49_11 R_wl
Cwl_50_11 word50_11 gnd C_wl
Rw51_11 word51_11 word50_11 R_wl
Cwl_51_11 word51_11 gnd C_wl
Rw52_11 word52_11 word51_11 R_wl
Cwl_52_11 word52_11 gnd C_wl
Rw53_11 word53_11 word52_11 R_wl
Cwl_53_11 word53_11 gnd C_wl
Rw54_11 word54_11 word53_11 R_wl
Cwl_54_11 word54_11 gnd C_wl
Rw55_11 word55_11 word54_11 R_wl
Cwl_55_11 word55_11 gnd C_wl
Rw56_11 word56_11 word55_11 R_wl
Cwl_56_11 word56_11 gnd C_wl
Rw57_11 word57_11 word56_11 R_wl
Cwl_57_11 word57_11 gnd C_wl
Rw58_11 word58_11 word57_11 R_wl
Cwl_58_11 word58_11 gnd C_wl
Rw59_11 word59_11 word58_11 R_wl
Cwl_59_11 word59_11 gnd C_wl
Rw60_11 word60_11 word59_11 R_wl
Cwl_60_11 word60_11 gnd C_wl
Rw61_11 word61_11 word60_11 R_wl
Cwl_61_11 word61_11 gnd C_wl
Rw62_11 word62_11 word61_11 R_wl
Cwl_62_11 word62_11 gnd C_wl
Rw63_11 word63_11 word62_11 R_wl
Cwl_63_11 word63_11 gnd C_wl
Rw64_11 word64_11 word63_11 R_wl
Cwl_64_11 word64_11 gnd C_wl
Rw65_11 word65_11 word64_11 R_wl
Cwl_65_11 word65_11 gnd C_wl
Rw66_11 word66_11 word65_11 R_wl
Cwl_66_11 word66_11 gnd C_wl
Rw67_11 word67_11 word66_11 R_wl
Cwl_67_11 word67_11 gnd C_wl
Rw68_11 word68_11 word67_11 R_wl
Cwl_68_11 word68_11 gnd C_wl
Rw69_11 word69_11 word68_11 R_wl
Cwl_69_11 word69_11 gnd C_wl
Rw70_11 word70_11 word69_11 R_wl
Cwl_70_11 word70_11 gnd C_wl
Rw71_11 word71_11 word70_11 R_wl
Cwl_71_11 word71_11 gnd C_wl
Rw72_11 word72_11 word71_11 R_wl
Cwl_72_11 word72_11 gnd C_wl
Rw73_11 word73_11 word72_11 R_wl
Cwl_73_11 word73_11 gnd C_wl
Rw74_11 word74_11 word73_11 R_wl
Cwl_74_11 word74_11 gnd C_wl
Rw75_11 word75_11 word74_11 R_wl
Cwl_75_11 word75_11 gnd C_wl
Rw76_11 word76_11 word75_11 R_wl
Cwl_76_11 word76_11 gnd C_wl
Rw77_11 word77_11 word76_11 R_wl
Cwl_77_11 word77_11 gnd C_wl
Rw78_11 word78_11 word77_11 R_wl
Cwl_78_11 word78_11 gnd C_wl
Rw79_11 word79_11 word78_11 R_wl
Cwl_79_11 word79_11 gnd C_wl
Rw80_11 word80_11 word79_11 R_wl
Cwl_80_11 word80_11 gnd C_wl
Rw81_11 word81_11 word80_11 R_wl
Cwl_81_11 word81_11 gnd C_wl
Rw82_11 word82_11 word81_11 R_wl
Cwl_82_11 word82_11 gnd C_wl
Rw83_11 word83_11 word82_11 R_wl
Cwl_83_11 word83_11 gnd C_wl
Rw84_11 word84_11 word83_11 R_wl
Cwl_84_11 word84_11 gnd C_wl
Rw85_11 word85_11 word84_11 R_wl
Cwl_85_11 word85_11 gnd C_wl
Rw86_11 word86_11 word85_11 R_wl
Cwl_86_11 word86_11 gnd C_wl
Rw87_11 word87_11 word86_11 R_wl
Cwl_87_11 word87_11 gnd C_wl
Rw88_11 word88_11 word87_11 R_wl
Cwl_88_11 word88_11 gnd C_wl
Rw89_11 word89_11 word88_11 R_wl
Cwl_89_11 word89_11 gnd C_wl
Rw90_11 word90_11 word89_11 R_wl
Cwl_90_11 word90_11 gnd C_wl
Rw91_11 word91_11 word90_11 R_wl
Cwl_91_11 word91_11 gnd C_wl
Rw92_11 word92_11 word91_11 R_wl
Cwl_92_11 word92_11 gnd C_wl
Rw93_11 word93_11 word92_11 R_wl
Cwl_93_11 word93_11 gnd C_wl
Rw94_11 word94_11 word93_11 R_wl
Cwl_94_11 word94_11 gnd C_wl
Rw95_11 word95_11 word94_11 R_wl
Cwl_95_11 word95_11 gnd C_wl
Rw96_11 word96_11 word95_11 R_wl
Cwl_96_11 word96_11 gnd C_wl
Rw97_11 word97_11 word96_11 R_wl
Cwl_97_11 word97_11 gnd C_wl
Rw98_11 word98_11 word97_11 R_wl
Cwl_98_11 word98_11 gnd C_wl
Rw99_11 word99_11 word98_11 R_wl
Cwl_99_11 word99_11 gnd C_wl
Vwl_12 word_12 0 0
Rw0_12 word_12 word0_12 R_wl
Cwl_0_12 word0_12 gnd C_wl
Rw1_12 word1_12 word0_12 R_wl
Cwl_1_12 word1_12 gnd C_wl
Rw2_12 word2_12 word1_12 R_wl
Cwl_2_12 word2_12 gnd C_wl
Rw3_12 word3_12 word2_12 R_wl
Cwl_3_12 word3_12 gnd C_wl
Rw4_12 word4_12 word3_12 R_wl
Cwl_4_12 word4_12 gnd C_wl
Rw5_12 word5_12 word4_12 R_wl
Cwl_5_12 word5_12 gnd C_wl
Rw6_12 word6_12 word5_12 R_wl
Cwl_6_12 word6_12 gnd C_wl
Rw7_12 word7_12 word6_12 R_wl
Cwl_7_12 word7_12 gnd C_wl
Rw8_12 word8_12 word7_12 R_wl
Cwl_8_12 word8_12 gnd C_wl
Rw9_12 word9_12 word8_12 R_wl
Cwl_9_12 word9_12 gnd C_wl
Rw10_12 word10_12 word9_12 R_wl
Cwl_10_12 word10_12 gnd C_wl
Rw11_12 word11_12 word10_12 R_wl
Cwl_11_12 word11_12 gnd C_wl
Rw12_12 word12_12 word11_12 R_wl
Cwl_12_12 word12_12 gnd C_wl
Rw13_12 word13_12 word12_12 R_wl
Cwl_13_12 word13_12 gnd C_wl
Rw14_12 word14_12 word13_12 R_wl
Cwl_14_12 word14_12 gnd C_wl
Rw15_12 word15_12 word14_12 R_wl
Cwl_15_12 word15_12 gnd C_wl
Rw16_12 word16_12 word15_12 R_wl
Cwl_16_12 word16_12 gnd C_wl
Rw17_12 word17_12 word16_12 R_wl
Cwl_17_12 word17_12 gnd C_wl
Rw18_12 word18_12 word17_12 R_wl
Cwl_18_12 word18_12 gnd C_wl
Rw19_12 word19_12 word18_12 R_wl
Cwl_19_12 word19_12 gnd C_wl
Rw20_12 word20_12 word19_12 R_wl
Cwl_20_12 word20_12 gnd C_wl
Rw21_12 word21_12 word20_12 R_wl
Cwl_21_12 word21_12 gnd C_wl
Rw22_12 word22_12 word21_12 R_wl
Cwl_22_12 word22_12 gnd C_wl
Rw23_12 word23_12 word22_12 R_wl
Cwl_23_12 word23_12 gnd C_wl
Rw24_12 word24_12 word23_12 R_wl
Cwl_24_12 word24_12 gnd C_wl
Rw25_12 word25_12 word24_12 R_wl
Cwl_25_12 word25_12 gnd C_wl
Rw26_12 word26_12 word25_12 R_wl
Cwl_26_12 word26_12 gnd C_wl
Rw27_12 word27_12 word26_12 R_wl
Cwl_27_12 word27_12 gnd C_wl
Rw28_12 word28_12 word27_12 R_wl
Cwl_28_12 word28_12 gnd C_wl
Rw29_12 word29_12 word28_12 R_wl
Cwl_29_12 word29_12 gnd C_wl
Rw30_12 word30_12 word29_12 R_wl
Cwl_30_12 word30_12 gnd C_wl
Rw31_12 word31_12 word30_12 R_wl
Cwl_31_12 word31_12 gnd C_wl
Rw32_12 word32_12 word31_12 R_wl
Cwl_32_12 word32_12 gnd C_wl
Rw33_12 word33_12 word32_12 R_wl
Cwl_33_12 word33_12 gnd C_wl
Rw34_12 word34_12 word33_12 R_wl
Cwl_34_12 word34_12 gnd C_wl
Rw35_12 word35_12 word34_12 R_wl
Cwl_35_12 word35_12 gnd C_wl
Rw36_12 word36_12 word35_12 R_wl
Cwl_36_12 word36_12 gnd C_wl
Rw37_12 word37_12 word36_12 R_wl
Cwl_37_12 word37_12 gnd C_wl
Rw38_12 word38_12 word37_12 R_wl
Cwl_38_12 word38_12 gnd C_wl
Rw39_12 word39_12 word38_12 R_wl
Cwl_39_12 word39_12 gnd C_wl
Rw40_12 word40_12 word39_12 R_wl
Cwl_40_12 word40_12 gnd C_wl
Rw41_12 word41_12 word40_12 R_wl
Cwl_41_12 word41_12 gnd C_wl
Rw42_12 word42_12 word41_12 R_wl
Cwl_42_12 word42_12 gnd C_wl
Rw43_12 word43_12 word42_12 R_wl
Cwl_43_12 word43_12 gnd C_wl
Rw44_12 word44_12 word43_12 R_wl
Cwl_44_12 word44_12 gnd C_wl
Rw45_12 word45_12 word44_12 R_wl
Cwl_45_12 word45_12 gnd C_wl
Rw46_12 word46_12 word45_12 R_wl
Cwl_46_12 word46_12 gnd C_wl
Rw47_12 word47_12 word46_12 R_wl
Cwl_47_12 word47_12 gnd C_wl
Rw48_12 word48_12 word47_12 R_wl
Cwl_48_12 word48_12 gnd C_wl
Rw49_12 word49_12 word48_12 R_wl
Cwl_49_12 word49_12 gnd C_wl
Rw50_12 word50_12 word49_12 R_wl
Cwl_50_12 word50_12 gnd C_wl
Rw51_12 word51_12 word50_12 R_wl
Cwl_51_12 word51_12 gnd C_wl
Rw52_12 word52_12 word51_12 R_wl
Cwl_52_12 word52_12 gnd C_wl
Rw53_12 word53_12 word52_12 R_wl
Cwl_53_12 word53_12 gnd C_wl
Rw54_12 word54_12 word53_12 R_wl
Cwl_54_12 word54_12 gnd C_wl
Rw55_12 word55_12 word54_12 R_wl
Cwl_55_12 word55_12 gnd C_wl
Rw56_12 word56_12 word55_12 R_wl
Cwl_56_12 word56_12 gnd C_wl
Rw57_12 word57_12 word56_12 R_wl
Cwl_57_12 word57_12 gnd C_wl
Rw58_12 word58_12 word57_12 R_wl
Cwl_58_12 word58_12 gnd C_wl
Rw59_12 word59_12 word58_12 R_wl
Cwl_59_12 word59_12 gnd C_wl
Rw60_12 word60_12 word59_12 R_wl
Cwl_60_12 word60_12 gnd C_wl
Rw61_12 word61_12 word60_12 R_wl
Cwl_61_12 word61_12 gnd C_wl
Rw62_12 word62_12 word61_12 R_wl
Cwl_62_12 word62_12 gnd C_wl
Rw63_12 word63_12 word62_12 R_wl
Cwl_63_12 word63_12 gnd C_wl
Rw64_12 word64_12 word63_12 R_wl
Cwl_64_12 word64_12 gnd C_wl
Rw65_12 word65_12 word64_12 R_wl
Cwl_65_12 word65_12 gnd C_wl
Rw66_12 word66_12 word65_12 R_wl
Cwl_66_12 word66_12 gnd C_wl
Rw67_12 word67_12 word66_12 R_wl
Cwl_67_12 word67_12 gnd C_wl
Rw68_12 word68_12 word67_12 R_wl
Cwl_68_12 word68_12 gnd C_wl
Rw69_12 word69_12 word68_12 R_wl
Cwl_69_12 word69_12 gnd C_wl
Rw70_12 word70_12 word69_12 R_wl
Cwl_70_12 word70_12 gnd C_wl
Rw71_12 word71_12 word70_12 R_wl
Cwl_71_12 word71_12 gnd C_wl
Rw72_12 word72_12 word71_12 R_wl
Cwl_72_12 word72_12 gnd C_wl
Rw73_12 word73_12 word72_12 R_wl
Cwl_73_12 word73_12 gnd C_wl
Rw74_12 word74_12 word73_12 R_wl
Cwl_74_12 word74_12 gnd C_wl
Rw75_12 word75_12 word74_12 R_wl
Cwl_75_12 word75_12 gnd C_wl
Rw76_12 word76_12 word75_12 R_wl
Cwl_76_12 word76_12 gnd C_wl
Rw77_12 word77_12 word76_12 R_wl
Cwl_77_12 word77_12 gnd C_wl
Rw78_12 word78_12 word77_12 R_wl
Cwl_78_12 word78_12 gnd C_wl
Rw79_12 word79_12 word78_12 R_wl
Cwl_79_12 word79_12 gnd C_wl
Rw80_12 word80_12 word79_12 R_wl
Cwl_80_12 word80_12 gnd C_wl
Rw81_12 word81_12 word80_12 R_wl
Cwl_81_12 word81_12 gnd C_wl
Rw82_12 word82_12 word81_12 R_wl
Cwl_82_12 word82_12 gnd C_wl
Rw83_12 word83_12 word82_12 R_wl
Cwl_83_12 word83_12 gnd C_wl
Rw84_12 word84_12 word83_12 R_wl
Cwl_84_12 word84_12 gnd C_wl
Rw85_12 word85_12 word84_12 R_wl
Cwl_85_12 word85_12 gnd C_wl
Rw86_12 word86_12 word85_12 R_wl
Cwl_86_12 word86_12 gnd C_wl
Rw87_12 word87_12 word86_12 R_wl
Cwl_87_12 word87_12 gnd C_wl
Rw88_12 word88_12 word87_12 R_wl
Cwl_88_12 word88_12 gnd C_wl
Rw89_12 word89_12 word88_12 R_wl
Cwl_89_12 word89_12 gnd C_wl
Rw90_12 word90_12 word89_12 R_wl
Cwl_90_12 word90_12 gnd C_wl
Rw91_12 word91_12 word90_12 R_wl
Cwl_91_12 word91_12 gnd C_wl
Rw92_12 word92_12 word91_12 R_wl
Cwl_92_12 word92_12 gnd C_wl
Rw93_12 word93_12 word92_12 R_wl
Cwl_93_12 word93_12 gnd C_wl
Rw94_12 word94_12 word93_12 R_wl
Cwl_94_12 word94_12 gnd C_wl
Rw95_12 word95_12 word94_12 R_wl
Cwl_95_12 word95_12 gnd C_wl
Rw96_12 word96_12 word95_12 R_wl
Cwl_96_12 word96_12 gnd C_wl
Rw97_12 word97_12 word96_12 R_wl
Cwl_97_12 word97_12 gnd C_wl
Rw98_12 word98_12 word97_12 R_wl
Cwl_98_12 word98_12 gnd C_wl
Rw99_12 word99_12 word98_12 R_wl
Cwl_99_12 word99_12 gnd C_wl
Vwl_13 word_13 0 0
Rw0_13 word_13 word0_13 R_wl
Cwl_0_13 word0_13 gnd C_wl
Rw1_13 word1_13 word0_13 R_wl
Cwl_1_13 word1_13 gnd C_wl
Rw2_13 word2_13 word1_13 R_wl
Cwl_2_13 word2_13 gnd C_wl
Rw3_13 word3_13 word2_13 R_wl
Cwl_3_13 word3_13 gnd C_wl
Rw4_13 word4_13 word3_13 R_wl
Cwl_4_13 word4_13 gnd C_wl
Rw5_13 word5_13 word4_13 R_wl
Cwl_5_13 word5_13 gnd C_wl
Rw6_13 word6_13 word5_13 R_wl
Cwl_6_13 word6_13 gnd C_wl
Rw7_13 word7_13 word6_13 R_wl
Cwl_7_13 word7_13 gnd C_wl
Rw8_13 word8_13 word7_13 R_wl
Cwl_8_13 word8_13 gnd C_wl
Rw9_13 word9_13 word8_13 R_wl
Cwl_9_13 word9_13 gnd C_wl
Rw10_13 word10_13 word9_13 R_wl
Cwl_10_13 word10_13 gnd C_wl
Rw11_13 word11_13 word10_13 R_wl
Cwl_11_13 word11_13 gnd C_wl
Rw12_13 word12_13 word11_13 R_wl
Cwl_12_13 word12_13 gnd C_wl
Rw13_13 word13_13 word12_13 R_wl
Cwl_13_13 word13_13 gnd C_wl
Rw14_13 word14_13 word13_13 R_wl
Cwl_14_13 word14_13 gnd C_wl
Rw15_13 word15_13 word14_13 R_wl
Cwl_15_13 word15_13 gnd C_wl
Rw16_13 word16_13 word15_13 R_wl
Cwl_16_13 word16_13 gnd C_wl
Rw17_13 word17_13 word16_13 R_wl
Cwl_17_13 word17_13 gnd C_wl
Rw18_13 word18_13 word17_13 R_wl
Cwl_18_13 word18_13 gnd C_wl
Rw19_13 word19_13 word18_13 R_wl
Cwl_19_13 word19_13 gnd C_wl
Rw20_13 word20_13 word19_13 R_wl
Cwl_20_13 word20_13 gnd C_wl
Rw21_13 word21_13 word20_13 R_wl
Cwl_21_13 word21_13 gnd C_wl
Rw22_13 word22_13 word21_13 R_wl
Cwl_22_13 word22_13 gnd C_wl
Rw23_13 word23_13 word22_13 R_wl
Cwl_23_13 word23_13 gnd C_wl
Rw24_13 word24_13 word23_13 R_wl
Cwl_24_13 word24_13 gnd C_wl
Rw25_13 word25_13 word24_13 R_wl
Cwl_25_13 word25_13 gnd C_wl
Rw26_13 word26_13 word25_13 R_wl
Cwl_26_13 word26_13 gnd C_wl
Rw27_13 word27_13 word26_13 R_wl
Cwl_27_13 word27_13 gnd C_wl
Rw28_13 word28_13 word27_13 R_wl
Cwl_28_13 word28_13 gnd C_wl
Rw29_13 word29_13 word28_13 R_wl
Cwl_29_13 word29_13 gnd C_wl
Rw30_13 word30_13 word29_13 R_wl
Cwl_30_13 word30_13 gnd C_wl
Rw31_13 word31_13 word30_13 R_wl
Cwl_31_13 word31_13 gnd C_wl
Rw32_13 word32_13 word31_13 R_wl
Cwl_32_13 word32_13 gnd C_wl
Rw33_13 word33_13 word32_13 R_wl
Cwl_33_13 word33_13 gnd C_wl
Rw34_13 word34_13 word33_13 R_wl
Cwl_34_13 word34_13 gnd C_wl
Rw35_13 word35_13 word34_13 R_wl
Cwl_35_13 word35_13 gnd C_wl
Rw36_13 word36_13 word35_13 R_wl
Cwl_36_13 word36_13 gnd C_wl
Rw37_13 word37_13 word36_13 R_wl
Cwl_37_13 word37_13 gnd C_wl
Rw38_13 word38_13 word37_13 R_wl
Cwl_38_13 word38_13 gnd C_wl
Rw39_13 word39_13 word38_13 R_wl
Cwl_39_13 word39_13 gnd C_wl
Rw40_13 word40_13 word39_13 R_wl
Cwl_40_13 word40_13 gnd C_wl
Rw41_13 word41_13 word40_13 R_wl
Cwl_41_13 word41_13 gnd C_wl
Rw42_13 word42_13 word41_13 R_wl
Cwl_42_13 word42_13 gnd C_wl
Rw43_13 word43_13 word42_13 R_wl
Cwl_43_13 word43_13 gnd C_wl
Rw44_13 word44_13 word43_13 R_wl
Cwl_44_13 word44_13 gnd C_wl
Rw45_13 word45_13 word44_13 R_wl
Cwl_45_13 word45_13 gnd C_wl
Rw46_13 word46_13 word45_13 R_wl
Cwl_46_13 word46_13 gnd C_wl
Rw47_13 word47_13 word46_13 R_wl
Cwl_47_13 word47_13 gnd C_wl
Rw48_13 word48_13 word47_13 R_wl
Cwl_48_13 word48_13 gnd C_wl
Rw49_13 word49_13 word48_13 R_wl
Cwl_49_13 word49_13 gnd C_wl
Rw50_13 word50_13 word49_13 R_wl
Cwl_50_13 word50_13 gnd C_wl
Rw51_13 word51_13 word50_13 R_wl
Cwl_51_13 word51_13 gnd C_wl
Rw52_13 word52_13 word51_13 R_wl
Cwl_52_13 word52_13 gnd C_wl
Rw53_13 word53_13 word52_13 R_wl
Cwl_53_13 word53_13 gnd C_wl
Rw54_13 word54_13 word53_13 R_wl
Cwl_54_13 word54_13 gnd C_wl
Rw55_13 word55_13 word54_13 R_wl
Cwl_55_13 word55_13 gnd C_wl
Rw56_13 word56_13 word55_13 R_wl
Cwl_56_13 word56_13 gnd C_wl
Rw57_13 word57_13 word56_13 R_wl
Cwl_57_13 word57_13 gnd C_wl
Rw58_13 word58_13 word57_13 R_wl
Cwl_58_13 word58_13 gnd C_wl
Rw59_13 word59_13 word58_13 R_wl
Cwl_59_13 word59_13 gnd C_wl
Rw60_13 word60_13 word59_13 R_wl
Cwl_60_13 word60_13 gnd C_wl
Rw61_13 word61_13 word60_13 R_wl
Cwl_61_13 word61_13 gnd C_wl
Rw62_13 word62_13 word61_13 R_wl
Cwl_62_13 word62_13 gnd C_wl
Rw63_13 word63_13 word62_13 R_wl
Cwl_63_13 word63_13 gnd C_wl
Rw64_13 word64_13 word63_13 R_wl
Cwl_64_13 word64_13 gnd C_wl
Rw65_13 word65_13 word64_13 R_wl
Cwl_65_13 word65_13 gnd C_wl
Rw66_13 word66_13 word65_13 R_wl
Cwl_66_13 word66_13 gnd C_wl
Rw67_13 word67_13 word66_13 R_wl
Cwl_67_13 word67_13 gnd C_wl
Rw68_13 word68_13 word67_13 R_wl
Cwl_68_13 word68_13 gnd C_wl
Rw69_13 word69_13 word68_13 R_wl
Cwl_69_13 word69_13 gnd C_wl
Rw70_13 word70_13 word69_13 R_wl
Cwl_70_13 word70_13 gnd C_wl
Rw71_13 word71_13 word70_13 R_wl
Cwl_71_13 word71_13 gnd C_wl
Rw72_13 word72_13 word71_13 R_wl
Cwl_72_13 word72_13 gnd C_wl
Rw73_13 word73_13 word72_13 R_wl
Cwl_73_13 word73_13 gnd C_wl
Rw74_13 word74_13 word73_13 R_wl
Cwl_74_13 word74_13 gnd C_wl
Rw75_13 word75_13 word74_13 R_wl
Cwl_75_13 word75_13 gnd C_wl
Rw76_13 word76_13 word75_13 R_wl
Cwl_76_13 word76_13 gnd C_wl
Rw77_13 word77_13 word76_13 R_wl
Cwl_77_13 word77_13 gnd C_wl
Rw78_13 word78_13 word77_13 R_wl
Cwl_78_13 word78_13 gnd C_wl
Rw79_13 word79_13 word78_13 R_wl
Cwl_79_13 word79_13 gnd C_wl
Rw80_13 word80_13 word79_13 R_wl
Cwl_80_13 word80_13 gnd C_wl
Rw81_13 word81_13 word80_13 R_wl
Cwl_81_13 word81_13 gnd C_wl
Rw82_13 word82_13 word81_13 R_wl
Cwl_82_13 word82_13 gnd C_wl
Rw83_13 word83_13 word82_13 R_wl
Cwl_83_13 word83_13 gnd C_wl
Rw84_13 word84_13 word83_13 R_wl
Cwl_84_13 word84_13 gnd C_wl
Rw85_13 word85_13 word84_13 R_wl
Cwl_85_13 word85_13 gnd C_wl
Rw86_13 word86_13 word85_13 R_wl
Cwl_86_13 word86_13 gnd C_wl
Rw87_13 word87_13 word86_13 R_wl
Cwl_87_13 word87_13 gnd C_wl
Rw88_13 word88_13 word87_13 R_wl
Cwl_88_13 word88_13 gnd C_wl
Rw89_13 word89_13 word88_13 R_wl
Cwl_89_13 word89_13 gnd C_wl
Rw90_13 word90_13 word89_13 R_wl
Cwl_90_13 word90_13 gnd C_wl
Rw91_13 word91_13 word90_13 R_wl
Cwl_91_13 word91_13 gnd C_wl
Rw92_13 word92_13 word91_13 R_wl
Cwl_92_13 word92_13 gnd C_wl
Rw93_13 word93_13 word92_13 R_wl
Cwl_93_13 word93_13 gnd C_wl
Rw94_13 word94_13 word93_13 R_wl
Cwl_94_13 word94_13 gnd C_wl
Rw95_13 word95_13 word94_13 R_wl
Cwl_95_13 word95_13 gnd C_wl
Rw96_13 word96_13 word95_13 R_wl
Cwl_96_13 word96_13 gnd C_wl
Rw97_13 word97_13 word96_13 R_wl
Cwl_97_13 word97_13 gnd C_wl
Rw98_13 word98_13 word97_13 R_wl
Cwl_98_13 word98_13 gnd C_wl
Rw99_13 word99_13 word98_13 R_wl
Cwl_99_13 word99_13 gnd C_wl
Vwl_14 word_14 0 0
Rw0_14 word_14 word0_14 R_wl
Cwl_0_14 word0_14 gnd C_wl
Rw1_14 word1_14 word0_14 R_wl
Cwl_1_14 word1_14 gnd C_wl
Rw2_14 word2_14 word1_14 R_wl
Cwl_2_14 word2_14 gnd C_wl
Rw3_14 word3_14 word2_14 R_wl
Cwl_3_14 word3_14 gnd C_wl
Rw4_14 word4_14 word3_14 R_wl
Cwl_4_14 word4_14 gnd C_wl
Rw5_14 word5_14 word4_14 R_wl
Cwl_5_14 word5_14 gnd C_wl
Rw6_14 word6_14 word5_14 R_wl
Cwl_6_14 word6_14 gnd C_wl
Rw7_14 word7_14 word6_14 R_wl
Cwl_7_14 word7_14 gnd C_wl
Rw8_14 word8_14 word7_14 R_wl
Cwl_8_14 word8_14 gnd C_wl
Rw9_14 word9_14 word8_14 R_wl
Cwl_9_14 word9_14 gnd C_wl
Rw10_14 word10_14 word9_14 R_wl
Cwl_10_14 word10_14 gnd C_wl
Rw11_14 word11_14 word10_14 R_wl
Cwl_11_14 word11_14 gnd C_wl
Rw12_14 word12_14 word11_14 R_wl
Cwl_12_14 word12_14 gnd C_wl
Rw13_14 word13_14 word12_14 R_wl
Cwl_13_14 word13_14 gnd C_wl
Rw14_14 word14_14 word13_14 R_wl
Cwl_14_14 word14_14 gnd C_wl
Rw15_14 word15_14 word14_14 R_wl
Cwl_15_14 word15_14 gnd C_wl
Rw16_14 word16_14 word15_14 R_wl
Cwl_16_14 word16_14 gnd C_wl
Rw17_14 word17_14 word16_14 R_wl
Cwl_17_14 word17_14 gnd C_wl
Rw18_14 word18_14 word17_14 R_wl
Cwl_18_14 word18_14 gnd C_wl
Rw19_14 word19_14 word18_14 R_wl
Cwl_19_14 word19_14 gnd C_wl
Rw20_14 word20_14 word19_14 R_wl
Cwl_20_14 word20_14 gnd C_wl
Rw21_14 word21_14 word20_14 R_wl
Cwl_21_14 word21_14 gnd C_wl
Rw22_14 word22_14 word21_14 R_wl
Cwl_22_14 word22_14 gnd C_wl
Rw23_14 word23_14 word22_14 R_wl
Cwl_23_14 word23_14 gnd C_wl
Rw24_14 word24_14 word23_14 R_wl
Cwl_24_14 word24_14 gnd C_wl
Rw25_14 word25_14 word24_14 R_wl
Cwl_25_14 word25_14 gnd C_wl
Rw26_14 word26_14 word25_14 R_wl
Cwl_26_14 word26_14 gnd C_wl
Rw27_14 word27_14 word26_14 R_wl
Cwl_27_14 word27_14 gnd C_wl
Rw28_14 word28_14 word27_14 R_wl
Cwl_28_14 word28_14 gnd C_wl
Rw29_14 word29_14 word28_14 R_wl
Cwl_29_14 word29_14 gnd C_wl
Rw30_14 word30_14 word29_14 R_wl
Cwl_30_14 word30_14 gnd C_wl
Rw31_14 word31_14 word30_14 R_wl
Cwl_31_14 word31_14 gnd C_wl
Rw32_14 word32_14 word31_14 R_wl
Cwl_32_14 word32_14 gnd C_wl
Rw33_14 word33_14 word32_14 R_wl
Cwl_33_14 word33_14 gnd C_wl
Rw34_14 word34_14 word33_14 R_wl
Cwl_34_14 word34_14 gnd C_wl
Rw35_14 word35_14 word34_14 R_wl
Cwl_35_14 word35_14 gnd C_wl
Rw36_14 word36_14 word35_14 R_wl
Cwl_36_14 word36_14 gnd C_wl
Rw37_14 word37_14 word36_14 R_wl
Cwl_37_14 word37_14 gnd C_wl
Rw38_14 word38_14 word37_14 R_wl
Cwl_38_14 word38_14 gnd C_wl
Rw39_14 word39_14 word38_14 R_wl
Cwl_39_14 word39_14 gnd C_wl
Rw40_14 word40_14 word39_14 R_wl
Cwl_40_14 word40_14 gnd C_wl
Rw41_14 word41_14 word40_14 R_wl
Cwl_41_14 word41_14 gnd C_wl
Rw42_14 word42_14 word41_14 R_wl
Cwl_42_14 word42_14 gnd C_wl
Rw43_14 word43_14 word42_14 R_wl
Cwl_43_14 word43_14 gnd C_wl
Rw44_14 word44_14 word43_14 R_wl
Cwl_44_14 word44_14 gnd C_wl
Rw45_14 word45_14 word44_14 R_wl
Cwl_45_14 word45_14 gnd C_wl
Rw46_14 word46_14 word45_14 R_wl
Cwl_46_14 word46_14 gnd C_wl
Rw47_14 word47_14 word46_14 R_wl
Cwl_47_14 word47_14 gnd C_wl
Rw48_14 word48_14 word47_14 R_wl
Cwl_48_14 word48_14 gnd C_wl
Rw49_14 word49_14 word48_14 R_wl
Cwl_49_14 word49_14 gnd C_wl
Rw50_14 word50_14 word49_14 R_wl
Cwl_50_14 word50_14 gnd C_wl
Rw51_14 word51_14 word50_14 R_wl
Cwl_51_14 word51_14 gnd C_wl
Rw52_14 word52_14 word51_14 R_wl
Cwl_52_14 word52_14 gnd C_wl
Rw53_14 word53_14 word52_14 R_wl
Cwl_53_14 word53_14 gnd C_wl
Rw54_14 word54_14 word53_14 R_wl
Cwl_54_14 word54_14 gnd C_wl
Rw55_14 word55_14 word54_14 R_wl
Cwl_55_14 word55_14 gnd C_wl
Rw56_14 word56_14 word55_14 R_wl
Cwl_56_14 word56_14 gnd C_wl
Rw57_14 word57_14 word56_14 R_wl
Cwl_57_14 word57_14 gnd C_wl
Rw58_14 word58_14 word57_14 R_wl
Cwl_58_14 word58_14 gnd C_wl
Rw59_14 word59_14 word58_14 R_wl
Cwl_59_14 word59_14 gnd C_wl
Rw60_14 word60_14 word59_14 R_wl
Cwl_60_14 word60_14 gnd C_wl
Rw61_14 word61_14 word60_14 R_wl
Cwl_61_14 word61_14 gnd C_wl
Rw62_14 word62_14 word61_14 R_wl
Cwl_62_14 word62_14 gnd C_wl
Rw63_14 word63_14 word62_14 R_wl
Cwl_63_14 word63_14 gnd C_wl
Rw64_14 word64_14 word63_14 R_wl
Cwl_64_14 word64_14 gnd C_wl
Rw65_14 word65_14 word64_14 R_wl
Cwl_65_14 word65_14 gnd C_wl
Rw66_14 word66_14 word65_14 R_wl
Cwl_66_14 word66_14 gnd C_wl
Rw67_14 word67_14 word66_14 R_wl
Cwl_67_14 word67_14 gnd C_wl
Rw68_14 word68_14 word67_14 R_wl
Cwl_68_14 word68_14 gnd C_wl
Rw69_14 word69_14 word68_14 R_wl
Cwl_69_14 word69_14 gnd C_wl
Rw70_14 word70_14 word69_14 R_wl
Cwl_70_14 word70_14 gnd C_wl
Rw71_14 word71_14 word70_14 R_wl
Cwl_71_14 word71_14 gnd C_wl
Rw72_14 word72_14 word71_14 R_wl
Cwl_72_14 word72_14 gnd C_wl
Rw73_14 word73_14 word72_14 R_wl
Cwl_73_14 word73_14 gnd C_wl
Rw74_14 word74_14 word73_14 R_wl
Cwl_74_14 word74_14 gnd C_wl
Rw75_14 word75_14 word74_14 R_wl
Cwl_75_14 word75_14 gnd C_wl
Rw76_14 word76_14 word75_14 R_wl
Cwl_76_14 word76_14 gnd C_wl
Rw77_14 word77_14 word76_14 R_wl
Cwl_77_14 word77_14 gnd C_wl
Rw78_14 word78_14 word77_14 R_wl
Cwl_78_14 word78_14 gnd C_wl
Rw79_14 word79_14 word78_14 R_wl
Cwl_79_14 word79_14 gnd C_wl
Rw80_14 word80_14 word79_14 R_wl
Cwl_80_14 word80_14 gnd C_wl
Rw81_14 word81_14 word80_14 R_wl
Cwl_81_14 word81_14 gnd C_wl
Rw82_14 word82_14 word81_14 R_wl
Cwl_82_14 word82_14 gnd C_wl
Rw83_14 word83_14 word82_14 R_wl
Cwl_83_14 word83_14 gnd C_wl
Rw84_14 word84_14 word83_14 R_wl
Cwl_84_14 word84_14 gnd C_wl
Rw85_14 word85_14 word84_14 R_wl
Cwl_85_14 word85_14 gnd C_wl
Rw86_14 word86_14 word85_14 R_wl
Cwl_86_14 word86_14 gnd C_wl
Rw87_14 word87_14 word86_14 R_wl
Cwl_87_14 word87_14 gnd C_wl
Rw88_14 word88_14 word87_14 R_wl
Cwl_88_14 word88_14 gnd C_wl
Rw89_14 word89_14 word88_14 R_wl
Cwl_89_14 word89_14 gnd C_wl
Rw90_14 word90_14 word89_14 R_wl
Cwl_90_14 word90_14 gnd C_wl
Rw91_14 word91_14 word90_14 R_wl
Cwl_91_14 word91_14 gnd C_wl
Rw92_14 word92_14 word91_14 R_wl
Cwl_92_14 word92_14 gnd C_wl
Rw93_14 word93_14 word92_14 R_wl
Cwl_93_14 word93_14 gnd C_wl
Rw94_14 word94_14 word93_14 R_wl
Cwl_94_14 word94_14 gnd C_wl
Rw95_14 word95_14 word94_14 R_wl
Cwl_95_14 word95_14 gnd C_wl
Rw96_14 word96_14 word95_14 R_wl
Cwl_96_14 word96_14 gnd C_wl
Rw97_14 word97_14 word96_14 R_wl
Cwl_97_14 word97_14 gnd C_wl
Rw98_14 word98_14 word97_14 R_wl
Cwl_98_14 word98_14 gnd C_wl
Rw99_14 word99_14 word98_14 R_wl
Cwl_99_14 word99_14 gnd C_wl
Vwl_15 word_15 0 0
Rw0_15 word_15 word0_15 R_wl
Cwl_0_15 word0_15 gnd C_wl
Rw1_15 word1_15 word0_15 R_wl
Cwl_1_15 word1_15 gnd C_wl
Rw2_15 word2_15 word1_15 R_wl
Cwl_2_15 word2_15 gnd C_wl
Rw3_15 word3_15 word2_15 R_wl
Cwl_3_15 word3_15 gnd C_wl
Rw4_15 word4_15 word3_15 R_wl
Cwl_4_15 word4_15 gnd C_wl
Rw5_15 word5_15 word4_15 R_wl
Cwl_5_15 word5_15 gnd C_wl
Rw6_15 word6_15 word5_15 R_wl
Cwl_6_15 word6_15 gnd C_wl
Rw7_15 word7_15 word6_15 R_wl
Cwl_7_15 word7_15 gnd C_wl
Rw8_15 word8_15 word7_15 R_wl
Cwl_8_15 word8_15 gnd C_wl
Rw9_15 word9_15 word8_15 R_wl
Cwl_9_15 word9_15 gnd C_wl
Rw10_15 word10_15 word9_15 R_wl
Cwl_10_15 word10_15 gnd C_wl
Rw11_15 word11_15 word10_15 R_wl
Cwl_11_15 word11_15 gnd C_wl
Rw12_15 word12_15 word11_15 R_wl
Cwl_12_15 word12_15 gnd C_wl
Rw13_15 word13_15 word12_15 R_wl
Cwl_13_15 word13_15 gnd C_wl
Rw14_15 word14_15 word13_15 R_wl
Cwl_14_15 word14_15 gnd C_wl
Rw15_15 word15_15 word14_15 R_wl
Cwl_15_15 word15_15 gnd C_wl
Rw16_15 word16_15 word15_15 R_wl
Cwl_16_15 word16_15 gnd C_wl
Rw17_15 word17_15 word16_15 R_wl
Cwl_17_15 word17_15 gnd C_wl
Rw18_15 word18_15 word17_15 R_wl
Cwl_18_15 word18_15 gnd C_wl
Rw19_15 word19_15 word18_15 R_wl
Cwl_19_15 word19_15 gnd C_wl
Rw20_15 word20_15 word19_15 R_wl
Cwl_20_15 word20_15 gnd C_wl
Rw21_15 word21_15 word20_15 R_wl
Cwl_21_15 word21_15 gnd C_wl
Rw22_15 word22_15 word21_15 R_wl
Cwl_22_15 word22_15 gnd C_wl
Rw23_15 word23_15 word22_15 R_wl
Cwl_23_15 word23_15 gnd C_wl
Rw24_15 word24_15 word23_15 R_wl
Cwl_24_15 word24_15 gnd C_wl
Rw25_15 word25_15 word24_15 R_wl
Cwl_25_15 word25_15 gnd C_wl
Rw26_15 word26_15 word25_15 R_wl
Cwl_26_15 word26_15 gnd C_wl
Rw27_15 word27_15 word26_15 R_wl
Cwl_27_15 word27_15 gnd C_wl
Rw28_15 word28_15 word27_15 R_wl
Cwl_28_15 word28_15 gnd C_wl
Rw29_15 word29_15 word28_15 R_wl
Cwl_29_15 word29_15 gnd C_wl
Rw30_15 word30_15 word29_15 R_wl
Cwl_30_15 word30_15 gnd C_wl
Rw31_15 word31_15 word30_15 R_wl
Cwl_31_15 word31_15 gnd C_wl
Rw32_15 word32_15 word31_15 R_wl
Cwl_32_15 word32_15 gnd C_wl
Rw33_15 word33_15 word32_15 R_wl
Cwl_33_15 word33_15 gnd C_wl
Rw34_15 word34_15 word33_15 R_wl
Cwl_34_15 word34_15 gnd C_wl
Rw35_15 word35_15 word34_15 R_wl
Cwl_35_15 word35_15 gnd C_wl
Rw36_15 word36_15 word35_15 R_wl
Cwl_36_15 word36_15 gnd C_wl
Rw37_15 word37_15 word36_15 R_wl
Cwl_37_15 word37_15 gnd C_wl
Rw38_15 word38_15 word37_15 R_wl
Cwl_38_15 word38_15 gnd C_wl
Rw39_15 word39_15 word38_15 R_wl
Cwl_39_15 word39_15 gnd C_wl
Rw40_15 word40_15 word39_15 R_wl
Cwl_40_15 word40_15 gnd C_wl
Rw41_15 word41_15 word40_15 R_wl
Cwl_41_15 word41_15 gnd C_wl
Rw42_15 word42_15 word41_15 R_wl
Cwl_42_15 word42_15 gnd C_wl
Rw43_15 word43_15 word42_15 R_wl
Cwl_43_15 word43_15 gnd C_wl
Rw44_15 word44_15 word43_15 R_wl
Cwl_44_15 word44_15 gnd C_wl
Rw45_15 word45_15 word44_15 R_wl
Cwl_45_15 word45_15 gnd C_wl
Rw46_15 word46_15 word45_15 R_wl
Cwl_46_15 word46_15 gnd C_wl
Rw47_15 word47_15 word46_15 R_wl
Cwl_47_15 word47_15 gnd C_wl
Rw48_15 word48_15 word47_15 R_wl
Cwl_48_15 word48_15 gnd C_wl
Rw49_15 word49_15 word48_15 R_wl
Cwl_49_15 word49_15 gnd C_wl
Rw50_15 word50_15 word49_15 R_wl
Cwl_50_15 word50_15 gnd C_wl
Rw51_15 word51_15 word50_15 R_wl
Cwl_51_15 word51_15 gnd C_wl
Rw52_15 word52_15 word51_15 R_wl
Cwl_52_15 word52_15 gnd C_wl
Rw53_15 word53_15 word52_15 R_wl
Cwl_53_15 word53_15 gnd C_wl
Rw54_15 word54_15 word53_15 R_wl
Cwl_54_15 word54_15 gnd C_wl
Rw55_15 word55_15 word54_15 R_wl
Cwl_55_15 word55_15 gnd C_wl
Rw56_15 word56_15 word55_15 R_wl
Cwl_56_15 word56_15 gnd C_wl
Rw57_15 word57_15 word56_15 R_wl
Cwl_57_15 word57_15 gnd C_wl
Rw58_15 word58_15 word57_15 R_wl
Cwl_58_15 word58_15 gnd C_wl
Rw59_15 word59_15 word58_15 R_wl
Cwl_59_15 word59_15 gnd C_wl
Rw60_15 word60_15 word59_15 R_wl
Cwl_60_15 word60_15 gnd C_wl
Rw61_15 word61_15 word60_15 R_wl
Cwl_61_15 word61_15 gnd C_wl
Rw62_15 word62_15 word61_15 R_wl
Cwl_62_15 word62_15 gnd C_wl
Rw63_15 word63_15 word62_15 R_wl
Cwl_63_15 word63_15 gnd C_wl
Rw64_15 word64_15 word63_15 R_wl
Cwl_64_15 word64_15 gnd C_wl
Rw65_15 word65_15 word64_15 R_wl
Cwl_65_15 word65_15 gnd C_wl
Rw66_15 word66_15 word65_15 R_wl
Cwl_66_15 word66_15 gnd C_wl
Rw67_15 word67_15 word66_15 R_wl
Cwl_67_15 word67_15 gnd C_wl
Rw68_15 word68_15 word67_15 R_wl
Cwl_68_15 word68_15 gnd C_wl
Rw69_15 word69_15 word68_15 R_wl
Cwl_69_15 word69_15 gnd C_wl
Rw70_15 word70_15 word69_15 R_wl
Cwl_70_15 word70_15 gnd C_wl
Rw71_15 word71_15 word70_15 R_wl
Cwl_71_15 word71_15 gnd C_wl
Rw72_15 word72_15 word71_15 R_wl
Cwl_72_15 word72_15 gnd C_wl
Rw73_15 word73_15 word72_15 R_wl
Cwl_73_15 word73_15 gnd C_wl
Rw74_15 word74_15 word73_15 R_wl
Cwl_74_15 word74_15 gnd C_wl
Rw75_15 word75_15 word74_15 R_wl
Cwl_75_15 word75_15 gnd C_wl
Rw76_15 word76_15 word75_15 R_wl
Cwl_76_15 word76_15 gnd C_wl
Rw77_15 word77_15 word76_15 R_wl
Cwl_77_15 word77_15 gnd C_wl
Rw78_15 word78_15 word77_15 R_wl
Cwl_78_15 word78_15 gnd C_wl
Rw79_15 word79_15 word78_15 R_wl
Cwl_79_15 word79_15 gnd C_wl
Rw80_15 word80_15 word79_15 R_wl
Cwl_80_15 word80_15 gnd C_wl
Rw81_15 word81_15 word80_15 R_wl
Cwl_81_15 word81_15 gnd C_wl
Rw82_15 word82_15 word81_15 R_wl
Cwl_82_15 word82_15 gnd C_wl
Rw83_15 word83_15 word82_15 R_wl
Cwl_83_15 word83_15 gnd C_wl
Rw84_15 word84_15 word83_15 R_wl
Cwl_84_15 word84_15 gnd C_wl
Rw85_15 word85_15 word84_15 R_wl
Cwl_85_15 word85_15 gnd C_wl
Rw86_15 word86_15 word85_15 R_wl
Cwl_86_15 word86_15 gnd C_wl
Rw87_15 word87_15 word86_15 R_wl
Cwl_87_15 word87_15 gnd C_wl
Rw88_15 word88_15 word87_15 R_wl
Cwl_88_15 word88_15 gnd C_wl
Rw89_15 word89_15 word88_15 R_wl
Cwl_89_15 word89_15 gnd C_wl
Rw90_15 word90_15 word89_15 R_wl
Cwl_90_15 word90_15 gnd C_wl
Rw91_15 word91_15 word90_15 R_wl
Cwl_91_15 word91_15 gnd C_wl
Rw92_15 word92_15 word91_15 R_wl
Cwl_92_15 word92_15 gnd C_wl
Rw93_15 word93_15 word92_15 R_wl
Cwl_93_15 word93_15 gnd C_wl
Rw94_15 word94_15 word93_15 R_wl
Cwl_94_15 word94_15 gnd C_wl
Rw95_15 word95_15 word94_15 R_wl
Cwl_95_15 word95_15 gnd C_wl
Rw96_15 word96_15 word95_15 R_wl
Cwl_96_15 word96_15 gnd C_wl
Rw97_15 word97_15 word96_15 R_wl
Cwl_97_15 word97_15 gnd C_wl
Rw98_15 word98_15 word97_15 R_wl
Cwl_98_15 word98_15 gnd C_wl
Rw99_15 word99_15 word98_15 R_wl
Cwl_99_15 word99_15 gnd C_wl
Vwl_16 word_16 0 0
Rw0_16 word_16 word0_16 R_wl
Cwl_0_16 word0_16 gnd C_wl
Rw1_16 word1_16 word0_16 R_wl
Cwl_1_16 word1_16 gnd C_wl
Rw2_16 word2_16 word1_16 R_wl
Cwl_2_16 word2_16 gnd C_wl
Rw3_16 word3_16 word2_16 R_wl
Cwl_3_16 word3_16 gnd C_wl
Rw4_16 word4_16 word3_16 R_wl
Cwl_4_16 word4_16 gnd C_wl
Rw5_16 word5_16 word4_16 R_wl
Cwl_5_16 word5_16 gnd C_wl
Rw6_16 word6_16 word5_16 R_wl
Cwl_6_16 word6_16 gnd C_wl
Rw7_16 word7_16 word6_16 R_wl
Cwl_7_16 word7_16 gnd C_wl
Rw8_16 word8_16 word7_16 R_wl
Cwl_8_16 word8_16 gnd C_wl
Rw9_16 word9_16 word8_16 R_wl
Cwl_9_16 word9_16 gnd C_wl
Rw10_16 word10_16 word9_16 R_wl
Cwl_10_16 word10_16 gnd C_wl
Rw11_16 word11_16 word10_16 R_wl
Cwl_11_16 word11_16 gnd C_wl
Rw12_16 word12_16 word11_16 R_wl
Cwl_12_16 word12_16 gnd C_wl
Rw13_16 word13_16 word12_16 R_wl
Cwl_13_16 word13_16 gnd C_wl
Rw14_16 word14_16 word13_16 R_wl
Cwl_14_16 word14_16 gnd C_wl
Rw15_16 word15_16 word14_16 R_wl
Cwl_15_16 word15_16 gnd C_wl
Rw16_16 word16_16 word15_16 R_wl
Cwl_16_16 word16_16 gnd C_wl
Rw17_16 word17_16 word16_16 R_wl
Cwl_17_16 word17_16 gnd C_wl
Rw18_16 word18_16 word17_16 R_wl
Cwl_18_16 word18_16 gnd C_wl
Rw19_16 word19_16 word18_16 R_wl
Cwl_19_16 word19_16 gnd C_wl
Rw20_16 word20_16 word19_16 R_wl
Cwl_20_16 word20_16 gnd C_wl
Rw21_16 word21_16 word20_16 R_wl
Cwl_21_16 word21_16 gnd C_wl
Rw22_16 word22_16 word21_16 R_wl
Cwl_22_16 word22_16 gnd C_wl
Rw23_16 word23_16 word22_16 R_wl
Cwl_23_16 word23_16 gnd C_wl
Rw24_16 word24_16 word23_16 R_wl
Cwl_24_16 word24_16 gnd C_wl
Rw25_16 word25_16 word24_16 R_wl
Cwl_25_16 word25_16 gnd C_wl
Rw26_16 word26_16 word25_16 R_wl
Cwl_26_16 word26_16 gnd C_wl
Rw27_16 word27_16 word26_16 R_wl
Cwl_27_16 word27_16 gnd C_wl
Rw28_16 word28_16 word27_16 R_wl
Cwl_28_16 word28_16 gnd C_wl
Rw29_16 word29_16 word28_16 R_wl
Cwl_29_16 word29_16 gnd C_wl
Rw30_16 word30_16 word29_16 R_wl
Cwl_30_16 word30_16 gnd C_wl
Rw31_16 word31_16 word30_16 R_wl
Cwl_31_16 word31_16 gnd C_wl
Rw32_16 word32_16 word31_16 R_wl
Cwl_32_16 word32_16 gnd C_wl
Rw33_16 word33_16 word32_16 R_wl
Cwl_33_16 word33_16 gnd C_wl
Rw34_16 word34_16 word33_16 R_wl
Cwl_34_16 word34_16 gnd C_wl
Rw35_16 word35_16 word34_16 R_wl
Cwl_35_16 word35_16 gnd C_wl
Rw36_16 word36_16 word35_16 R_wl
Cwl_36_16 word36_16 gnd C_wl
Rw37_16 word37_16 word36_16 R_wl
Cwl_37_16 word37_16 gnd C_wl
Rw38_16 word38_16 word37_16 R_wl
Cwl_38_16 word38_16 gnd C_wl
Rw39_16 word39_16 word38_16 R_wl
Cwl_39_16 word39_16 gnd C_wl
Rw40_16 word40_16 word39_16 R_wl
Cwl_40_16 word40_16 gnd C_wl
Rw41_16 word41_16 word40_16 R_wl
Cwl_41_16 word41_16 gnd C_wl
Rw42_16 word42_16 word41_16 R_wl
Cwl_42_16 word42_16 gnd C_wl
Rw43_16 word43_16 word42_16 R_wl
Cwl_43_16 word43_16 gnd C_wl
Rw44_16 word44_16 word43_16 R_wl
Cwl_44_16 word44_16 gnd C_wl
Rw45_16 word45_16 word44_16 R_wl
Cwl_45_16 word45_16 gnd C_wl
Rw46_16 word46_16 word45_16 R_wl
Cwl_46_16 word46_16 gnd C_wl
Rw47_16 word47_16 word46_16 R_wl
Cwl_47_16 word47_16 gnd C_wl
Rw48_16 word48_16 word47_16 R_wl
Cwl_48_16 word48_16 gnd C_wl
Rw49_16 word49_16 word48_16 R_wl
Cwl_49_16 word49_16 gnd C_wl
Rw50_16 word50_16 word49_16 R_wl
Cwl_50_16 word50_16 gnd C_wl
Rw51_16 word51_16 word50_16 R_wl
Cwl_51_16 word51_16 gnd C_wl
Rw52_16 word52_16 word51_16 R_wl
Cwl_52_16 word52_16 gnd C_wl
Rw53_16 word53_16 word52_16 R_wl
Cwl_53_16 word53_16 gnd C_wl
Rw54_16 word54_16 word53_16 R_wl
Cwl_54_16 word54_16 gnd C_wl
Rw55_16 word55_16 word54_16 R_wl
Cwl_55_16 word55_16 gnd C_wl
Rw56_16 word56_16 word55_16 R_wl
Cwl_56_16 word56_16 gnd C_wl
Rw57_16 word57_16 word56_16 R_wl
Cwl_57_16 word57_16 gnd C_wl
Rw58_16 word58_16 word57_16 R_wl
Cwl_58_16 word58_16 gnd C_wl
Rw59_16 word59_16 word58_16 R_wl
Cwl_59_16 word59_16 gnd C_wl
Rw60_16 word60_16 word59_16 R_wl
Cwl_60_16 word60_16 gnd C_wl
Rw61_16 word61_16 word60_16 R_wl
Cwl_61_16 word61_16 gnd C_wl
Rw62_16 word62_16 word61_16 R_wl
Cwl_62_16 word62_16 gnd C_wl
Rw63_16 word63_16 word62_16 R_wl
Cwl_63_16 word63_16 gnd C_wl
Rw64_16 word64_16 word63_16 R_wl
Cwl_64_16 word64_16 gnd C_wl
Rw65_16 word65_16 word64_16 R_wl
Cwl_65_16 word65_16 gnd C_wl
Rw66_16 word66_16 word65_16 R_wl
Cwl_66_16 word66_16 gnd C_wl
Rw67_16 word67_16 word66_16 R_wl
Cwl_67_16 word67_16 gnd C_wl
Rw68_16 word68_16 word67_16 R_wl
Cwl_68_16 word68_16 gnd C_wl
Rw69_16 word69_16 word68_16 R_wl
Cwl_69_16 word69_16 gnd C_wl
Rw70_16 word70_16 word69_16 R_wl
Cwl_70_16 word70_16 gnd C_wl
Rw71_16 word71_16 word70_16 R_wl
Cwl_71_16 word71_16 gnd C_wl
Rw72_16 word72_16 word71_16 R_wl
Cwl_72_16 word72_16 gnd C_wl
Rw73_16 word73_16 word72_16 R_wl
Cwl_73_16 word73_16 gnd C_wl
Rw74_16 word74_16 word73_16 R_wl
Cwl_74_16 word74_16 gnd C_wl
Rw75_16 word75_16 word74_16 R_wl
Cwl_75_16 word75_16 gnd C_wl
Rw76_16 word76_16 word75_16 R_wl
Cwl_76_16 word76_16 gnd C_wl
Rw77_16 word77_16 word76_16 R_wl
Cwl_77_16 word77_16 gnd C_wl
Rw78_16 word78_16 word77_16 R_wl
Cwl_78_16 word78_16 gnd C_wl
Rw79_16 word79_16 word78_16 R_wl
Cwl_79_16 word79_16 gnd C_wl
Rw80_16 word80_16 word79_16 R_wl
Cwl_80_16 word80_16 gnd C_wl
Rw81_16 word81_16 word80_16 R_wl
Cwl_81_16 word81_16 gnd C_wl
Rw82_16 word82_16 word81_16 R_wl
Cwl_82_16 word82_16 gnd C_wl
Rw83_16 word83_16 word82_16 R_wl
Cwl_83_16 word83_16 gnd C_wl
Rw84_16 word84_16 word83_16 R_wl
Cwl_84_16 word84_16 gnd C_wl
Rw85_16 word85_16 word84_16 R_wl
Cwl_85_16 word85_16 gnd C_wl
Rw86_16 word86_16 word85_16 R_wl
Cwl_86_16 word86_16 gnd C_wl
Rw87_16 word87_16 word86_16 R_wl
Cwl_87_16 word87_16 gnd C_wl
Rw88_16 word88_16 word87_16 R_wl
Cwl_88_16 word88_16 gnd C_wl
Rw89_16 word89_16 word88_16 R_wl
Cwl_89_16 word89_16 gnd C_wl
Rw90_16 word90_16 word89_16 R_wl
Cwl_90_16 word90_16 gnd C_wl
Rw91_16 word91_16 word90_16 R_wl
Cwl_91_16 word91_16 gnd C_wl
Rw92_16 word92_16 word91_16 R_wl
Cwl_92_16 word92_16 gnd C_wl
Rw93_16 word93_16 word92_16 R_wl
Cwl_93_16 word93_16 gnd C_wl
Rw94_16 word94_16 word93_16 R_wl
Cwl_94_16 word94_16 gnd C_wl
Rw95_16 word95_16 word94_16 R_wl
Cwl_95_16 word95_16 gnd C_wl
Rw96_16 word96_16 word95_16 R_wl
Cwl_96_16 word96_16 gnd C_wl
Rw97_16 word97_16 word96_16 R_wl
Cwl_97_16 word97_16 gnd C_wl
Rw98_16 word98_16 word97_16 R_wl
Cwl_98_16 word98_16 gnd C_wl
Rw99_16 word99_16 word98_16 R_wl
Cwl_99_16 word99_16 gnd C_wl
Vwl_17 word_17 0 0
Rw0_17 word_17 word0_17 R_wl
Cwl_0_17 word0_17 gnd C_wl
Rw1_17 word1_17 word0_17 R_wl
Cwl_1_17 word1_17 gnd C_wl
Rw2_17 word2_17 word1_17 R_wl
Cwl_2_17 word2_17 gnd C_wl
Rw3_17 word3_17 word2_17 R_wl
Cwl_3_17 word3_17 gnd C_wl
Rw4_17 word4_17 word3_17 R_wl
Cwl_4_17 word4_17 gnd C_wl
Rw5_17 word5_17 word4_17 R_wl
Cwl_5_17 word5_17 gnd C_wl
Rw6_17 word6_17 word5_17 R_wl
Cwl_6_17 word6_17 gnd C_wl
Rw7_17 word7_17 word6_17 R_wl
Cwl_7_17 word7_17 gnd C_wl
Rw8_17 word8_17 word7_17 R_wl
Cwl_8_17 word8_17 gnd C_wl
Rw9_17 word9_17 word8_17 R_wl
Cwl_9_17 word9_17 gnd C_wl
Rw10_17 word10_17 word9_17 R_wl
Cwl_10_17 word10_17 gnd C_wl
Rw11_17 word11_17 word10_17 R_wl
Cwl_11_17 word11_17 gnd C_wl
Rw12_17 word12_17 word11_17 R_wl
Cwl_12_17 word12_17 gnd C_wl
Rw13_17 word13_17 word12_17 R_wl
Cwl_13_17 word13_17 gnd C_wl
Rw14_17 word14_17 word13_17 R_wl
Cwl_14_17 word14_17 gnd C_wl
Rw15_17 word15_17 word14_17 R_wl
Cwl_15_17 word15_17 gnd C_wl
Rw16_17 word16_17 word15_17 R_wl
Cwl_16_17 word16_17 gnd C_wl
Rw17_17 word17_17 word16_17 R_wl
Cwl_17_17 word17_17 gnd C_wl
Rw18_17 word18_17 word17_17 R_wl
Cwl_18_17 word18_17 gnd C_wl
Rw19_17 word19_17 word18_17 R_wl
Cwl_19_17 word19_17 gnd C_wl
Rw20_17 word20_17 word19_17 R_wl
Cwl_20_17 word20_17 gnd C_wl
Rw21_17 word21_17 word20_17 R_wl
Cwl_21_17 word21_17 gnd C_wl
Rw22_17 word22_17 word21_17 R_wl
Cwl_22_17 word22_17 gnd C_wl
Rw23_17 word23_17 word22_17 R_wl
Cwl_23_17 word23_17 gnd C_wl
Rw24_17 word24_17 word23_17 R_wl
Cwl_24_17 word24_17 gnd C_wl
Rw25_17 word25_17 word24_17 R_wl
Cwl_25_17 word25_17 gnd C_wl
Rw26_17 word26_17 word25_17 R_wl
Cwl_26_17 word26_17 gnd C_wl
Rw27_17 word27_17 word26_17 R_wl
Cwl_27_17 word27_17 gnd C_wl
Rw28_17 word28_17 word27_17 R_wl
Cwl_28_17 word28_17 gnd C_wl
Rw29_17 word29_17 word28_17 R_wl
Cwl_29_17 word29_17 gnd C_wl
Rw30_17 word30_17 word29_17 R_wl
Cwl_30_17 word30_17 gnd C_wl
Rw31_17 word31_17 word30_17 R_wl
Cwl_31_17 word31_17 gnd C_wl
Rw32_17 word32_17 word31_17 R_wl
Cwl_32_17 word32_17 gnd C_wl
Rw33_17 word33_17 word32_17 R_wl
Cwl_33_17 word33_17 gnd C_wl
Rw34_17 word34_17 word33_17 R_wl
Cwl_34_17 word34_17 gnd C_wl
Rw35_17 word35_17 word34_17 R_wl
Cwl_35_17 word35_17 gnd C_wl
Rw36_17 word36_17 word35_17 R_wl
Cwl_36_17 word36_17 gnd C_wl
Rw37_17 word37_17 word36_17 R_wl
Cwl_37_17 word37_17 gnd C_wl
Rw38_17 word38_17 word37_17 R_wl
Cwl_38_17 word38_17 gnd C_wl
Rw39_17 word39_17 word38_17 R_wl
Cwl_39_17 word39_17 gnd C_wl
Rw40_17 word40_17 word39_17 R_wl
Cwl_40_17 word40_17 gnd C_wl
Rw41_17 word41_17 word40_17 R_wl
Cwl_41_17 word41_17 gnd C_wl
Rw42_17 word42_17 word41_17 R_wl
Cwl_42_17 word42_17 gnd C_wl
Rw43_17 word43_17 word42_17 R_wl
Cwl_43_17 word43_17 gnd C_wl
Rw44_17 word44_17 word43_17 R_wl
Cwl_44_17 word44_17 gnd C_wl
Rw45_17 word45_17 word44_17 R_wl
Cwl_45_17 word45_17 gnd C_wl
Rw46_17 word46_17 word45_17 R_wl
Cwl_46_17 word46_17 gnd C_wl
Rw47_17 word47_17 word46_17 R_wl
Cwl_47_17 word47_17 gnd C_wl
Rw48_17 word48_17 word47_17 R_wl
Cwl_48_17 word48_17 gnd C_wl
Rw49_17 word49_17 word48_17 R_wl
Cwl_49_17 word49_17 gnd C_wl
Rw50_17 word50_17 word49_17 R_wl
Cwl_50_17 word50_17 gnd C_wl
Rw51_17 word51_17 word50_17 R_wl
Cwl_51_17 word51_17 gnd C_wl
Rw52_17 word52_17 word51_17 R_wl
Cwl_52_17 word52_17 gnd C_wl
Rw53_17 word53_17 word52_17 R_wl
Cwl_53_17 word53_17 gnd C_wl
Rw54_17 word54_17 word53_17 R_wl
Cwl_54_17 word54_17 gnd C_wl
Rw55_17 word55_17 word54_17 R_wl
Cwl_55_17 word55_17 gnd C_wl
Rw56_17 word56_17 word55_17 R_wl
Cwl_56_17 word56_17 gnd C_wl
Rw57_17 word57_17 word56_17 R_wl
Cwl_57_17 word57_17 gnd C_wl
Rw58_17 word58_17 word57_17 R_wl
Cwl_58_17 word58_17 gnd C_wl
Rw59_17 word59_17 word58_17 R_wl
Cwl_59_17 word59_17 gnd C_wl
Rw60_17 word60_17 word59_17 R_wl
Cwl_60_17 word60_17 gnd C_wl
Rw61_17 word61_17 word60_17 R_wl
Cwl_61_17 word61_17 gnd C_wl
Rw62_17 word62_17 word61_17 R_wl
Cwl_62_17 word62_17 gnd C_wl
Rw63_17 word63_17 word62_17 R_wl
Cwl_63_17 word63_17 gnd C_wl
Rw64_17 word64_17 word63_17 R_wl
Cwl_64_17 word64_17 gnd C_wl
Rw65_17 word65_17 word64_17 R_wl
Cwl_65_17 word65_17 gnd C_wl
Rw66_17 word66_17 word65_17 R_wl
Cwl_66_17 word66_17 gnd C_wl
Rw67_17 word67_17 word66_17 R_wl
Cwl_67_17 word67_17 gnd C_wl
Rw68_17 word68_17 word67_17 R_wl
Cwl_68_17 word68_17 gnd C_wl
Rw69_17 word69_17 word68_17 R_wl
Cwl_69_17 word69_17 gnd C_wl
Rw70_17 word70_17 word69_17 R_wl
Cwl_70_17 word70_17 gnd C_wl
Rw71_17 word71_17 word70_17 R_wl
Cwl_71_17 word71_17 gnd C_wl
Rw72_17 word72_17 word71_17 R_wl
Cwl_72_17 word72_17 gnd C_wl
Rw73_17 word73_17 word72_17 R_wl
Cwl_73_17 word73_17 gnd C_wl
Rw74_17 word74_17 word73_17 R_wl
Cwl_74_17 word74_17 gnd C_wl
Rw75_17 word75_17 word74_17 R_wl
Cwl_75_17 word75_17 gnd C_wl
Rw76_17 word76_17 word75_17 R_wl
Cwl_76_17 word76_17 gnd C_wl
Rw77_17 word77_17 word76_17 R_wl
Cwl_77_17 word77_17 gnd C_wl
Rw78_17 word78_17 word77_17 R_wl
Cwl_78_17 word78_17 gnd C_wl
Rw79_17 word79_17 word78_17 R_wl
Cwl_79_17 word79_17 gnd C_wl
Rw80_17 word80_17 word79_17 R_wl
Cwl_80_17 word80_17 gnd C_wl
Rw81_17 word81_17 word80_17 R_wl
Cwl_81_17 word81_17 gnd C_wl
Rw82_17 word82_17 word81_17 R_wl
Cwl_82_17 word82_17 gnd C_wl
Rw83_17 word83_17 word82_17 R_wl
Cwl_83_17 word83_17 gnd C_wl
Rw84_17 word84_17 word83_17 R_wl
Cwl_84_17 word84_17 gnd C_wl
Rw85_17 word85_17 word84_17 R_wl
Cwl_85_17 word85_17 gnd C_wl
Rw86_17 word86_17 word85_17 R_wl
Cwl_86_17 word86_17 gnd C_wl
Rw87_17 word87_17 word86_17 R_wl
Cwl_87_17 word87_17 gnd C_wl
Rw88_17 word88_17 word87_17 R_wl
Cwl_88_17 word88_17 gnd C_wl
Rw89_17 word89_17 word88_17 R_wl
Cwl_89_17 word89_17 gnd C_wl
Rw90_17 word90_17 word89_17 R_wl
Cwl_90_17 word90_17 gnd C_wl
Rw91_17 word91_17 word90_17 R_wl
Cwl_91_17 word91_17 gnd C_wl
Rw92_17 word92_17 word91_17 R_wl
Cwl_92_17 word92_17 gnd C_wl
Rw93_17 word93_17 word92_17 R_wl
Cwl_93_17 word93_17 gnd C_wl
Rw94_17 word94_17 word93_17 R_wl
Cwl_94_17 word94_17 gnd C_wl
Rw95_17 word95_17 word94_17 R_wl
Cwl_95_17 word95_17 gnd C_wl
Rw96_17 word96_17 word95_17 R_wl
Cwl_96_17 word96_17 gnd C_wl
Rw97_17 word97_17 word96_17 R_wl
Cwl_97_17 word97_17 gnd C_wl
Rw98_17 word98_17 word97_17 R_wl
Cwl_98_17 word98_17 gnd C_wl
Rw99_17 word99_17 word98_17 R_wl
Cwl_99_17 word99_17 gnd C_wl
Vwl_18 word_18 0 0
Rw0_18 word_18 word0_18 R_wl
Cwl_0_18 word0_18 gnd C_wl
Rw1_18 word1_18 word0_18 R_wl
Cwl_1_18 word1_18 gnd C_wl
Rw2_18 word2_18 word1_18 R_wl
Cwl_2_18 word2_18 gnd C_wl
Rw3_18 word3_18 word2_18 R_wl
Cwl_3_18 word3_18 gnd C_wl
Rw4_18 word4_18 word3_18 R_wl
Cwl_4_18 word4_18 gnd C_wl
Rw5_18 word5_18 word4_18 R_wl
Cwl_5_18 word5_18 gnd C_wl
Rw6_18 word6_18 word5_18 R_wl
Cwl_6_18 word6_18 gnd C_wl
Rw7_18 word7_18 word6_18 R_wl
Cwl_7_18 word7_18 gnd C_wl
Rw8_18 word8_18 word7_18 R_wl
Cwl_8_18 word8_18 gnd C_wl
Rw9_18 word9_18 word8_18 R_wl
Cwl_9_18 word9_18 gnd C_wl
Rw10_18 word10_18 word9_18 R_wl
Cwl_10_18 word10_18 gnd C_wl
Rw11_18 word11_18 word10_18 R_wl
Cwl_11_18 word11_18 gnd C_wl
Rw12_18 word12_18 word11_18 R_wl
Cwl_12_18 word12_18 gnd C_wl
Rw13_18 word13_18 word12_18 R_wl
Cwl_13_18 word13_18 gnd C_wl
Rw14_18 word14_18 word13_18 R_wl
Cwl_14_18 word14_18 gnd C_wl
Rw15_18 word15_18 word14_18 R_wl
Cwl_15_18 word15_18 gnd C_wl
Rw16_18 word16_18 word15_18 R_wl
Cwl_16_18 word16_18 gnd C_wl
Rw17_18 word17_18 word16_18 R_wl
Cwl_17_18 word17_18 gnd C_wl
Rw18_18 word18_18 word17_18 R_wl
Cwl_18_18 word18_18 gnd C_wl
Rw19_18 word19_18 word18_18 R_wl
Cwl_19_18 word19_18 gnd C_wl
Rw20_18 word20_18 word19_18 R_wl
Cwl_20_18 word20_18 gnd C_wl
Rw21_18 word21_18 word20_18 R_wl
Cwl_21_18 word21_18 gnd C_wl
Rw22_18 word22_18 word21_18 R_wl
Cwl_22_18 word22_18 gnd C_wl
Rw23_18 word23_18 word22_18 R_wl
Cwl_23_18 word23_18 gnd C_wl
Rw24_18 word24_18 word23_18 R_wl
Cwl_24_18 word24_18 gnd C_wl
Rw25_18 word25_18 word24_18 R_wl
Cwl_25_18 word25_18 gnd C_wl
Rw26_18 word26_18 word25_18 R_wl
Cwl_26_18 word26_18 gnd C_wl
Rw27_18 word27_18 word26_18 R_wl
Cwl_27_18 word27_18 gnd C_wl
Rw28_18 word28_18 word27_18 R_wl
Cwl_28_18 word28_18 gnd C_wl
Rw29_18 word29_18 word28_18 R_wl
Cwl_29_18 word29_18 gnd C_wl
Rw30_18 word30_18 word29_18 R_wl
Cwl_30_18 word30_18 gnd C_wl
Rw31_18 word31_18 word30_18 R_wl
Cwl_31_18 word31_18 gnd C_wl
Rw32_18 word32_18 word31_18 R_wl
Cwl_32_18 word32_18 gnd C_wl
Rw33_18 word33_18 word32_18 R_wl
Cwl_33_18 word33_18 gnd C_wl
Rw34_18 word34_18 word33_18 R_wl
Cwl_34_18 word34_18 gnd C_wl
Rw35_18 word35_18 word34_18 R_wl
Cwl_35_18 word35_18 gnd C_wl
Rw36_18 word36_18 word35_18 R_wl
Cwl_36_18 word36_18 gnd C_wl
Rw37_18 word37_18 word36_18 R_wl
Cwl_37_18 word37_18 gnd C_wl
Rw38_18 word38_18 word37_18 R_wl
Cwl_38_18 word38_18 gnd C_wl
Rw39_18 word39_18 word38_18 R_wl
Cwl_39_18 word39_18 gnd C_wl
Rw40_18 word40_18 word39_18 R_wl
Cwl_40_18 word40_18 gnd C_wl
Rw41_18 word41_18 word40_18 R_wl
Cwl_41_18 word41_18 gnd C_wl
Rw42_18 word42_18 word41_18 R_wl
Cwl_42_18 word42_18 gnd C_wl
Rw43_18 word43_18 word42_18 R_wl
Cwl_43_18 word43_18 gnd C_wl
Rw44_18 word44_18 word43_18 R_wl
Cwl_44_18 word44_18 gnd C_wl
Rw45_18 word45_18 word44_18 R_wl
Cwl_45_18 word45_18 gnd C_wl
Rw46_18 word46_18 word45_18 R_wl
Cwl_46_18 word46_18 gnd C_wl
Rw47_18 word47_18 word46_18 R_wl
Cwl_47_18 word47_18 gnd C_wl
Rw48_18 word48_18 word47_18 R_wl
Cwl_48_18 word48_18 gnd C_wl
Rw49_18 word49_18 word48_18 R_wl
Cwl_49_18 word49_18 gnd C_wl
Rw50_18 word50_18 word49_18 R_wl
Cwl_50_18 word50_18 gnd C_wl
Rw51_18 word51_18 word50_18 R_wl
Cwl_51_18 word51_18 gnd C_wl
Rw52_18 word52_18 word51_18 R_wl
Cwl_52_18 word52_18 gnd C_wl
Rw53_18 word53_18 word52_18 R_wl
Cwl_53_18 word53_18 gnd C_wl
Rw54_18 word54_18 word53_18 R_wl
Cwl_54_18 word54_18 gnd C_wl
Rw55_18 word55_18 word54_18 R_wl
Cwl_55_18 word55_18 gnd C_wl
Rw56_18 word56_18 word55_18 R_wl
Cwl_56_18 word56_18 gnd C_wl
Rw57_18 word57_18 word56_18 R_wl
Cwl_57_18 word57_18 gnd C_wl
Rw58_18 word58_18 word57_18 R_wl
Cwl_58_18 word58_18 gnd C_wl
Rw59_18 word59_18 word58_18 R_wl
Cwl_59_18 word59_18 gnd C_wl
Rw60_18 word60_18 word59_18 R_wl
Cwl_60_18 word60_18 gnd C_wl
Rw61_18 word61_18 word60_18 R_wl
Cwl_61_18 word61_18 gnd C_wl
Rw62_18 word62_18 word61_18 R_wl
Cwl_62_18 word62_18 gnd C_wl
Rw63_18 word63_18 word62_18 R_wl
Cwl_63_18 word63_18 gnd C_wl
Rw64_18 word64_18 word63_18 R_wl
Cwl_64_18 word64_18 gnd C_wl
Rw65_18 word65_18 word64_18 R_wl
Cwl_65_18 word65_18 gnd C_wl
Rw66_18 word66_18 word65_18 R_wl
Cwl_66_18 word66_18 gnd C_wl
Rw67_18 word67_18 word66_18 R_wl
Cwl_67_18 word67_18 gnd C_wl
Rw68_18 word68_18 word67_18 R_wl
Cwl_68_18 word68_18 gnd C_wl
Rw69_18 word69_18 word68_18 R_wl
Cwl_69_18 word69_18 gnd C_wl
Rw70_18 word70_18 word69_18 R_wl
Cwl_70_18 word70_18 gnd C_wl
Rw71_18 word71_18 word70_18 R_wl
Cwl_71_18 word71_18 gnd C_wl
Rw72_18 word72_18 word71_18 R_wl
Cwl_72_18 word72_18 gnd C_wl
Rw73_18 word73_18 word72_18 R_wl
Cwl_73_18 word73_18 gnd C_wl
Rw74_18 word74_18 word73_18 R_wl
Cwl_74_18 word74_18 gnd C_wl
Rw75_18 word75_18 word74_18 R_wl
Cwl_75_18 word75_18 gnd C_wl
Rw76_18 word76_18 word75_18 R_wl
Cwl_76_18 word76_18 gnd C_wl
Rw77_18 word77_18 word76_18 R_wl
Cwl_77_18 word77_18 gnd C_wl
Rw78_18 word78_18 word77_18 R_wl
Cwl_78_18 word78_18 gnd C_wl
Rw79_18 word79_18 word78_18 R_wl
Cwl_79_18 word79_18 gnd C_wl
Rw80_18 word80_18 word79_18 R_wl
Cwl_80_18 word80_18 gnd C_wl
Rw81_18 word81_18 word80_18 R_wl
Cwl_81_18 word81_18 gnd C_wl
Rw82_18 word82_18 word81_18 R_wl
Cwl_82_18 word82_18 gnd C_wl
Rw83_18 word83_18 word82_18 R_wl
Cwl_83_18 word83_18 gnd C_wl
Rw84_18 word84_18 word83_18 R_wl
Cwl_84_18 word84_18 gnd C_wl
Rw85_18 word85_18 word84_18 R_wl
Cwl_85_18 word85_18 gnd C_wl
Rw86_18 word86_18 word85_18 R_wl
Cwl_86_18 word86_18 gnd C_wl
Rw87_18 word87_18 word86_18 R_wl
Cwl_87_18 word87_18 gnd C_wl
Rw88_18 word88_18 word87_18 R_wl
Cwl_88_18 word88_18 gnd C_wl
Rw89_18 word89_18 word88_18 R_wl
Cwl_89_18 word89_18 gnd C_wl
Rw90_18 word90_18 word89_18 R_wl
Cwl_90_18 word90_18 gnd C_wl
Rw91_18 word91_18 word90_18 R_wl
Cwl_91_18 word91_18 gnd C_wl
Rw92_18 word92_18 word91_18 R_wl
Cwl_92_18 word92_18 gnd C_wl
Rw93_18 word93_18 word92_18 R_wl
Cwl_93_18 word93_18 gnd C_wl
Rw94_18 word94_18 word93_18 R_wl
Cwl_94_18 word94_18 gnd C_wl
Rw95_18 word95_18 word94_18 R_wl
Cwl_95_18 word95_18 gnd C_wl
Rw96_18 word96_18 word95_18 R_wl
Cwl_96_18 word96_18 gnd C_wl
Rw97_18 word97_18 word96_18 R_wl
Cwl_97_18 word97_18 gnd C_wl
Rw98_18 word98_18 word97_18 R_wl
Cwl_98_18 word98_18 gnd C_wl
Rw99_18 word99_18 word98_18 R_wl
Cwl_99_18 word99_18 gnd C_wl
Vwl_19 word_19 0 0
Rw0_19 word_19 word0_19 R_wl
Cwl_0_19 word0_19 gnd C_wl
Rw1_19 word1_19 word0_19 R_wl
Cwl_1_19 word1_19 gnd C_wl
Rw2_19 word2_19 word1_19 R_wl
Cwl_2_19 word2_19 gnd C_wl
Rw3_19 word3_19 word2_19 R_wl
Cwl_3_19 word3_19 gnd C_wl
Rw4_19 word4_19 word3_19 R_wl
Cwl_4_19 word4_19 gnd C_wl
Rw5_19 word5_19 word4_19 R_wl
Cwl_5_19 word5_19 gnd C_wl
Rw6_19 word6_19 word5_19 R_wl
Cwl_6_19 word6_19 gnd C_wl
Rw7_19 word7_19 word6_19 R_wl
Cwl_7_19 word7_19 gnd C_wl
Rw8_19 word8_19 word7_19 R_wl
Cwl_8_19 word8_19 gnd C_wl
Rw9_19 word9_19 word8_19 R_wl
Cwl_9_19 word9_19 gnd C_wl
Rw10_19 word10_19 word9_19 R_wl
Cwl_10_19 word10_19 gnd C_wl
Rw11_19 word11_19 word10_19 R_wl
Cwl_11_19 word11_19 gnd C_wl
Rw12_19 word12_19 word11_19 R_wl
Cwl_12_19 word12_19 gnd C_wl
Rw13_19 word13_19 word12_19 R_wl
Cwl_13_19 word13_19 gnd C_wl
Rw14_19 word14_19 word13_19 R_wl
Cwl_14_19 word14_19 gnd C_wl
Rw15_19 word15_19 word14_19 R_wl
Cwl_15_19 word15_19 gnd C_wl
Rw16_19 word16_19 word15_19 R_wl
Cwl_16_19 word16_19 gnd C_wl
Rw17_19 word17_19 word16_19 R_wl
Cwl_17_19 word17_19 gnd C_wl
Rw18_19 word18_19 word17_19 R_wl
Cwl_18_19 word18_19 gnd C_wl
Rw19_19 word19_19 word18_19 R_wl
Cwl_19_19 word19_19 gnd C_wl
Rw20_19 word20_19 word19_19 R_wl
Cwl_20_19 word20_19 gnd C_wl
Rw21_19 word21_19 word20_19 R_wl
Cwl_21_19 word21_19 gnd C_wl
Rw22_19 word22_19 word21_19 R_wl
Cwl_22_19 word22_19 gnd C_wl
Rw23_19 word23_19 word22_19 R_wl
Cwl_23_19 word23_19 gnd C_wl
Rw24_19 word24_19 word23_19 R_wl
Cwl_24_19 word24_19 gnd C_wl
Rw25_19 word25_19 word24_19 R_wl
Cwl_25_19 word25_19 gnd C_wl
Rw26_19 word26_19 word25_19 R_wl
Cwl_26_19 word26_19 gnd C_wl
Rw27_19 word27_19 word26_19 R_wl
Cwl_27_19 word27_19 gnd C_wl
Rw28_19 word28_19 word27_19 R_wl
Cwl_28_19 word28_19 gnd C_wl
Rw29_19 word29_19 word28_19 R_wl
Cwl_29_19 word29_19 gnd C_wl
Rw30_19 word30_19 word29_19 R_wl
Cwl_30_19 word30_19 gnd C_wl
Rw31_19 word31_19 word30_19 R_wl
Cwl_31_19 word31_19 gnd C_wl
Rw32_19 word32_19 word31_19 R_wl
Cwl_32_19 word32_19 gnd C_wl
Rw33_19 word33_19 word32_19 R_wl
Cwl_33_19 word33_19 gnd C_wl
Rw34_19 word34_19 word33_19 R_wl
Cwl_34_19 word34_19 gnd C_wl
Rw35_19 word35_19 word34_19 R_wl
Cwl_35_19 word35_19 gnd C_wl
Rw36_19 word36_19 word35_19 R_wl
Cwl_36_19 word36_19 gnd C_wl
Rw37_19 word37_19 word36_19 R_wl
Cwl_37_19 word37_19 gnd C_wl
Rw38_19 word38_19 word37_19 R_wl
Cwl_38_19 word38_19 gnd C_wl
Rw39_19 word39_19 word38_19 R_wl
Cwl_39_19 word39_19 gnd C_wl
Rw40_19 word40_19 word39_19 R_wl
Cwl_40_19 word40_19 gnd C_wl
Rw41_19 word41_19 word40_19 R_wl
Cwl_41_19 word41_19 gnd C_wl
Rw42_19 word42_19 word41_19 R_wl
Cwl_42_19 word42_19 gnd C_wl
Rw43_19 word43_19 word42_19 R_wl
Cwl_43_19 word43_19 gnd C_wl
Rw44_19 word44_19 word43_19 R_wl
Cwl_44_19 word44_19 gnd C_wl
Rw45_19 word45_19 word44_19 R_wl
Cwl_45_19 word45_19 gnd C_wl
Rw46_19 word46_19 word45_19 R_wl
Cwl_46_19 word46_19 gnd C_wl
Rw47_19 word47_19 word46_19 R_wl
Cwl_47_19 word47_19 gnd C_wl
Rw48_19 word48_19 word47_19 R_wl
Cwl_48_19 word48_19 gnd C_wl
Rw49_19 word49_19 word48_19 R_wl
Cwl_49_19 word49_19 gnd C_wl
Rw50_19 word50_19 word49_19 R_wl
Cwl_50_19 word50_19 gnd C_wl
Rw51_19 word51_19 word50_19 R_wl
Cwl_51_19 word51_19 gnd C_wl
Rw52_19 word52_19 word51_19 R_wl
Cwl_52_19 word52_19 gnd C_wl
Rw53_19 word53_19 word52_19 R_wl
Cwl_53_19 word53_19 gnd C_wl
Rw54_19 word54_19 word53_19 R_wl
Cwl_54_19 word54_19 gnd C_wl
Rw55_19 word55_19 word54_19 R_wl
Cwl_55_19 word55_19 gnd C_wl
Rw56_19 word56_19 word55_19 R_wl
Cwl_56_19 word56_19 gnd C_wl
Rw57_19 word57_19 word56_19 R_wl
Cwl_57_19 word57_19 gnd C_wl
Rw58_19 word58_19 word57_19 R_wl
Cwl_58_19 word58_19 gnd C_wl
Rw59_19 word59_19 word58_19 R_wl
Cwl_59_19 word59_19 gnd C_wl
Rw60_19 word60_19 word59_19 R_wl
Cwl_60_19 word60_19 gnd C_wl
Rw61_19 word61_19 word60_19 R_wl
Cwl_61_19 word61_19 gnd C_wl
Rw62_19 word62_19 word61_19 R_wl
Cwl_62_19 word62_19 gnd C_wl
Rw63_19 word63_19 word62_19 R_wl
Cwl_63_19 word63_19 gnd C_wl
Rw64_19 word64_19 word63_19 R_wl
Cwl_64_19 word64_19 gnd C_wl
Rw65_19 word65_19 word64_19 R_wl
Cwl_65_19 word65_19 gnd C_wl
Rw66_19 word66_19 word65_19 R_wl
Cwl_66_19 word66_19 gnd C_wl
Rw67_19 word67_19 word66_19 R_wl
Cwl_67_19 word67_19 gnd C_wl
Rw68_19 word68_19 word67_19 R_wl
Cwl_68_19 word68_19 gnd C_wl
Rw69_19 word69_19 word68_19 R_wl
Cwl_69_19 word69_19 gnd C_wl
Rw70_19 word70_19 word69_19 R_wl
Cwl_70_19 word70_19 gnd C_wl
Rw71_19 word71_19 word70_19 R_wl
Cwl_71_19 word71_19 gnd C_wl
Rw72_19 word72_19 word71_19 R_wl
Cwl_72_19 word72_19 gnd C_wl
Rw73_19 word73_19 word72_19 R_wl
Cwl_73_19 word73_19 gnd C_wl
Rw74_19 word74_19 word73_19 R_wl
Cwl_74_19 word74_19 gnd C_wl
Rw75_19 word75_19 word74_19 R_wl
Cwl_75_19 word75_19 gnd C_wl
Rw76_19 word76_19 word75_19 R_wl
Cwl_76_19 word76_19 gnd C_wl
Rw77_19 word77_19 word76_19 R_wl
Cwl_77_19 word77_19 gnd C_wl
Rw78_19 word78_19 word77_19 R_wl
Cwl_78_19 word78_19 gnd C_wl
Rw79_19 word79_19 word78_19 R_wl
Cwl_79_19 word79_19 gnd C_wl
Rw80_19 word80_19 word79_19 R_wl
Cwl_80_19 word80_19 gnd C_wl
Rw81_19 word81_19 word80_19 R_wl
Cwl_81_19 word81_19 gnd C_wl
Rw82_19 word82_19 word81_19 R_wl
Cwl_82_19 word82_19 gnd C_wl
Rw83_19 word83_19 word82_19 R_wl
Cwl_83_19 word83_19 gnd C_wl
Rw84_19 word84_19 word83_19 R_wl
Cwl_84_19 word84_19 gnd C_wl
Rw85_19 word85_19 word84_19 R_wl
Cwl_85_19 word85_19 gnd C_wl
Rw86_19 word86_19 word85_19 R_wl
Cwl_86_19 word86_19 gnd C_wl
Rw87_19 word87_19 word86_19 R_wl
Cwl_87_19 word87_19 gnd C_wl
Rw88_19 word88_19 word87_19 R_wl
Cwl_88_19 word88_19 gnd C_wl
Rw89_19 word89_19 word88_19 R_wl
Cwl_89_19 word89_19 gnd C_wl
Rw90_19 word90_19 word89_19 R_wl
Cwl_90_19 word90_19 gnd C_wl
Rw91_19 word91_19 word90_19 R_wl
Cwl_91_19 word91_19 gnd C_wl
Rw92_19 word92_19 word91_19 R_wl
Cwl_92_19 word92_19 gnd C_wl
Rw93_19 word93_19 word92_19 R_wl
Cwl_93_19 word93_19 gnd C_wl
Rw94_19 word94_19 word93_19 R_wl
Cwl_94_19 word94_19 gnd C_wl
Rw95_19 word95_19 word94_19 R_wl
Cwl_95_19 word95_19 gnd C_wl
Rw96_19 word96_19 word95_19 R_wl
Cwl_96_19 word96_19 gnd C_wl
Rw97_19 word97_19 word96_19 R_wl
Cwl_97_19 word97_19 gnd C_wl
Rw98_19 word98_19 word97_19 R_wl
Cwl_98_19 word98_19 gnd C_wl
Rw99_19 word99_19 word98_19 R_wl
Cwl_99_19 word99_19 gnd C_wl
Vwl_20 word_20 0 0
Rw0_20 word_20 word0_20 R_wl
Cwl_0_20 word0_20 gnd C_wl
Rw1_20 word1_20 word0_20 R_wl
Cwl_1_20 word1_20 gnd C_wl
Rw2_20 word2_20 word1_20 R_wl
Cwl_2_20 word2_20 gnd C_wl
Rw3_20 word3_20 word2_20 R_wl
Cwl_3_20 word3_20 gnd C_wl
Rw4_20 word4_20 word3_20 R_wl
Cwl_4_20 word4_20 gnd C_wl
Rw5_20 word5_20 word4_20 R_wl
Cwl_5_20 word5_20 gnd C_wl
Rw6_20 word6_20 word5_20 R_wl
Cwl_6_20 word6_20 gnd C_wl
Rw7_20 word7_20 word6_20 R_wl
Cwl_7_20 word7_20 gnd C_wl
Rw8_20 word8_20 word7_20 R_wl
Cwl_8_20 word8_20 gnd C_wl
Rw9_20 word9_20 word8_20 R_wl
Cwl_9_20 word9_20 gnd C_wl
Rw10_20 word10_20 word9_20 R_wl
Cwl_10_20 word10_20 gnd C_wl
Rw11_20 word11_20 word10_20 R_wl
Cwl_11_20 word11_20 gnd C_wl
Rw12_20 word12_20 word11_20 R_wl
Cwl_12_20 word12_20 gnd C_wl
Rw13_20 word13_20 word12_20 R_wl
Cwl_13_20 word13_20 gnd C_wl
Rw14_20 word14_20 word13_20 R_wl
Cwl_14_20 word14_20 gnd C_wl
Rw15_20 word15_20 word14_20 R_wl
Cwl_15_20 word15_20 gnd C_wl
Rw16_20 word16_20 word15_20 R_wl
Cwl_16_20 word16_20 gnd C_wl
Rw17_20 word17_20 word16_20 R_wl
Cwl_17_20 word17_20 gnd C_wl
Rw18_20 word18_20 word17_20 R_wl
Cwl_18_20 word18_20 gnd C_wl
Rw19_20 word19_20 word18_20 R_wl
Cwl_19_20 word19_20 gnd C_wl
Rw20_20 word20_20 word19_20 R_wl
Cwl_20_20 word20_20 gnd C_wl
Rw21_20 word21_20 word20_20 R_wl
Cwl_21_20 word21_20 gnd C_wl
Rw22_20 word22_20 word21_20 R_wl
Cwl_22_20 word22_20 gnd C_wl
Rw23_20 word23_20 word22_20 R_wl
Cwl_23_20 word23_20 gnd C_wl
Rw24_20 word24_20 word23_20 R_wl
Cwl_24_20 word24_20 gnd C_wl
Rw25_20 word25_20 word24_20 R_wl
Cwl_25_20 word25_20 gnd C_wl
Rw26_20 word26_20 word25_20 R_wl
Cwl_26_20 word26_20 gnd C_wl
Rw27_20 word27_20 word26_20 R_wl
Cwl_27_20 word27_20 gnd C_wl
Rw28_20 word28_20 word27_20 R_wl
Cwl_28_20 word28_20 gnd C_wl
Rw29_20 word29_20 word28_20 R_wl
Cwl_29_20 word29_20 gnd C_wl
Rw30_20 word30_20 word29_20 R_wl
Cwl_30_20 word30_20 gnd C_wl
Rw31_20 word31_20 word30_20 R_wl
Cwl_31_20 word31_20 gnd C_wl
Rw32_20 word32_20 word31_20 R_wl
Cwl_32_20 word32_20 gnd C_wl
Rw33_20 word33_20 word32_20 R_wl
Cwl_33_20 word33_20 gnd C_wl
Rw34_20 word34_20 word33_20 R_wl
Cwl_34_20 word34_20 gnd C_wl
Rw35_20 word35_20 word34_20 R_wl
Cwl_35_20 word35_20 gnd C_wl
Rw36_20 word36_20 word35_20 R_wl
Cwl_36_20 word36_20 gnd C_wl
Rw37_20 word37_20 word36_20 R_wl
Cwl_37_20 word37_20 gnd C_wl
Rw38_20 word38_20 word37_20 R_wl
Cwl_38_20 word38_20 gnd C_wl
Rw39_20 word39_20 word38_20 R_wl
Cwl_39_20 word39_20 gnd C_wl
Rw40_20 word40_20 word39_20 R_wl
Cwl_40_20 word40_20 gnd C_wl
Rw41_20 word41_20 word40_20 R_wl
Cwl_41_20 word41_20 gnd C_wl
Rw42_20 word42_20 word41_20 R_wl
Cwl_42_20 word42_20 gnd C_wl
Rw43_20 word43_20 word42_20 R_wl
Cwl_43_20 word43_20 gnd C_wl
Rw44_20 word44_20 word43_20 R_wl
Cwl_44_20 word44_20 gnd C_wl
Rw45_20 word45_20 word44_20 R_wl
Cwl_45_20 word45_20 gnd C_wl
Rw46_20 word46_20 word45_20 R_wl
Cwl_46_20 word46_20 gnd C_wl
Rw47_20 word47_20 word46_20 R_wl
Cwl_47_20 word47_20 gnd C_wl
Rw48_20 word48_20 word47_20 R_wl
Cwl_48_20 word48_20 gnd C_wl
Rw49_20 word49_20 word48_20 R_wl
Cwl_49_20 word49_20 gnd C_wl
Rw50_20 word50_20 word49_20 R_wl
Cwl_50_20 word50_20 gnd C_wl
Rw51_20 word51_20 word50_20 R_wl
Cwl_51_20 word51_20 gnd C_wl
Rw52_20 word52_20 word51_20 R_wl
Cwl_52_20 word52_20 gnd C_wl
Rw53_20 word53_20 word52_20 R_wl
Cwl_53_20 word53_20 gnd C_wl
Rw54_20 word54_20 word53_20 R_wl
Cwl_54_20 word54_20 gnd C_wl
Rw55_20 word55_20 word54_20 R_wl
Cwl_55_20 word55_20 gnd C_wl
Rw56_20 word56_20 word55_20 R_wl
Cwl_56_20 word56_20 gnd C_wl
Rw57_20 word57_20 word56_20 R_wl
Cwl_57_20 word57_20 gnd C_wl
Rw58_20 word58_20 word57_20 R_wl
Cwl_58_20 word58_20 gnd C_wl
Rw59_20 word59_20 word58_20 R_wl
Cwl_59_20 word59_20 gnd C_wl
Rw60_20 word60_20 word59_20 R_wl
Cwl_60_20 word60_20 gnd C_wl
Rw61_20 word61_20 word60_20 R_wl
Cwl_61_20 word61_20 gnd C_wl
Rw62_20 word62_20 word61_20 R_wl
Cwl_62_20 word62_20 gnd C_wl
Rw63_20 word63_20 word62_20 R_wl
Cwl_63_20 word63_20 gnd C_wl
Rw64_20 word64_20 word63_20 R_wl
Cwl_64_20 word64_20 gnd C_wl
Rw65_20 word65_20 word64_20 R_wl
Cwl_65_20 word65_20 gnd C_wl
Rw66_20 word66_20 word65_20 R_wl
Cwl_66_20 word66_20 gnd C_wl
Rw67_20 word67_20 word66_20 R_wl
Cwl_67_20 word67_20 gnd C_wl
Rw68_20 word68_20 word67_20 R_wl
Cwl_68_20 word68_20 gnd C_wl
Rw69_20 word69_20 word68_20 R_wl
Cwl_69_20 word69_20 gnd C_wl
Rw70_20 word70_20 word69_20 R_wl
Cwl_70_20 word70_20 gnd C_wl
Rw71_20 word71_20 word70_20 R_wl
Cwl_71_20 word71_20 gnd C_wl
Rw72_20 word72_20 word71_20 R_wl
Cwl_72_20 word72_20 gnd C_wl
Rw73_20 word73_20 word72_20 R_wl
Cwl_73_20 word73_20 gnd C_wl
Rw74_20 word74_20 word73_20 R_wl
Cwl_74_20 word74_20 gnd C_wl
Rw75_20 word75_20 word74_20 R_wl
Cwl_75_20 word75_20 gnd C_wl
Rw76_20 word76_20 word75_20 R_wl
Cwl_76_20 word76_20 gnd C_wl
Rw77_20 word77_20 word76_20 R_wl
Cwl_77_20 word77_20 gnd C_wl
Rw78_20 word78_20 word77_20 R_wl
Cwl_78_20 word78_20 gnd C_wl
Rw79_20 word79_20 word78_20 R_wl
Cwl_79_20 word79_20 gnd C_wl
Rw80_20 word80_20 word79_20 R_wl
Cwl_80_20 word80_20 gnd C_wl
Rw81_20 word81_20 word80_20 R_wl
Cwl_81_20 word81_20 gnd C_wl
Rw82_20 word82_20 word81_20 R_wl
Cwl_82_20 word82_20 gnd C_wl
Rw83_20 word83_20 word82_20 R_wl
Cwl_83_20 word83_20 gnd C_wl
Rw84_20 word84_20 word83_20 R_wl
Cwl_84_20 word84_20 gnd C_wl
Rw85_20 word85_20 word84_20 R_wl
Cwl_85_20 word85_20 gnd C_wl
Rw86_20 word86_20 word85_20 R_wl
Cwl_86_20 word86_20 gnd C_wl
Rw87_20 word87_20 word86_20 R_wl
Cwl_87_20 word87_20 gnd C_wl
Rw88_20 word88_20 word87_20 R_wl
Cwl_88_20 word88_20 gnd C_wl
Rw89_20 word89_20 word88_20 R_wl
Cwl_89_20 word89_20 gnd C_wl
Rw90_20 word90_20 word89_20 R_wl
Cwl_90_20 word90_20 gnd C_wl
Rw91_20 word91_20 word90_20 R_wl
Cwl_91_20 word91_20 gnd C_wl
Rw92_20 word92_20 word91_20 R_wl
Cwl_92_20 word92_20 gnd C_wl
Rw93_20 word93_20 word92_20 R_wl
Cwl_93_20 word93_20 gnd C_wl
Rw94_20 word94_20 word93_20 R_wl
Cwl_94_20 word94_20 gnd C_wl
Rw95_20 word95_20 word94_20 R_wl
Cwl_95_20 word95_20 gnd C_wl
Rw96_20 word96_20 word95_20 R_wl
Cwl_96_20 word96_20 gnd C_wl
Rw97_20 word97_20 word96_20 R_wl
Cwl_97_20 word97_20 gnd C_wl
Rw98_20 word98_20 word97_20 R_wl
Cwl_98_20 word98_20 gnd C_wl
Rw99_20 word99_20 word98_20 R_wl
Cwl_99_20 word99_20 gnd C_wl
Vwl_21 word_21 0 0
Rw0_21 word_21 word0_21 R_wl
Cwl_0_21 word0_21 gnd C_wl
Rw1_21 word1_21 word0_21 R_wl
Cwl_1_21 word1_21 gnd C_wl
Rw2_21 word2_21 word1_21 R_wl
Cwl_2_21 word2_21 gnd C_wl
Rw3_21 word3_21 word2_21 R_wl
Cwl_3_21 word3_21 gnd C_wl
Rw4_21 word4_21 word3_21 R_wl
Cwl_4_21 word4_21 gnd C_wl
Rw5_21 word5_21 word4_21 R_wl
Cwl_5_21 word5_21 gnd C_wl
Rw6_21 word6_21 word5_21 R_wl
Cwl_6_21 word6_21 gnd C_wl
Rw7_21 word7_21 word6_21 R_wl
Cwl_7_21 word7_21 gnd C_wl
Rw8_21 word8_21 word7_21 R_wl
Cwl_8_21 word8_21 gnd C_wl
Rw9_21 word9_21 word8_21 R_wl
Cwl_9_21 word9_21 gnd C_wl
Rw10_21 word10_21 word9_21 R_wl
Cwl_10_21 word10_21 gnd C_wl
Rw11_21 word11_21 word10_21 R_wl
Cwl_11_21 word11_21 gnd C_wl
Rw12_21 word12_21 word11_21 R_wl
Cwl_12_21 word12_21 gnd C_wl
Rw13_21 word13_21 word12_21 R_wl
Cwl_13_21 word13_21 gnd C_wl
Rw14_21 word14_21 word13_21 R_wl
Cwl_14_21 word14_21 gnd C_wl
Rw15_21 word15_21 word14_21 R_wl
Cwl_15_21 word15_21 gnd C_wl
Rw16_21 word16_21 word15_21 R_wl
Cwl_16_21 word16_21 gnd C_wl
Rw17_21 word17_21 word16_21 R_wl
Cwl_17_21 word17_21 gnd C_wl
Rw18_21 word18_21 word17_21 R_wl
Cwl_18_21 word18_21 gnd C_wl
Rw19_21 word19_21 word18_21 R_wl
Cwl_19_21 word19_21 gnd C_wl
Rw20_21 word20_21 word19_21 R_wl
Cwl_20_21 word20_21 gnd C_wl
Rw21_21 word21_21 word20_21 R_wl
Cwl_21_21 word21_21 gnd C_wl
Rw22_21 word22_21 word21_21 R_wl
Cwl_22_21 word22_21 gnd C_wl
Rw23_21 word23_21 word22_21 R_wl
Cwl_23_21 word23_21 gnd C_wl
Rw24_21 word24_21 word23_21 R_wl
Cwl_24_21 word24_21 gnd C_wl
Rw25_21 word25_21 word24_21 R_wl
Cwl_25_21 word25_21 gnd C_wl
Rw26_21 word26_21 word25_21 R_wl
Cwl_26_21 word26_21 gnd C_wl
Rw27_21 word27_21 word26_21 R_wl
Cwl_27_21 word27_21 gnd C_wl
Rw28_21 word28_21 word27_21 R_wl
Cwl_28_21 word28_21 gnd C_wl
Rw29_21 word29_21 word28_21 R_wl
Cwl_29_21 word29_21 gnd C_wl
Rw30_21 word30_21 word29_21 R_wl
Cwl_30_21 word30_21 gnd C_wl
Rw31_21 word31_21 word30_21 R_wl
Cwl_31_21 word31_21 gnd C_wl
Rw32_21 word32_21 word31_21 R_wl
Cwl_32_21 word32_21 gnd C_wl
Rw33_21 word33_21 word32_21 R_wl
Cwl_33_21 word33_21 gnd C_wl
Rw34_21 word34_21 word33_21 R_wl
Cwl_34_21 word34_21 gnd C_wl
Rw35_21 word35_21 word34_21 R_wl
Cwl_35_21 word35_21 gnd C_wl
Rw36_21 word36_21 word35_21 R_wl
Cwl_36_21 word36_21 gnd C_wl
Rw37_21 word37_21 word36_21 R_wl
Cwl_37_21 word37_21 gnd C_wl
Rw38_21 word38_21 word37_21 R_wl
Cwl_38_21 word38_21 gnd C_wl
Rw39_21 word39_21 word38_21 R_wl
Cwl_39_21 word39_21 gnd C_wl
Rw40_21 word40_21 word39_21 R_wl
Cwl_40_21 word40_21 gnd C_wl
Rw41_21 word41_21 word40_21 R_wl
Cwl_41_21 word41_21 gnd C_wl
Rw42_21 word42_21 word41_21 R_wl
Cwl_42_21 word42_21 gnd C_wl
Rw43_21 word43_21 word42_21 R_wl
Cwl_43_21 word43_21 gnd C_wl
Rw44_21 word44_21 word43_21 R_wl
Cwl_44_21 word44_21 gnd C_wl
Rw45_21 word45_21 word44_21 R_wl
Cwl_45_21 word45_21 gnd C_wl
Rw46_21 word46_21 word45_21 R_wl
Cwl_46_21 word46_21 gnd C_wl
Rw47_21 word47_21 word46_21 R_wl
Cwl_47_21 word47_21 gnd C_wl
Rw48_21 word48_21 word47_21 R_wl
Cwl_48_21 word48_21 gnd C_wl
Rw49_21 word49_21 word48_21 R_wl
Cwl_49_21 word49_21 gnd C_wl
Rw50_21 word50_21 word49_21 R_wl
Cwl_50_21 word50_21 gnd C_wl
Rw51_21 word51_21 word50_21 R_wl
Cwl_51_21 word51_21 gnd C_wl
Rw52_21 word52_21 word51_21 R_wl
Cwl_52_21 word52_21 gnd C_wl
Rw53_21 word53_21 word52_21 R_wl
Cwl_53_21 word53_21 gnd C_wl
Rw54_21 word54_21 word53_21 R_wl
Cwl_54_21 word54_21 gnd C_wl
Rw55_21 word55_21 word54_21 R_wl
Cwl_55_21 word55_21 gnd C_wl
Rw56_21 word56_21 word55_21 R_wl
Cwl_56_21 word56_21 gnd C_wl
Rw57_21 word57_21 word56_21 R_wl
Cwl_57_21 word57_21 gnd C_wl
Rw58_21 word58_21 word57_21 R_wl
Cwl_58_21 word58_21 gnd C_wl
Rw59_21 word59_21 word58_21 R_wl
Cwl_59_21 word59_21 gnd C_wl
Rw60_21 word60_21 word59_21 R_wl
Cwl_60_21 word60_21 gnd C_wl
Rw61_21 word61_21 word60_21 R_wl
Cwl_61_21 word61_21 gnd C_wl
Rw62_21 word62_21 word61_21 R_wl
Cwl_62_21 word62_21 gnd C_wl
Rw63_21 word63_21 word62_21 R_wl
Cwl_63_21 word63_21 gnd C_wl
Rw64_21 word64_21 word63_21 R_wl
Cwl_64_21 word64_21 gnd C_wl
Rw65_21 word65_21 word64_21 R_wl
Cwl_65_21 word65_21 gnd C_wl
Rw66_21 word66_21 word65_21 R_wl
Cwl_66_21 word66_21 gnd C_wl
Rw67_21 word67_21 word66_21 R_wl
Cwl_67_21 word67_21 gnd C_wl
Rw68_21 word68_21 word67_21 R_wl
Cwl_68_21 word68_21 gnd C_wl
Rw69_21 word69_21 word68_21 R_wl
Cwl_69_21 word69_21 gnd C_wl
Rw70_21 word70_21 word69_21 R_wl
Cwl_70_21 word70_21 gnd C_wl
Rw71_21 word71_21 word70_21 R_wl
Cwl_71_21 word71_21 gnd C_wl
Rw72_21 word72_21 word71_21 R_wl
Cwl_72_21 word72_21 gnd C_wl
Rw73_21 word73_21 word72_21 R_wl
Cwl_73_21 word73_21 gnd C_wl
Rw74_21 word74_21 word73_21 R_wl
Cwl_74_21 word74_21 gnd C_wl
Rw75_21 word75_21 word74_21 R_wl
Cwl_75_21 word75_21 gnd C_wl
Rw76_21 word76_21 word75_21 R_wl
Cwl_76_21 word76_21 gnd C_wl
Rw77_21 word77_21 word76_21 R_wl
Cwl_77_21 word77_21 gnd C_wl
Rw78_21 word78_21 word77_21 R_wl
Cwl_78_21 word78_21 gnd C_wl
Rw79_21 word79_21 word78_21 R_wl
Cwl_79_21 word79_21 gnd C_wl
Rw80_21 word80_21 word79_21 R_wl
Cwl_80_21 word80_21 gnd C_wl
Rw81_21 word81_21 word80_21 R_wl
Cwl_81_21 word81_21 gnd C_wl
Rw82_21 word82_21 word81_21 R_wl
Cwl_82_21 word82_21 gnd C_wl
Rw83_21 word83_21 word82_21 R_wl
Cwl_83_21 word83_21 gnd C_wl
Rw84_21 word84_21 word83_21 R_wl
Cwl_84_21 word84_21 gnd C_wl
Rw85_21 word85_21 word84_21 R_wl
Cwl_85_21 word85_21 gnd C_wl
Rw86_21 word86_21 word85_21 R_wl
Cwl_86_21 word86_21 gnd C_wl
Rw87_21 word87_21 word86_21 R_wl
Cwl_87_21 word87_21 gnd C_wl
Rw88_21 word88_21 word87_21 R_wl
Cwl_88_21 word88_21 gnd C_wl
Rw89_21 word89_21 word88_21 R_wl
Cwl_89_21 word89_21 gnd C_wl
Rw90_21 word90_21 word89_21 R_wl
Cwl_90_21 word90_21 gnd C_wl
Rw91_21 word91_21 word90_21 R_wl
Cwl_91_21 word91_21 gnd C_wl
Rw92_21 word92_21 word91_21 R_wl
Cwl_92_21 word92_21 gnd C_wl
Rw93_21 word93_21 word92_21 R_wl
Cwl_93_21 word93_21 gnd C_wl
Rw94_21 word94_21 word93_21 R_wl
Cwl_94_21 word94_21 gnd C_wl
Rw95_21 word95_21 word94_21 R_wl
Cwl_95_21 word95_21 gnd C_wl
Rw96_21 word96_21 word95_21 R_wl
Cwl_96_21 word96_21 gnd C_wl
Rw97_21 word97_21 word96_21 R_wl
Cwl_97_21 word97_21 gnd C_wl
Rw98_21 word98_21 word97_21 R_wl
Cwl_98_21 word98_21 gnd C_wl
Rw99_21 word99_21 word98_21 R_wl
Cwl_99_21 word99_21 gnd C_wl
Vwl_22 word_22 0 0
Rw0_22 word_22 word0_22 R_wl
Cwl_0_22 word0_22 gnd C_wl
Rw1_22 word1_22 word0_22 R_wl
Cwl_1_22 word1_22 gnd C_wl
Rw2_22 word2_22 word1_22 R_wl
Cwl_2_22 word2_22 gnd C_wl
Rw3_22 word3_22 word2_22 R_wl
Cwl_3_22 word3_22 gnd C_wl
Rw4_22 word4_22 word3_22 R_wl
Cwl_4_22 word4_22 gnd C_wl
Rw5_22 word5_22 word4_22 R_wl
Cwl_5_22 word5_22 gnd C_wl
Rw6_22 word6_22 word5_22 R_wl
Cwl_6_22 word6_22 gnd C_wl
Rw7_22 word7_22 word6_22 R_wl
Cwl_7_22 word7_22 gnd C_wl
Rw8_22 word8_22 word7_22 R_wl
Cwl_8_22 word8_22 gnd C_wl
Rw9_22 word9_22 word8_22 R_wl
Cwl_9_22 word9_22 gnd C_wl
Rw10_22 word10_22 word9_22 R_wl
Cwl_10_22 word10_22 gnd C_wl
Rw11_22 word11_22 word10_22 R_wl
Cwl_11_22 word11_22 gnd C_wl
Rw12_22 word12_22 word11_22 R_wl
Cwl_12_22 word12_22 gnd C_wl
Rw13_22 word13_22 word12_22 R_wl
Cwl_13_22 word13_22 gnd C_wl
Rw14_22 word14_22 word13_22 R_wl
Cwl_14_22 word14_22 gnd C_wl
Rw15_22 word15_22 word14_22 R_wl
Cwl_15_22 word15_22 gnd C_wl
Rw16_22 word16_22 word15_22 R_wl
Cwl_16_22 word16_22 gnd C_wl
Rw17_22 word17_22 word16_22 R_wl
Cwl_17_22 word17_22 gnd C_wl
Rw18_22 word18_22 word17_22 R_wl
Cwl_18_22 word18_22 gnd C_wl
Rw19_22 word19_22 word18_22 R_wl
Cwl_19_22 word19_22 gnd C_wl
Rw20_22 word20_22 word19_22 R_wl
Cwl_20_22 word20_22 gnd C_wl
Rw21_22 word21_22 word20_22 R_wl
Cwl_21_22 word21_22 gnd C_wl
Rw22_22 word22_22 word21_22 R_wl
Cwl_22_22 word22_22 gnd C_wl
Rw23_22 word23_22 word22_22 R_wl
Cwl_23_22 word23_22 gnd C_wl
Rw24_22 word24_22 word23_22 R_wl
Cwl_24_22 word24_22 gnd C_wl
Rw25_22 word25_22 word24_22 R_wl
Cwl_25_22 word25_22 gnd C_wl
Rw26_22 word26_22 word25_22 R_wl
Cwl_26_22 word26_22 gnd C_wl
Rw27_22 word27_22 word26_22 R_wl
Cwl_27_22 word27_22 gnd C_wl
Rw28_22 word28_22 word27_22 R_wl
Cwl_28_22 word28_22 gnd C_wl
Rw29_22 word29_22 word28_22 R_wl
Cwl_29_22 word29_22 gnd C_wl
Rw30_22 word30_22 word29_22 R_wl
Cwl_30_22 word30_22 gnd C_wl
Rw31_22 word31_22 word30_22 R_wl
Cwl_31_22 word31_22 gnd C_wl
Rw32_22 word32_22 word31_22 R_wl
Cwl_32_22 word32_22 gnd C_wl
Rw33_22 word33_22 word32_22 R_wl
Cwl_33_22 word33_22 gnd C_wl
Rw34_22 word34_22 word33_22 R_wl
Cwl_34_22 word34_22 gnd C_wl
Rw35_22 word35_22 word34_22 R_wl
Cwl_35_22 word35_22 gnd C_wl
Rw36_22 word36_22 word35_22 R_wl
Cwl_36_22 word36_22 gnd C_wl
Rw37_22 word37_22 word36_22 R_wl
Cwl_37_22 word37_22 gnd C_wl
Rw38_22 word38_22 word37_22 R_wl
Cwl_38_22 word38_22 gnd C_wl
Rw39_22 word39_22 word38_22 R_wl
Cwl_39_22 word39_22 gnd C_wl
Rw40_22 word40_22 word39_22 R_wl
Cwl_40_22 word40_22 gnd C_wl
Rw41_22 word41_22 word40_22 R_wl
Cwl_41_22 word41_22 gnd C_wl
Rw42_22 word42_22 word41_22 R_wl
Cwl_42_22 word42_22 gnd C_wl
Rw43_22 word43_22 word42_22 R_wl
Cwl_43_22 word43_22 gnd C_wl
Rw44_22 word44_22 word43_22 R_wl
Cwl_44_22 word44_22 gnd C_wl
Rw45_22 word45_22 word44_22 R_wl
Cwl_45_22 word45_22 gnd C_wl
Rw46_22 word46_22 word45_22 R_wl
Cwl_46_22 word46_22 gnd C_wl
Rw47_22 word47_22 word46_22 R_wl
Cwl_47_22 word47_22 gnd C_wl
Rw48_22 word48_22 word47_22 R_wl
Cwl_48_22 word48_22 gnd C_wl
Rw49_22 word49_22 word48_22 R_wl
Cwl_49_22 word49_22 gnd C_wl
Rw50_22 word50_22 word49_22 R_wl
Cwl_50_22 word50_22 gnd C_wl
Rw51_22 word51_22 word50_22 R_wl
Cwl_51_22 word51_22 gnd C_wl
Rw52_22 word52_22 word51_22 R_wl
Cwl_52_22 word52_22 gnd C_wl
Rw53_22 word53_22 word52_22 R_wl
Cwl_53_22 word53_22 gnd C_wl
Rw54_22 word54_22 word53_22 R_wl
Cwl_54_22 word54_22 gnd C_wl
Rw55_22 word55_22 word54_22 R_wl
Cwl_55_22 word55_22 gnd C_wl
Rw56_22 word56_22 word55_22 R_wl
Cwl_56_22 word56_22 gnd C_wl
Rw57_22 word57_22 word56_22 R_wl
Cwl_57_22 word57_22 gnd C_wl
Rw58_22 word58_22 word57_22 R_wl
Cwl_58_22 word58_22 gnd C_wl
Rw59_22 word59_22 word58_22 R_wl
Cwl_59_22 word59_22 gnd C_wl
Rw60_22 word60_22 word59_22 R_wl
Cwl_60_22 word60_22 gnd C_wl
Rw61_22 word61_22 word60_22 R_wl
Cwl_61_22 word61_22 gnd C_wl
Rw62_22 word62_22 word61_22 R_wl
Cwl_62_22 word62_22 gnd C_wl
Rw63_22 word63_22 word62_22 R_wl
Cwl_63_22 word63_22 gnd C_wl
Rw64_22 word64_22 word63_22 R_wl
Cwl_64_22 word64_22 gnd C_wl
Rw65_22 word65_22 word64_22 R_wl
Cwl_65_22 word65_22 gnd C_wl
Rw66_22 word66_22 word65_22 R_wl
Cwl_66_22 word66_22 gnd C_wl
Rw67_22 word67_22 word66_22 R_wl
Cwl_67_22 word67_22 gnd C_wl
Rw68_22 word68_22 word67_22 R_wl
Cwl_68_22 word68_22 gnd C_wl
Rw69_22 word69_22 word68_22 R_wl
Cwl_69_22 word69_22 gnd C_wl
Rw70_22 word70_22 word69_22 R_wl
Cwl_70_22 word70_22 gnd C_wl
Rw71_22 word71_22 word70_22 R_wl
Cwl_71_22 word71_22 gnd C_wl
Rw72_22 word72_22 word71_22 R_wl
Cwl_72_22 word72_22 gnd C_wl
Rw73_22 word73_22 word72_22 R_wl
Cwl_73_22 word73_22 gnd C_wl
Rw74_22 word74_22 word73_22 R_wl
Cwl_74_22 word74_22 gnd C_wl
Rw75_22 word75_22 word74_22 R_wl
Cwl_75_22 word75_22 gnd C_wl
Rw76_22 word76_22 word75_22 R_wl
Cwl_76_22 word76_22 gnd C_wl
Rw77_22 word77_22 word76_22 R_wl
Cwl_77_22 word77_22 gnd C_wl
Rw78_22 word78_22 word77_22 R_wl
Cwl_78_22 word78_22 gnd C_wl
Rw79_22 word79_22 word78_22 R_wl
Cwl_79_22 word79_22 gnd C_wl
Rw80_22 word80_22 word79_22 R_wl
Cwl_80_22 word80_22 gnd C_wl
Rw81_22 word81_22 word80_22 R_wl
Cwl_81_22 word81_22 gnd C_wl
Rw82_22 word82_22 word81_22 R_wl
Cwl_82_22 word82_22 gnd C_wl
Rw83_22 word83_22 word82_22 R_wl
Cwl_83_22 word83_22 gnd C_wl
Rw84_22 word84_22 word83_22 R_wl
Cwl_84_22 word84_22 gnd C_wl
Rw85_22 word85_22 word84_22 R_wl
Cwl_85_22 word85_22 gnd C_wl
Rw86_22 word86_22 word85_22 R_wl
Cwl_86_22 word86_22 gnd C_wl
Rw87_22 word87_22 word86_22 R_wl
Cwl_87_22 word87_22 gnd C_wl
Rw88_22 word88_22 word87_22 R_wl
Cwl_88_22 word88_22 gnd C_wl
Rw89_22 word89_22 word88_22 R_wl
Cwl_89_22 word89_22 gnd C_wl
Rw90_22 word90_22 word89_22 R_wl
Cwl_90_22 word90_22 gnd C_wl
Rw91_22 word91_22 word90_22 R_wl
Cwl_91_22 word91_22 gnd C_wl
Rw92_22 word92_22 word91_22 R_wl
Cwl_92_22 word92_22 gnd C_wl
Rw93_22 word93_22 word92_22 R_wl
Cwl_93_22 word93_22 gnd C_wl
Rw94_22 word94_22 word93_22 R_wl
Cwl_94_22 word94_22 gnd C_wl
Rw95_22 word95_22 word94_22 R_wl
Cwl_95_22 word95_22 gnd C_wl
Rw96_22 word96_22 word95_22 R_wl
Cwl_96_22 word96_22 gnd C_wl
Rw97_22 word97_22 word96_22 R_wl
Cwl_97_22 word97_22 gnd C_wl
Rw98_22 word98_22 word97_22 R_wl
Cwl_98_22 word98_22 gnd C_wl
Rw99_22 word99_22 word98_22 R_wl
Cwl_99_22 word99_22 gnd C_wl
Vwl_23 word_23 0 0
Rw0_23 word_23 word0_23 R_wl
Cwl_0_23 word0_23 gnd C_wl
Rw1_23 word1_23 word0_23 R_wl
Cwl_1_23 word1_23 gnd C_wl
Rw2_23 word2_23 word1_23 R_wl
Cwl_2_23 word2_23 gnd C_wl
Rw3_23 word3_23 word2_23 R_wl
Cwl_3_23 word3_23 gnd C_wl
Rw4_23 word4_23 word3_23 R_wl
Cwl_4_23 word4_23 gnd C_wl
Rw5_23 word5_23 word4_23 R_wl
Cwl_5_23 word5_23 gnd C_wl
Rw6_23 word6_23 word5_23 R_wl
Cwl_6_23 word6_23 gnd C_wl
Rw7_23 word7_23 word6_23 R_wl
Cwl_7_23 word7_23 gnd C_wl
Rw8_23 word8_23 word7_23 R_wl
Cwl_8_23 word8_23 gnd C_wl
Rw9_23 word9_23 word8_23 R_wl
Cwl_9_23 word9_23 gnd C_wl
Rw10_23 word10_23 word9_23 R_wl
Cwl_10_23 word10_23 gnd C_wl
Rw11_23 word11_23 word10_23 R_wl
Cwl_11_23 word11_23 gnd C_wl
Rw12_23 word12_23 word11_23 R_wl
Cwl_12_23 word12_23 gnd C_wl
Rw13_23 word13_23 word12_23 R_wl
Cwl_13_23 word13_23 gnd C_wl
Rw14_23 word14_23 word13_23 R_wl
Cwl_14_23 word14_23 gnd C_wl
Rw15_23 word15_23 word14_23 R_wl
Cwl_15_23 word15_23 gnd C_wl
Rw16_23 word16_23 word15_23 R_wl
Cwl_16_23 word16_23 gnd C_wl
Rw17_23 word17_23 word16_23 R_wl
Cwl_17_23 word17_23 gnd C_wl
Rw18_23 word18_23 word17_23 R_wl
Cwl_18_23 word18_23 gnd C_wl
Rw19_23 word19_23 word18_23 R_wl
Cwl_19_23 word19_23 gnd C_wl
Rw20_23 word20_23 word19_23 R_wl
Cwl_20_23 word20_23 gnd C_wl
Rw21_23 word21_23 word20_23 R_wl
Cwl_21_23 word21_23 gnd C_wl
Rw22_23 word22_23 word21_23 R_wl
Cwl_22_23 word22_23 gnd C_wl
Rw23_23 word23_23 word22_23 R_wl
Cwl_23_23 word23_23 gnd C_wl
Rw24_23 word24_23 word23_23 R_wl
Cwl_24_23 word24_23 gnd C_wl
Rw25_23 word25_23 word24_23 R_wl
Cwl_25_23 word25_23 gnd C_wl
Rw26_23 word26_23 word25_23 R_wl
Cwl_26_23 word26_23 gnd C_wl
Rw27_23 word27_23 word26_23 R_wl
Cwl_27_23 word27_23 gnd C_wl
Rw28_23 word28_23 word27_23 R_wl
Cwl_28_23 word28_23 gnd C_wl
Rw29_23 word29_23 word28_23 R_wl
Cwl_29_23 word29_23 gnd C_wl
Rw30_23 word30_23 word29_23 R_wl
Cwl_30_23 word30_23 gnd C_wl
Rw31_23 word31_23 word30_23 R_wl
Cwl_31_23 word31_23 gnd C_wl
Rw32_23 word32_23 word31_23 R_wl
Cwl_32_23 word32_23 gnd C_wl
Rw33_23 word33_23 word32_23 R_wl
Cwl_33_23 word33_23 gnd C_wl
Rw34_23 word34_23 word33_23 R_wl
Cwl_34_23 word34_23 gnd C_wl
Rw35_23 word35_23 word34_23 R_wl
Cwl_35_23 word35_23 gnd C_wl
Rw36_23 word36_23 word35_23 R_wl
Cwl_36_23 word36_23 gnd C_wl
Rw37_23 word37_23 word36_23 R_wl
Cwl_37_23 word37_23 gnd C_wl
Rw38_23 word38_23 word37_23 R_wl
Cwl_38_23 word38_23 gnd C_wl
Rw39_23 word39_23 word38_23 R_wl
Cwl_39_23 word39_23 gnd C_wl
Rw40_23 word40_23 word39_23 R_wl
Cwl_40_23 word40_23 gnd C_wl
Rw41_23 word41_23 word40_23 R_wl
Cwl_41_23 word41_23 gnd C_wl
Rw42_23 word42_23 word41_23 R_wl
Cwl_42_23 word42_23 gnd C_wl
Rw43_23 word43_23 word42_23 R_wl
Cwl_43_23 word43_23 gnd C_wl
Rw44_23 word44_23 word43_23 R_wl
Cwl_44_23 word44_23 gnd C_wl
Rw45_23 word45_23 word44_23 R_wl
Cwl_45_23 word45_23 gnd C_wl
Rw46_23 word46_23 word45_23 R_wl
Cwl_46_23 word46_23 gnd C_wl
Rw47_23 word47_23 word46_23 R_wl
Cwl_47_23 word47_23 gnd C_wl
Rw48_23 word48_23 word47_23 R_wl
Cwl_48_23 word48_23 gnd C_wl
Rw49_23 word49_23 word48_23 R_wl
Cwl_49_23 word49_23 gnd C_wl
Rw50_23 word50_23 word49_23 R_wl
Cwl_50_23 word50_23 gnd C_wl
Rw51_23 word51_23 word50_23 R_wl
Cwl_51_23 word51_23 gnd C_wl
Rw52_23 word52_23 word51_23 R_wl
Cwl_52_23 word52_23 gnd C_wl
Rw53_23 word53_23 word52_23 R_wl
Cwl_53_23 word53_23 gnd C_wl
Rw54_23 word54_23 word53_23 R_wl
Cwl_54_23 word54_23 gnd C_wl
Rw55_23 word55_23 word54_23 R_wl
Cwl_55_23 word55_23 gnd C_wl
Rw56_23 word56_23 word55_23 R_wl
Cwl_56_23 word56_23 gnd C_wl
Rw57_23 word57_23 word56_23 R_wl
Cwl_57_23 word57_23 gnd C_wl
Rw58_23 word58_23 word57_23 R_wl
Cwl_58_23 word58_23 gnd C_wl
Rw59_23 word59_23 word58_23 R_wl
Cwl_59_23 word59_23 gnd C_wl
Rw60_23 word60_23 word59_23 R_wl
Cwl_60_23 word60_23 gnd C_wl
Rw61_23 word61_23 word60_23 R_wl
Cwl_61_23 word61_23 gnd C_wl
Rw62_23 word62_23 word61_23 R_wl
Cwl_62_23 word62_23 gnd C_wl
Rw63_23 word63_23 word62_23 R_wl
Cwl_63_23 word63_23 gnd C_wl
Rw64_23 word64_23 word63_23 R_wl
Cwl_64_23 word64_23 gnd C_wl
Rw65_23 word65_23 word64_23 R_wl
Cwl_65_23 word65_23 gnd C_wl
Rw66_23 word66_23 word65_23 R_wl
Cwl_66_23 word66_23 gnd C_wl
Rw67_23 word67_23 word66_23 R_wl
Cwl_67_23 word67_23 gnd C_wl
Rw68_23 word68_23 word67_23 R_wl
Cwl_68_23 word68_23 gnd C_wl
Rw69_23 word69_23 word68_23 R_wl
Cwl_69_23 word69_23 gnd C_wl
Rw70_23 word70_23 word69_23 R_wl
Cwl_70_23 word70_23 gnd C_wl
Rw71_23 word71_23 word70_23 R_wl
Cwl_71_23 word71_23 gnd C_wl
Rw72_23 word72_23 word71_23 R_wl
Cwl_72_23 word72_23 gnd C_wl
Rw73_23 word73_23 word72_23 R_wl
Cwl_73_23 word73_23 gnd C_wl
Rw74_23 word74_23 word73_23 R_wl
Cwl_74_23 word74_23 gnd C_wl
Rw75_23 word75_23 word74_23 R_wl
Cwl_75_23 word75_23 gnd C_wl
Rw76_23 word76_23 word75_23 R_wl
Cwl_76_23 word76_23 gnd C_wl
Rw77_23 word77_23 word76_23 R_wl
Cwl_77_23 word77_23 gnd C_wl
Rw78_23 word78_23 word77_23 R_wl
Cwl_78_23 word78_23 gnd C_wl
Rw79_23 word79_23 word78_23 R_wl
Cwl_79_23 word79_23 gnd C_wl
Rw80_23 word80_23 word79_23 R_wl
Cwl_80_23 word80_23 gnd C_wl
Rw81_23 word81_23 word80_23 R_wl
Cwl_81_23 word81_23 gnd C_wl
Rw82_23 word82_23 word81_23 R_wl
Cwl_82_23 word82_23 gnd C_wl
Rw83_23 word83_23 word82_23 R_wl
Cwl_83_23 word83_23 gnd C_wl
Rw84_23 word84_23 word83_23 R_wl
Cwl_84_23 word84_23 gnd C_wl
Rw85_23 word85_23 word84_23 R_wl
Cwl_85_23 word85_23 gnd C_wl
Rw86_23 word86_23 word85_23 R_wl
Cwl_86_23 word86_23 gnd C_wl
Rw87_23 word87_23 word86_23 R_wl
Cwl_87_23 word87_23 gnd C_wl
Rw88_23 word88_23 word87_23 R_wl
Cwl_88_23 word88_23 gnd C_wl
Rw89_23 word89_23 word88_23 R_wl
Cwl_89_23 word89_23 gnd C_wl
Rw90_23 word90_23 word89_23 R_wl
Cwl_90_23 word90_23 gnd C_wl
Rw91_23 word91_23 word90_23 R_wl
Cwl_91_23 word91_23 gnd C_wl
Rw92_23 word92_23 word91_23 R_wl
Cwl_92_23 word92_23 gnd C_wl
Rw93_23 word93_23 word92_23 R_wl
Cwl_93_23 word93_23 gnd C_wl
Rw94_23 word94_23 word93_23 R_wl
Cwl_94_23 word94_23 gnd C_wl
Rw95_23 word95_23 word94_23 R_wl
Cwl_95_23 word95_23 gnd C_wl
Rw96_23 word96_23 word95_23 R_wl
Cwl_96_23 word96_23 gnd C_wl
Rw97_23 word97_23 word96_23 R_wl
Cwl_97_23 word97_23 gnd C_wl
Rw98_23 word98_23 word97_23 R_wl
Cwl_98_23 word98_23 gnd C_wl
Rw99_23 word99_23 word98_23 R_wl
Cwl_99_23 word99_23 gnd C_wl
Vwl_24 word_24 0 0
Rw0_24 word_24 word0_24 R_wl
Cwl_0_24 word0_24 gnd C_wl
Rw1_24 word1_24 word0_24 R_wl
Cwl_1_24 word1_24 gnd C_wl
Rw2_24 word2_24 word1_24 R_wl
Cwl_2_24 word2_24 gnd C_wl
Rw3_24 word3_24 word2_24 R_wl
Cwl_3_24 word3_24 gnd C_wl
Rw4_24 word4_24 word3_24 R_wl
Cwl_4_24 word4_24 gnd C_wl
Rw5_24 word5_24 word4_24 R_wl
Cwl_5_24 word5_24 gnd C_wl
Rw6_24 word6_24 word5_24 R_wl
Cwl_6_24 word6_24 gnd C_wl
Rw7_24 word7_24 word6_24 R_wl
Cwl_7_24 word7_24 gnd C_wl
Rw8_24 word8_24 word7_24 R_wl
Cwl_8_24 word8_24 gnd C_wl
Rw9_24 word9_24 word8_24 R_wl
Cwl_9_24 word9_24 gnd C_wl
Rw10_24 word10_24 word9_24 R_wl
Cwl_10_24 word10_24 gnd C_wl
Rw11_24 word11_24 word10_24 R_wl
Cwl_11_24 word11_24 gnd C_wl
Rw12_24 word12_24 word11_24 R_wl
Cwl_12_24 word12_24 gnd C_wl
Rw13_24 word13_24 word12_24 R_wl
Cwl_13_24 word13_24 gnd C_wl
Rw14_24 word14_24 word13_24 R_wl
Cwl_14_24 word14_24 gnd C_wl
Rw15_24 word15_24 word14_24 R_wl
Cwl_15_24 word15_24 gnd C_wl
Rw16_24 word16_24 word15_24 R_wl
Cwl_16_24 word16_24 gnd C_wl
Rw17_24 word17_24 word16_24 R_wl
Cwl_17_24 word17_24 gnd C_wl
Rw18_24 word18_24 word17_24 R_wl
Cwl_18_24 word18_24 gnd C_wl
Rw19_24 word19_24 word18_24 R_wl
Cwl_19_24 word19_24 gnd C_wl
Rw20_24 word20_24 word19_24 R_wl
Cwl_20_24 word20_24 gnd C_wl
Rw21_24 word21_24 word20_24 R_wl
Cwl_21_24 word21_24 gnd C_wl
Rw22_24 word22_24 word21_24 R_wl
Cwl_22_24 word22_24 gnd C_wl
Rw23_24 word23_24 word22_24 R_wl
Cwl_23_24 word23_24 gnd C_wl
Rw24_24 word24_24 word23_24 R_wl
Cwl_24_24 word24_24 gnd C_wl
Rw25_24 word25_24 word24_24 R_wl
Cwl_25_24 word25_24 gnd C_wl
Rw26_24 word26_24 word25_24 R_wl
Cwl_26_24 word26_24 gnd C_wl
Rw27_24 word27_24 word26_24 R_wl
Cwl_27_24 word27_24 gnd C_wl
Rw28_24 word28_24 word27_24 R_wl
Cwl_28_24 word28_24 gnd C_wl
Rw29_24 word29_24 word28_24 R_wl
Cwl_29_24 word29_24 gnd C_wl
Rw30_24 word30_24 word29_24 R_wl
Cwl_30_24 word30_24 gnd C_wl
Rw31_24 word31_24 word30_24 R_wl
Cwl_31_24 word31_24 gnd C_wl
Rw32_24 word32_24 word31_24 R_wl
Cwl_32_24 word32_24 gnd C_wl
Rw33_24 word33_24 word32_24 R_wl
Cwl_33_24 word33_24 gnd C_wl
Rw34_24 word34_24 word33_24 R_wl
Cwl_34_24 word34_24 gnd C_wl
Rw35_24 word35_24 word34_24 R_wl
Cwl_35_24 word35_24 gnd C_wl
Rw36_24 word36_24 word35_24 R_wl
Cwl_36_24 word36_24 gnd C_wl
Rw37_24 word37_24 word36_24 R_wl
Cwl_37_24 word37_24 gnd C_wl
Rw38_24 word38_24 word37_24 R_wl
Cwl_38_24 word38_24 gnd C_wl
Rw39_24 word39_24 word38_24 R_wl
Cwl_39_24 word39_24 gnd C_wl
Rw40_24 word40_24 word39_24 R_wl
Cwl_40_24 word40_24 gnd C_wl
Rw41_24 word41_24 word40_24 R_wl
Cwl_41_24 word41_24 gnd C_wl
Rw42_24 word42_24 word41_24 R_wl
Cwl_42_24 word42_24 gnd C_wl
Rw43_24 word43_24 word42_24 R_wl
Cwl_43_24 word43_24 gnd C_wl
Rw44_24 word44_24 word43_24 R_wl
Cwl_44_24 word44_24 gnd C_wl
Rw45_24 word45_24 word44_24 R_wl
Cwl_45_24 word45_24 gnd C_wl
Rw46_24 word46_24 word45_24 R_wl
Cwl_46_24 word46_24 gnd C_wl
Rw47_24 word47_24 word46_24 R_wl
Cwl_47_24 word47_24 gnd C_wl
Rw48_24 word48_24 word47_24 R_wl
Cwl_48_24 word48_24 gnd C_wl
Rw49_24 word49_24 word48_24 R_wl
Cwl_49_24 word49_24 gnd C_wl
Rw50_24 word50_24 word49_24 R_wl
Cwl_50_24 word50_24 gnd C_wl
Rw51_24 word51_24 word50_24 R_wl
Cwl_51_24 word51_24 gnd C_wl
Rw52_24 word52_24 word51_24 R_wl
Cwl_52_24 word52_24 gnd C_wl
Rw53_24 word53_24 word52_24 R_wl
Cwl_53_24 word53_24 gnd C_wl
Rw54_24 word54_24 word53_24 R_wl
Cwl_54_24 word54_24 gnd C_wl
Rw55_24 word55_24 word54_24 R_wl
Cwl_55_24 word55_24 gnd C_wl
Rw56_24 word56_24 word55_24 R_wl
Cwl_56_24 word56_24 gnd C_wl
Rw57_24 word57_24 word56_24 R_wl
Cwl_57_24 word57_24 gnd C_wl
Rw58_24 word58_24 word57_24 R_wl
Cwl_58_24 word58_24 gnd C_wl
Rw59_24 word59_24 word58_24 R_wl
Cwl_59_24 word59_24 gnd C_wl
Rw60_24 word60_24 word59_24 R_wl
Cwl_60_24 word60_24 gnd C_wl
Rw61_24 word61_24 word60_24 R_wl
Cwl_61_24 word61_24 gnd C_wl
Rw62_24 word62_24 word61_24 R_wl
Cwl_62_24 word62_24 gnd C_wl
Rw63_24 word63_24 word62_24 R_wl
Cwl_63_24 word63_24 gnd C_wl
Rw64_24 word64_24 word63_24 R_wl
Cwl_64_24 word64_24 gnd C_wl
Rw65_24 word65_24 word64_24 R_wl
Cwl_65_24 word65_24 gnd C_wl
Rw66_24 word66_24 word65_24 R_wl
Cwl_66_24 word66_24 gnd C_wl
Rw67_24 word67_24 word66_24 R_wl
Cwl_67_24 word67_24 gnd C_wl
Rw68_24 word68_24 word67_24 R_wl
Cwl_68_24 word68_24 gnd C_wl
Rw69_24 word69_24 word68_24 R_wl
Cwl_69_24 word69_24 gnd C_wl
Rw70_24 word70_24 word69_24 R_wl
Cwl_70_24 word70_24 gnd C_wl
Rw71_24 word71_24 word70_24 R_wl
Cwl_71_24 word71_24 gnd C_wl
Rw72_24 word72_24 word71_24 R_wl
Cwl_72_24 word72_24 gnd C_wl
Rw73_24 word73_24 word72_24 R_wl
Cwl_73_24 word73_24 gnd C_wl
Rw74_24 word74_24 word73_24 R_wl
Cwl_74_24 word74_24 gnd C_wl
Rw75_24 word75_24 word74_24 R_wl
Cwl_75_24 word75_24 gnd C_wl
Rw76_24 word76_24 word75_24 R_wl
Cwl_76_24 word76_24 gnd C_wl
Rw77_24 word77_24 word76_24 R_wl
Cwl_77_24 word77_24 gnd C_wl
Rw78_24 word78_24 word77_24 R_wl
Cwl_78_24 word78_24 gnd C_wl
Rw79_24 word79_24 word78_24 R_wl
Cwl_79_24 word79_24 gnd C_wl
Rw80_24 word80_24 word79_24 R_wl
Cwl_80_24 word80_24 gnd C_wl
Rw81_24 word81_24 word80_24 R_wl
Cwl_81_24 word81_24 gnd C_wl
Rw82_24 word82_24 word81_24 R_wl
Cwl_82_24 word82_24 gnd C_wl
Rw83_24 word83_24 word82_24 R_wl
Cwl_83_24 word83_24 gnd C_wl
Rw84_24 word84_24 word83_24 R_wl
Cwl_84_24 word84_24 gnd C_wl
Rw85_24 word85_24 word84_24 R_wl
Cwl_85_24 word85_24 gnd C_wl
Rw86_24 word86_24 word85_24 R_wl
Cwl_86_24 word86_24 gnd C_wl
Rw87_24 word87_24 word86_24 R_wl
Cwl_87_24 word87_24 gnd C_wl
Rw88_24 word88_24 word87_24 R_wl
Cwl_88_24 word88_24 gnd C_wl
Rw89_24 word89_24 word88_24 R_wl
Cwl_89_24 word89_24 gnd C_wl
Rw90_24 word90_24 word89_24 R_wl
Cwl_90_24 word90_24 gnd C_wl
Rw91_24 word91_24 word90_24 R_wl
Cwl_91_24 word91_24 gnd C_wl
Rw92_24 word92_24 word91_24 R_wl
Cwl_92_24 word92_24 gnd C_wl
Rw93_24 word93_24 word92_24 R_wl
Cwl_93_24 word93_24 gnd C_wl
Rw94_24 word94_24 word93_24 R_wl
Cwl_94_24 word94_24 gnd C_wl
Rw95_24 word95_24 word94_24 R_wl
Cwl_95_24 word95_24 gnd C_wl
Rw96_24 word96_24 word95_24 R_wl
Cwl_96_24 word96_24 gnd C_wl
Rw97_24 word97_24 word96_24 R_wl
Cwl_97_24 word97_24 gnd C_wl
Rw98_24 word98_24 word97_24 R_wl
Cwl_98_24 word98_24 gnd C_wl
Rw99_24 word99_24 word98_24 R_wl
Cwl_99_24 word99_24 gnd C_wl
Vwl_25 word_25 0 0
Rw0_25 word_25 word0_25 R_wl
Cwl_0_25 word0_25 gnd C_wl
Rw1_25 word1_25 word0_25 R_wl
Cwl_1_25 word1_25 gnd C_wl
Rw2_25 word2_25 word1_25 R_wl
Cwl_2_25 word2_25 gnd C_wl
Rw3_25 word3_25 word2_25 R_wl
Cwl_3_25 word3_25 gnd C_wl
Rw4_25 word4_25 word3_25 R_wl
Cwl_4_25 word4_25 gnd C_wl
Rw5_25 word5_25 word4_25 R_wl
Cwl_5_25 word5_25 gnd C_wl
Rw6_25 word6_25 word5_25 R_wl
Cwl_6_25 word6_25 gnd C_wl
Rw7_25 word7_25 word6_25 R_wl
Cwl_7_25 word7_25 gnd C_wl
Rw8_25 word8_25 word7_25 R_wl
Cwl_8_25 word8_25 gnd C_wl
Rw9_25 word9_25 word8_25 R_wl
Cwl_9_25 word9_25 gnd C_wl
Rw10_25 word10_25 word9_25 R_wl
Cwl_10_25 word10_25 gnd C_wl
Rw11_25 word11_25 word10_25 R_wl
Cwl_11_25 word11_25 gnd C_wl
Rw12_25 word12_25 word11_25 R_wl
Cwl_12_25 word12_25 gnd C_wl
Rw13_25 word13_25 word12_25 R_wl
Cwl_13_25 word13_25 gnd C_wl
Rw14_25 word14_25 word13_25 R_wl
Cwl_14_25 word14_25 gnd C_wl
Rw15_25 word15_25 word14_25 R_wl
Cwl_15_25 word15_25 gnd C_wl
Rw16_25 word16_25 word15_25 R_wl
Cwl_16_25 word16_25 gnd C_wl
Rw17_25 word17_25 word16_25 R_wl
Cwl_17_25 word17_25 gnd C_wl
Rw18_25 word18_25 word17_25 R_wl
Cwl_18_25 word18_25 gnd C_wl
Rw19_25 word19_25 word18_25 R_wl
Cwl_19_25 word19_25 gnd C_wl
Rw20_25 word20_25 word19_25 R_wl
Cwl_20_25 word20_25 gnd C_wl
Rw21_25 word21_25 word20_25 R_wl
Cwl_21_25 word21_25 gnd C_wl
Rw22_25 word22_25 word21_25 R_wl
Cwl_22_25 word22_25 gnd C_wl
Rw23_25 word23_25 word22_25 R_wl
Cwl_23_25 word23_25 gnd C_wl
Rw24_25 word24_25 word23_25 R_wl
Cwl_24_25 word24_25 gnd C_wl
Rw25_25 word25_25 word24_25 R_wl
Cwl_25_25 word25_25 gnd C_wl
Rw26_25 word26_25 word25_25 R_wl
Cwl_26_25 word26_25 gnd C_wl
Rw27_25 word27_25 word26_25 R_wl
Cwl_27_25 word27_25 gnd C_wl
Rw28_25 word28_25 word27_25 R_wl
Cwl_28_25 word28_25 gnd C_wl
Rw29_25 word29_25 word28_25 R_wl
Cwl_29_25 word29_25 gnd C_wl
Rw30_25 word30_25 word29_25 R_wl
Cwl_30_25 word30_25 gnd C_wl
Rw31_25 word31_25 word30_25 R_wl
Cwl_31_25 word31_25 gnd C_wl
Rw32_25 word32_25 word31_25 R_wl
Cwl_32_25 word32_25 gnd C_wl
Rw33_25 word33_25 word32_25 R_wl
Cwl_33_25 word33_25 gnd C_wl
Rw34_25 word34_25 word33_25 R_wl
Cwl_34_25 word34_25 gnd C_wl
Rw35_25 word35_25 word34_25 R_wl
Cwl_35_25 word35_25 gnd C_wl
Rw36_25 word36_25 word35_25 R_wl
Cwl_36_25 word36_25 gnd C_wl
Rw37_25 word37_25 word36_25 R_wl
Cwl_37_25 word37_25 gnd C_wl
Rw38_25 word38_25 word37_25 R_wl
Cwl_38_25 word38_25 gnd C_wl
Rw39_25 word39_25 word38_25 R_wl
Cwl_39_25 word39_25 gnd C_wl
Rw40_25 word40_25 word39_25 R_wl
Cwl_40_25 word40_25 gnd C_wl
Rw41_25 word41_25 word40_25 R_wl
Cwl_41_25 word41_25 gnd C_wl
Rw42_25 word42_25 word41_25 R_wl
Cwl_42_25 word42_25 gnd C_wl
Rw43_25 word43_25 word42_25 R_wl
Cwl_43_25 word43_25 gnd C_wl
Rw44_25 word44_25 word43_25 R_wl
Cwl_44_25 word44_25 gnd C_wl
Rw45_25 word45_25 word44_25 R_wl
Cwl_45_25 word45_25 gnd C_wl
Rw46_25 word46_25 word45_25 R_wl
Cwl_46_25 word46_25 gnd C_wl
Rw47_25 word47_25 word46_25 R_wl
Cwl_47_25 word47_25 gnd C_wl
Rw48_25 word48_25 word47_25 R_wl
Cwl_48_25 word48_25 gnd C_wl
Rw49_25 word49_25 word48_25 R_wl
Cwl_49_25 word49_25 gnd C_wl
Rw50_25 word50_25 word49_25 R_wl
Cwl_50_25 word50_25 gnd C_wl
Rw51_25 word51_25 word50_25 R_wl
Cwl_51_25 word51_25 gnd C_wl
Rw52_25 word52_25 word51_25 R_wl
Cwl_52_25 word52_25 gnd C_wl
Rw53_25 word53_25 word52_25 R_wl
Cwl_53_25 word53_25 gnd C_wl
Rw54_25 word54_25 word53_25 R_wl
Cwl_54_25 word54_25 gnd C_wl
Rw55_25 word55_25 word54_25 R_wl
Cwl_55_25 word55_25 gnd C_wl
Rw56_25 word56_25 word55_25 R_wl
Cwl_56_25 word56_25 gnd C_wl
Rw57_25 word57_25 word56_25 R_wl
Cwl_57_25 word57_25 gnd C_wl
Rw58_25 word58_25 word57_25 R_wl
Cwl_58_25 word58_25 gnd C_wl
Rw59_25 word59_25 word58_25 R_wl
Cwl_59_25 word59_25 gnd C_wl
Rw60_25 word60_25 word59_25 R_wl
Cwl_60_25 word60_25 gnd C_wl
Rw61_25 word61_25 word60_25 R_wl
Cwl_61_25 word61_25 gnd C_wl
Rw62_25 word62_25 word61_25 R_wl
Cwl_62_25 word62_25 gnd C_wl
Rw63_25 word63_25 word62_25 R_wl
Cwl_63_25 word63_25 gnd C_wl
Rw64_25 word64_25 word63_25 R_wl
Cwl_64_25 word64_25 gnd C_wl
Rw65_25 word65_25 word64_25 R_wl
Cwl_65_25 word65_25 gnd C_wl
Rw66_25 word66_25 word65_25 R_wl
Cwl_66_25 word66_25 gnd C_wl
Rw67_25 word67_25 word66_25 R_wl
Cwl_67_25 word67_25 gnd C_wl
Rw68_25 word68_25 word67_25 R_wl
Cwl_68_25 word68_25 gnd C_wl
Rw69_25 word69_25 word68_25 R_wl
Cwl_69_25 word69_25 gnd C_wl
Rw70_25 word70_25 word69_25 R_wl
Cwl_70_25 word70_25 gnd C_wl
Rw71_25 word71_25 word70_25 R_wl
Cwl_71_25 word71_25 gnd C_wl
Rw72_25 word72_25 word71_25 R_wl
Cwl_72_25 word72_25 gnd C_wl
Rw73_25 word73_25 word72_25 R_wl
Cwl_73_25 word73_25 gnd C_wl
Rw74_25 word74_25 word73_25 R_wl
Cwl_74_25 word74_25 gnd C_wl
Rw75_25 word75_25 word74_25 R_wl
Cwl_75_25 word75_25 gnd C_wl
Rw76_25 word76_25 word75_25 R_wl
Cwl_76_25 word76_25 gnd C_wl
Rw77_25 word77_25 word76_25 R_wl
Cwl_77_25 word77_25 gnd C_wl
Rw78_25 word78_25 word77_25 R_wl
Cwl_78_25 word78_25 gnd C_wl
Rw79_25 word79_25 word78_25 R_wl
Cwl_79_25 word79_25 gnd C_wl
Rw80_25 word80_25 word79_25 R_wl
Cwl_80_25 word80_25 gnd C_wl
Rw81_25 word81_25 word80_25 R_wl
Cwl_81_25 word81_25 gnd C_wl
Rw82_25 word82_25 word81_25 R_wl
Cwl_82_25 word82_25 gnd C_wl
Rw83_25 word83_25 word82_25 R_wl
Cwl_83_25 word83_25 gnd C_wl
Rw84_25 word84_25 word83_25 R_wl
Cwl_84_25 word84_25 gnd C_wl
Rw85_25 word85_25 word84_25 R_wl
Cwl_85_25 word85_25 gnd C_wl
Rw86_25 word86_25 word85_25 R_wl
Cwl_86_25 word86_25 gnd C_wl
Rw87_25 word87_25 word86_25 R_wl
Cwl_87_25 word87_25 gnd C_wl
Rw88_25 word88_25 word87_25 R_wl
Cwl_88_25 word88_25 gnd C_wl
Rw89_25 word89_25 word88_25 R_wl
Cwl_89_25 word89_25 gnd C_wl
Rw90_25 word90_25 word89_25 R_wl
Cwl_90_25 word90_25 gnd C_wl
Rw91_25 word91_25 word90_25 R_wl
Cwl_91_25 word91_25 gnd C_wl
Rw92_25 word92_25 word91_25 R_wl
Cwl_92_25 word92_25 gnd C_wl
Rw93_25 word93_25 word92_25 R_wl
Cwl_93_25 word93_25 gnd C_wl
Rw94_25 word94_25 word93_25 R_wl
Cwl_94_25 word94_25 gnd C_wl
Rw95_25 word95_25 word94_25 R_wl
Cwl_95_25 word95_25 gnd C_wl
Rw96_25 word96_25 word95_25 R_wl
Cwl_96_25 word96_25 gnd C_wl
Rw97_25 word97_25 word96_25 R_wl
Cwl_97_25 word97_25 gnd C_wl
Rw98_25 word98_25 word97_25 R_wl
Cwl_98_25 word98_25 gnd C_wl
Rw99_25 word99_25 word98_25 R_wl
Cwl_99_25 word99_25 gnd C_wl
Vwl_26 word_26 0 0
Rw0_26 word_26 word0_26 R_wl
Cwl_0_26 word0_26 gnd C_wl
Rw1_26 word1_26 word0_26 R_wl
Cwl_1_26 word1_26 gnd C_wl
Rw2_26 word2_26 word1_26 R_wl
Cwl_2_26 word2_26 gnd C_wl
Rw3_26 word3_26 word2_26 R_wl
Cwl_3_26 word3_26 gnd C_wl
Rw4_26 word4_26 word3_26 R_wl
Cwl_4_26 word4_26 gnd C_wl
Rw5_26 word5_26 word4_26 R_wl
Cwl_5_26 word5_26 gnd C_wl
Rw6_26 word6_26 word5_26 R_wl
Cwl_6_26 word6_26 gnd C_wl
Rw7_26 word7_26 word6_26 R_wl
Cwl_7_26 word7_26 gnd C_wl
Rw8_26 word8_26 word7_26 R_wl
Cwl_8_26 word8_26 gnd C_wl
Rw9_26 word9_26 word8_26 R_wl
Cwl_9_26 word9_26 gnd C_wl
Rw10_26 word10_26 word9_26 R_wl
Cwl_10_26 word10_26 gnd C_wl
Rw11_26 word11_26 word10_26 R_wl
Cwl_11_26 word11_26 gnd C_wl
Rw12_26 word12_26 word11_26 R_wl
Cwl_12_26 word12_26 gnd C_wl
Rw13_26 word13_26 word12_26 R_wl
Cwl_13_26 word13_26 gnd C_wl
Rw14_26 word14_26 word13_26 R_wl
Cwl_14_26 word14_26 gnd C_wl
Rw15_26 word15_26 word14_26 R_wl
Cwl_15_26 word15_26 gnd C_wl
Rw16_26 word16_26 word15_26 R_wl
Cwl_16_26 word16_26 gnd C_wl
Rw17_26 word17_26 word16_26 R_wl
Cwl_17_26 word17_26 gnd C_wl
Rw18_26 word18_26 word17_26 R_wl
Cwl_18_26 word18_26 gnd C_wl
Rw19_26 word19_26 word18_26 R_wl
Cwl_19_26 word19_26 gnd C_wl
Rw20_26 word20_26 word19_26 R_wl
Cwl_20_26 word20_26 gnd C_wl
Rw21_26 word21_26 word20_26 R_wl
Cwl_21_26 word21_26 gnd C_wl
Rw22_26 word22_26 word21_26 R_wl
Cwl_22_26 word22_26 gnd C_wl
Rw23_26 word23_26 word22_26 R_wl
Cwl_23_26 word23_26 gnd C_wl
Rw24_26 word24_26 word23_26 R_wl
Cwl_24_26 word24_26 gnd C_wl
Rw25_26 word25_26 word24_26 R_wl
Cwl_25_26 word25_26 gnd C_wl
Rw26_26 word26_26 word25_26 R_wl
Cwl_26_26 word26_26 gnd C_wl
Rw27_26 word27_26 word26_26 R_wl
Cwl_27_26 word27_26 gnd C_wl
Rw28_26 word28_26 word27_26 R_wl
Cwl_28_26 word28_26 gnd C_wl
Rw29_26 word29_26 word28_26 R_wl
Cwl_29_26 word29_26 gnd C_wl
Rw30_26 word30_26 word29_26 R_wl
Cwl_30_26 word30_26 gnd C_wl
Rw31_26 word31_26 word30_26 R_wl
Cwl_31_26 word31_26 gnd C_wl
Rw32_26 word32_26 word31_26 R_wl
Cwl_32_26 word32_26 gnd C_wl
Rw33_26 word33_26 word32_26 R_wl
Cwl_33_26 word33_26 gnd C_wl
Rw34_26 word34_26 word33_26 R_wl
Cwl_34_26 word34_26 gnd C_wl
Rw35_26 word35_26 word34_26 R_wl
Cwl_35_26 word35_26 gnd C_wl
Rw36_26 word36_26 word35_26 R_wl
Cwl_36_26 word36_26 gnd C_wl
Rw37_26 word37_26 word36_26 R_wl
Cwl_37_26 word37_26 gnd C_wl
Rw38_26 word38_26 word37_26 R_wl
Cwl_38_26 word38_26 gnd C_wl
Rw39_26 word39_26 word38_26 R_wl
Cwl_39_26 word39_26 gnd C_wl
Rw40_26 word40_26 word39_26 R_wl
Cwl_40_26 word40_26 gnd C_wl
Rw41_26 word41_26 word40_26 R_wl
Cwl_41_26 word41_26 gnd C_wl
Rw42_26 word42_26 word41_26 R_wl
Cwl_42_26 word42_26 gnd C_wl
Rw43_26 word43_26 word42_26 R_wl
Cwl_43_26 word43_26 gnd C_wl
Rw44_26 word44_26 word43_26 R_wl
Cwl_44_26 word44_26 gnd C_wl
Rw45_26 word45_26 word44_26 R_wl
Cwl_45_26 word45_26 gnd C_wl
Rw46_26 word46_26 word45_26 R_wl
Cwl_46_26 word46_26 gnd C_wl
Rw47_26 word47_26 word46_26 R_wl
Cwl_47_26 word47_26 gnd C_wl
Rw48_26 word48_26 word47_26 R_wl
Cwl_48_26 word48_26 gnd C_wl
Rw49_26 word49_26 word48_26 R_wl
Cwl_49_26 word49_26 gnd C_wl
Rw50_26 word50_26 word49_26 R_wl
Cwl_50_26 word50_26 gnd C_wl
Rw51_26 word51_26 word50_26 R_wl
Cwl_51_26 word51_26 gnd C_wl
Rw52_26 word52_26 word51_26 R_wl
Cwl_52_26 word52_26 gnd C_wl
Rw53_26 word53_26 word52_26 R_wl
Cwl_53_26 word53_26 gnd C_wl
Rw54_26 word54_26 word53_26 R_wl
Cwl_54_26 word54_26 gnd C_wl
Rw55_26 word55_26 word54_26 R_wl
Cwl_55_26 word55_26 gnd C_wl
Rw56_26 word56_26 word55_26 R_wl
Cwl_56_26 word56_26 gnd C_wl
Rw57_26 word57_26 word56_26 R_wl
Cwl_57_26 word57_26 gnd C_wl
Rw58_26 word58_26 word57_26 R_wl
Cwl_58_26 word58_26 gnd C_wl
Rw59_26 word59_26 word58_26 R_wl
Cwl_59_26 word59_26 gnd C_wl
Rw60_26 word60_26 word59_26 R_wl
Cwl_60_26 word60_26 gnd C_wl
Rw61_26 word61_26 word60_26 R_wl
Cwl_61_26 word61_26 gnd C_wl
Rw62_26 word62_26 word61_26 R_wl
Cwl_62_26 word62_26 gnd C_wl
Rw63_26 word63_26 word62_26 R_wl
Cwl_63_26 word63_26 gnd C_wl
Rw64_26 word64_26 word63_26 R_wl
Cwl_64_26 word64_26 gnd C_wl
Rw65_26 word65_26 word64_26 R_wl
Cwl_65_26 word65_26 gnd C_wl
Rw66_26 word66_26 word65_26 R_wl
Cwl_66_26 word66_26 gnd C_wl
Rw67_26 word67_26 word66_26 R_wl
Cwl_67_26 word67_26 gnd C_wl
Rw68_26 word68_26 word67_26 R_wl
Cwl_68_26 word68_26 gnd C_wl
Rw69_26 word69_26 word68_26 R_wl
Cwl_69_26 word69_26 gnd C_wl
Rw70_26 word70_26 word69_26 R_wl
Cwl_70_26 word70_26 gnd C_wl
Rw71_26 word71_26 word70_26 R_wl
Cwl_71_26 word71_26 gnd C_wl
Rw72_26 word72_26 word71_26 R_wl
Cwl_72_26 word72_26 gnd C_wl
Rw73_26 word73_26 word72_26 R_wl
Cwl_73_26 word73_26 gnd C_wl
Rw74_26 word74_26 word73_26 R_wl
Cwl_74_26 word74_26 gnd C_wl
Rw75_26 word75_26 word74_26 R_wl
Cwl_75_26 word75_26 gnd C_wl
Rw76_26 word76_26 word75_26 R_wl
Cwl_76_26 word76_26 gnd C_wl
Rw77_26 word77_26 word76_26 R_wl
Cwl_77_26 word77_26 gnd C_wl
Rw78_26 word78_26 word77_26 R_wl
Cwl_78_26 word78_26 gnd C_wl
Rw79_26 word79_26 word78_26 R_wl
Cwl_79_26 word79_26 gnd C_wl
Rw80_26 word80_26 word79_26 R_wl
Cwl_80_26 word80_26 gnd C_wl
Rw81_26 word81_26 word80_26 R_wl
Cwl_81_26 word81_26 gnd C_wl
Rw82_26 word82_26 word81_26 R_wl
Cwl_82_26 word82_26 gnd C_wl
Rw83_26 word83_26 word82_26 R_wl
Cwl_83_26 word83_26 gnd C_wl
Rw84_26 word84_26 word83_26 R_wl
Cwl_84_26 word84_26 gnd C_wl
Rw85_26 word85_26 word84_26 R_wl
Cwl_85_26 word85_26 gnd C_wl
Rw86_26 word86_26 word85_26 R_wl
Cwl_86_26 word86_26 gnd C_wl
Rw87_26 word87_26 word86_26 R_wl
Cwl_87_26 word87_26 gnd C_wl
Rw88_26 word88_26 word87_26 R_wl
Cwl_88_26 word88_26 gnd C_wl
Rw89_26 word89_26 word88_26 R_wl
Cwl_89_26 word89_26 gnd C_wl
Rw90_26 word90_26 word89_26 R_wl
Cwl_90_26 word90_26 gnd C_wl
Rw91_26 word91_26 word90_26 R_wl
Cwl_91_26 word91_26 gnd C_wl
Rw92_26 word92_26 word91_26 R_wl
Cwl_92_26 word92_26 gnd C_wl
Rw93_26 word93_26 word92_26 R_wl
Cwl_93_26 word93_26 gnd C_wl
Rw94_26 word94_26 word93_26 R_wl
Cwl_94_26 word94_26 gnd C_wl
Rw95_26 word95_26 word94_26 R_wl
Cwl_95_26 word95_26 gnd C_wl
Rw96_26 word96_26 word95_26 R_wl
Cwl_96_26 word96_26 gnd C_wl
Rw97_26 word97_26 word96_26 R_wl
Cwl_97_26 word97_26 gnd C_wl
Rw98_26 word98_26 word97_26 R_wl
Cwl_98_26 word98_26 gnd C_wl
Rw99_26 word99_26 word98_26 R_wl
Cwl_99_26 word99_26 gnd C_wl
Vwl_27 word_27 0 0
Rw0_27 word_27 word0_27 R_wl
Cwl_0_27 word0_27 gnd C_wl
Rw1_27 word1_27 word0_27 R_wl
Cwl_1_27 word1_27 gnd C_wl
Rw2_27 word2_27 word1_27 R_wl
Cwl_2_27 word2_27 gnd C_wl
Rw3_27 word3_27 word2_27 R_wl
Cwl_3_27 word3_27 gnd C_wl
Rw4_27 word4_27 word3_27 R_wl
Cwl_4_27 word4_27 gnd C_wl
Rw5_27 word5_27 word4_27 R_wl
Cwl_5_27 word5_27 gnd C_wl
Rw6_27 word6_27 word5_27 R_wl
Cwl_6_27 word6_27 gnd C_wl
Rw7_27 word7_27 word6_27 R_wl
Cwl_7_27 word7_27 gnd C_wl
Rw8_27 word8_27 word7_27 R_wl
Cwl_8_27 word8_27 gnd C_wl
Rw9_27 word9_27 word8_27 R_wl
Cwl_9_27 word9_27 gnd C_wl
Rw10_27 word10_27 word9_27 R_wl
Cwl_10_27 word10_27 gnd C_wl
Rw11_27 word11_27 word10_27 R_wl
Cwl_11_27 word11_27 gnd C_wl
Rw12_27 word12_27 word11_27 R_wl
Cwl_12_27 word12_27 gnd C_wl
Rw13_27 word13_27 word12_27 R_wl
Cwl_13_27 word13_27 gnd C_wl
Rw14_27 word14_27 word13_27 R_wl
Cwl_14_27 word14_27 gnd C_wl
Rw15_27 word15_27 word14_27 R_wl
Cwl_15_27 word15_27 gnd C_wl
Rw16_27 word16_27 word15_27 R_wl
Cwl_16_27 word16_27 gnd C_wl
Rw17_27 word17_27 word16_27 R_wl
Cwl_17_27 word17_27 gnd C_wl
Rw18_27 word18_27 word17_27 R_wl
Cwl_18_27 word18_27 gnd C_wl
Rw19_27 word19_27 word18_27 R_wl
Cwl_19_27 word19_27 gnd C_wl
Rw20_27 word20_27 word19_27 R_wl
Cwl_20_27 word20_27 gnd C_wl
Rw21_27 word21_27 word20_27 R_wl
Cwl_21_27 word21_27 gnd C_wl
Rw22_27 word22_27 word21_27 R_wl
Cwl_22_27 word22_27 gnd C_wl
Rw23_27 word23_27 word22_27 R_wl
Cwl_23_27 word23_27 gnd C_wl
Rw24_27 word24_27 word23_27 R_wl
Cwl_24_27 word24_27 gnd C_wl
Rw25_27 word25_27 word24_27 R_wl
Cwl_25_27 word25_27 gnd C_wl
Rw26_27 word26_27 word25_27 R_wl
Cwl_26_27 word26_27 gnd C_wl
Rw27_27 word27_27 word26_27 R_wl
Cwl_27_27 word27_27 gnd C_wl
Rw28_27 word28_27 word27_27 R_wl
Cwl_28_27 word28_27 gnd C_wl
Rw29_27 word29_27 word28_27 R_wl
Cwl_29_27 word29_27 gnd C_wl
Rw30_27 word30_27 word29_27 R_wl
Cwl_30_27 word30_27 gnd C_wl
Rw31_27 word31_27 word30_27 R_wl
Cwl_31_27 word31_27 gnd C_wl
Rw32_27 word32_27 word31_27 R_wl
Cwl_32_27 word32_27 gnd C_wl
Rw33_27 word33_27 word32_27 R_wl
Cwl_33_27 word33_27 gnd C_wl
Rw34_27 word34_27 word33_27 R_wl
Cwl_34_27 word34_27 gnd C_wl
Rw35_27 word35_27 word34_27 R_wl
Cwl_35_27 word35_27 gnd C_wl
Rw36_27 word36_27 word35_27 R_wl
Cwl_36_27 word36_27 gnd C_wl
Rw37_27 word37_27 word36_27 R_wl
Cwl_37_27 word37_27 gnd C_wl
Rw38_27 word38_27 word37_27 R_wl
Cwl_38_27 word38_27 gnd C_wl
Rw39_27 word39_27 word38_27 R_wl
Cwl_39_27 word39_27 gnd C_wl
Rw40_27 word40_27 word39_27 R_wl
Cwl_40_27 word40_27 gnd C_wl
Rw41_27 word41_27 word40_27 R_wl
Cwl_41_27 word41_27 gnd C_wl
Rw42_27 word42_27 word41_27 R_wl
Cwl_42_27 word42_27 gnd C_wl
Rw43_27 word43_27 word42_27 R_wl
Cwl_43_27 word43_27 gnd C_wl
Rw44_27 word44_27 word43_27 R_wl
Cwl_44_27 word44_27 gnd C_wl
Rw45_27 word45_27 word44_27 R_wl
Cwl_45_27 word45_27 gnd C_wl
Rw46_27 word46_27 word45_27 R_wl
Cwl_46_27 word46_27 gnd C_wl
Rw47_27 word47_27 word46_27 R_wl
Cwl_47_27 word47_27 gnd C_wl
Rw48_27 word48_27 word47_27 R_wl
Cwl_48_27 word48_27 gnd C_wl
Rw49_27 word49_27 word48_27 R_wl
Cwl_49_27 word49_27 gnd C_wl
Rw50_27 word50_27 word49_27 R_wl
Cwl_50_27 word50_27 gnd C_wl
Rw51_27 word51_27 word50_27 R_wl
Cwl_51_27 word51_27 gnd C_wl
Rw52_27 word52_27 word51_27 R_wl
Cwl_52_27 word52_27 gnd C_wl
Rw53_27 word53_27 word52_27 R_wl
Cwl_53_27 word53_27 gnd C_wl
Rw54_27 word54_27 word53_27 R_wl
Cwl_54_27 word54_27 gnd C_wl
Rw55_27 word55_27 word54_27 R_wl
Cwl_55_27 word55_27 gnd C_wl
Rw56_27 word56_27 word55_27 R_wl
Cwl_56_27 word56_27 gnd C_wl
Rw57_27 word57_27 word56_27 R_wl
Cwl_57_27 word57_27 gnd C_wl
Rw58_27 word58_27 word57_27 R_wl
Cwl_58_27 word58_27 gnd C_wl
Rw59_27 word59_27 word58_27 R_wl
Cwl_59_27 word59_27 gnd C_wl
Rw60_27 word60_27 word59_27 R_wl
Cwl_60_27 word60_27 gnd C_wl
Rw61_27 word61_27 word60_27 R_wl
Cwl_61_27 word61_27 gnd C_wl
Rw62_27 word62_27 word61_27 R_wl
Cwl_62_27 word62_27 gnd C_wl
Rw63_27 word63_27 word62_27 R_wl
Cwl_63_27 word63_27 gnd C_wl
Rw64_27 word64_27 word63_27 R_wl
Cwl_64_27 word64_27 gnd C_wl
Rw65_27 word65_27 word64_27 R_wl
Cwl_65_27 word65_27 gnd C_wl
Rw66_27 word66_27 word65_27 R_wl
Cwl_66_27 word66_27 gnd C_wl
Rw67_27 word67_27 word66_27 R_wl
Cwl_67_27 word67_27 gnd C_wl
Rw68_27 word68_27 word67_27 R_wl
Cwl_68_27 word68_27 gnd C_wl
Rw69_27 word69_27 word68_27 R_wl
Cwl_69_27 word69_27 gnd C_wl
Rw70_27 word70_27 word69_27 R_wl
Cwl_70_27 word70_27 gnd C_wl
Rw71_27 word71_27 word70_27 R_wl
Cwl_71_27 word71_27 gnd C_wl
Rw72_27 word72_27 word71_27 R_wl
Cwl_72_27 word72_27 gnd C_wl
Rw73_27 word73_27 word72_27 R_wl
Cwl_73_27 word73_27 gnd C_wl
Rw74_27 word74_27 word73_27 R_wl
Cwl_74_27 word74_27 gnd C_wl
Rw75_27 word75_27 word74_27 R_wl
Cwl_75_27 word75_27 gnd C_wl
Rw76_27 word76_27 word75_27 R_wl
Cwl_76_27 word76_27 gnd C_wl
Rw77_27 word77_27 word76_27 R_wl
Cwl_77_27 word77_27 gnd C_wl
Rw78_27 word78_27 word77_27 R_wl
Cwl_78_27 word78_27 gnd C_wl
Rw79_27 word79_27 word78_27 R_wl
Cwl_79_27 word79_27 gnd C_wl
Rw80_27 word80_27 word79_27 R_wl
Cwl_80_27 word80_27 gnd C_wl
Rw81_27 word81_27 word80_27 R_wl
Cwl_81_27 word81_27 gnd C_wl
Rw82_27 word82_27 word81_27 R_wl
Cwl_82_27 word82_27 gnd C_wl
Rw83_27 word83_27 word82_27 R_wl
Cwl_83_27 word83_27 gnd C_wl
Rw84_27 word84_27 word83_27 R_wl
Cwl_84_27 word84_27 gnd C_wl
Rw85_27 word85_27 word84_27 R_wl
Cwl_85_27 word85_27 gnd C_wl
Rw86_27 word86_27 word85_27 R_wl
Cwl_86_27 word86_27 gnd C_wl
Rw87_27 word87_27 word86_27 R_wl
Cwl_87_27 word87_27 gnd C_wl
Rw88_27 word88_27 word87_27 R_wl
Cwl_88_27 word88_27 gnd C_wl
Rw89_27 word89_27 word88_27 R_wl
Cwl_89_27 word89_27 gnd C_wl
Rw90_27 word90_27 word89_27 R_wl
Cwl_90_27 word90_27 gnd C_wl
Rw91_27 word91_27 word90_27 R_wl
Cwl_91_27 word91_27 gnd C_wl
Rw92_27 word92_27 word91_27 R_wl
Cwl_92_27 word92_27 gnd C_wl
Rw93_27 word93_27 word92_27 R_wl
Cwl_93_27 word93_27 gnd C_wl
Rw94_27 word94_27 word93_27 R_wl
Cwl_94_27 word94_27 gnd C_wl
Rw95_27 word95_27 word94_27 R_wl
Cwl_95_27 word95_27 gnd C_wl
Rw96_27 word96_27 word95_27 R_wl
Cwl_96_27 word96_27 gnd C_wl
Rw97_27 word97_27 word96_27 R_wl
Cwl_97_27 word97_27 gnd C_wl
Rw98_27 word98_27 word97_27 R_wl
Cwl_98_27 word98_27 gnd C_wl
Rw99_27 word99_27 word98_27 R_wl
Cwl_99_27 word99_27 gnd C_wl
Vwl_28 word_28 0 0
Rw0_28 word_28 word0_28 R_wl
Cwl_0_28 word0_28 gnd C_wl
Rw1_28 word1_28 word0_28 R_wl
Cwl_1_28 word1_28 gnd C_wl
Rw2_28 word2_28 word1_28 R_wl
Cwl_2_28 word2_28 gnd C_wl
Rw3_28 word3_28 word2_28 R_wl
Cwl_3_28 word3_28 gnd C_wl
Rw4_28 word4_28 word3_28 R_wl
Cwl_4_28 word4_28 gnd C_wl
Rw5_28 word5_28 word4_28 R_wl
Cwl_5_28 word5_28 gnd C_wl
Rw6_28 word6_28 word5_28 R_wl
Cwl_6_28 word6_28 gnd C_wl
Rw7_28 word7_28 word6_28 R_wl
Cwl_7_28 word7_28 gnd C_wl
Rw8_28 word8_28 word7_28 R_wl
Cwl_8_28 word8_28 gnd C_wl
Rw9_28 word9_28 word8_28 R_wl
Cwl_9_28 word9_28 gnd C_wl
Rw10_28 word10_28 word9_28 R_wl
Cwl_10_28 word10_28 gnd C_wl
Rw11_28 word11_28 word10_28 R_wl
Cwl_11_28 word11_28 gnd C_wl
Rw12_28 word12_28 word11_28 R_wl
Cwl_12_28 word12_28 gnd C_wl
Rw13_28 word13_28 word12_28 R_wl
Cwl_13_28 word13_28 gnd C_wl
Rw14_28 word14_28 word13_28 R_wl
Cwl_14_28 word14_28 gnd C_wl
Rw15_28 word15_28 word14_28 R_wl
Cwl_15_28 word15_28 gnd C_wl
Rw16_28 word16_28 word15_28 R_wl
Cwl_16_28 word16_28 gnd C_wl
Rw17_28 word17_28 word16_28 R_wl
Cwl_17_28 word17_28 gnd C_wl
Rw18_28 word18_28 word17_28 R_wl
Cwl_18_28 word18_28 gnd C_wl
Rw19_28 word19_28 word18_28 R_wl
Cwl_19_28 word19_28 gnd C_wl
Rw20_28 word20_28 word19_28 R_wl
Cwl_20_28 word20_28 gnd C_wl
Rw21_28 word21_28 word20_28 R_wl
Cwl_21_28 word21_28 gnd C_wl
Rw22_28 word22_28 word21_28 R_wl
Cwl_22_28 word22_28 gnd C_wl
Rw23_28 word23_28 word22_28 R_wl
Cwl_23_28 word23_28 gnd C_wl
Rw24_28 word24_28 word23_28 R_wl
Cwl_24_28 word24_28 gnd C_wl
Rw25_28 word25_28 word24_28 R_wl
Cwl_25_28 word25_28 gnd C_wl
Rw26_28 word26_28 word25_28 R_wl
Cwl_26_28 word26_28 gnd C_wl
Rw27_28 word27_28 word26_28 R_wl
Cwl_27_28 word27_28 gnd C_wl
Rw28_28 word28_28 word27_28 R_wl
Cwl_28_28 word28_28 gnd C_wl
Rw29_28 word29_28 word28_28 R_wl
Cwl_29_28 word29_28 gnd C_wl
Rw30_28 word30_28 word29_28 R_wl
Cwl_30_28 word30_28 gnd C_wl
Rw31_28 word31_28 word30_28 R_wl
Cwl_31_28 word31_28 gnd C_wl
Rw32_28 word32_28 word31_28 R_wl
Cwl_32_28 word32_28 gnd C_wl
Rw33_28 word33_28 word32_28 R_wl
Cwl_33_28 word33_28 gnd C_wl
Rw34_28 word34_28 word33_28 R_wl
Cwl_34_28 word34_28 gnd C_wl
Rw35_28 word35_28 word34_28 R_wl
Cwl_35_28 word35_28 gnd C_wl
Rw36_28 word36_28 word35_28 R_wl
Cwl_36_28 word36_28 gnd C_wl
Rw37_28 word37_28 word36_28 R_wl
Cwl_37_28 word37_28 gnd C_wl
Rw38_28 word38_28 word37_28 R_wl
Cwl_38_28 word38_28 gnd C_wl
Rw39_28 word39_28 word38_28 R_wl
Cwl_39_28 word39_28 gnd C_wl
Rw40_28 word40_28 word39_28 R_wl
Cwl_40_28 word40_28 gnd C_wl
Rw41_28 word41_28 word40_28 R_wl
Cwl_41_28 word41_28 gnd C_wl
Rw42_28 word42_28 word41_28 R_wl
Cwl_42_28 word42_28 gnd C_wl
Rw43_28 word43_28 word42_28 R_wl
Cwl_43_28 word43_28 gnd C_wl
Rw44_28 word44_28 word43_28 R_wl
Cwl_44_28 word44_28 gnd C_wl
Rw45_28 word45_28 word44_28 R_wl
Cwl_45_28 word45_28 gnd C_wl
Rw46_28 word46_28 word45_28 R_wl
Cwl_46_28 word46_28 gnd C_wl
Rw47_28 word47_28 word46_28 R_wl
Cwl_47_28 word47_28 gnd C_wl
Rw48_28 word48_28 word47_28 R_wl
Cwl_48_28 word48_28 gnd C_wl
Rw49_28 word49_28 word48_28 R_wl
Cwl_49_28 word49_28 gnd C_wl
Rw50_28 word50_28 word49_28 R_wl
Cwl_50_28 word50_28 gnd C_wl
Rw51_28 word51_28 word50_28 R_wl
Cwl_51_28 word51_28 gnd C_wl
Rw52_28 word52_28 word51_28 R_wl
Cwl_52_28 word52_28 gnd C_wl
Rw53_28 word53_28 word52_28 R_wl
Cwl_53_28 word53_28 gnd C_wl
Rw54_28 word54_28 word53_28 R_wl
Cwl_54_28 word54_28 gnd C_wl
Rw55_28 word55_28 word54_28 R_wl
Cwl_55_28 word55_28 gnd C_wl
Rw56_28 word56_28 word55_28 R_wl
Cwl_56_28 word56_28 gnd C_wl
Rw57_28 word57_28 word56_28 R_wl
Cwl_57_28 word57_28 gnd C_wl
Rw58_28 word58_28 word57_28 R_wl
Cwl_58_28 word58_28 gnd C_wl
Rw59_28 word59_28 word58_28 R_wl
Cwl_59_28 word59_28 gnd C_wl
Rw60_28 word60_28 word59_28 R_wl
Cwl_60_28 word60_28 gnd C_wl
Rw61_28 word61_28 word60_28 R_wl
Cwl_61_28 word61_28 gnd C_wl
Rw62_28 word62_28 word61_28 R_wl
Cwl_62_28 word62_28 gnd C_wl
Rw63_28 word63_28 word62_28 R_wl
Cwl_63_28 word63_28 gnd C_wl
Rw64_28 word64_28 word63_28 R_wl
Cwl_64_28 word64_28 gnd C_wl
Rw65_28 word65_28 word64_28 R_wl
Cwl_65_28 word65_28 gnd C_wl
Rw66_28 word66_28 word65_28 R_wl
Cwl_66_28 word66_28 gnd C_wl
Rw67_28 word67_28 word66_28 R_wl
Cwl_67_28 word67_28 gnd C_wl
Rw68_28 word68_28 word67_28 R_wl
Cwl_68_28 word68_28 gnd C_wl
Rw69_28 word69_28 word68_28 R_wl
Cwl_69_28 word69_28 gnd C_wl
Rw70_28 word70_28 word69_28 R_wl
Cwl_70_28 word70_28 gnd C_wl
Rw71_28 word71_28 word70_28 R_wl
Cwl_71_28 word71_28 gnd C_wl
Rw72_28 word72_28 word71_28 R_wl
Cwl_72_28 word72_28 gnd C_wl
Rw73_28 word73_28 word72_28 R_wl
Cwl_73_28 word73_28 gnd C_wl
Rw74_28 word74_28 word73_28 R_wl
Cwl_74_28 word74_28 gnd C_wl
Rw75_28 word75_28 word74_28 R_wl
Cwl_75_28 word75_28 gnd C_wl
Rw76_28 word76_28 word75_28 R_wl
Cwl_76_28 word76_28 gnd C_wl
Rw77_28 word77_28 word76_28 R_wl
Cwl_77_28 word77_28 gnd C_wl
Rw78_28 word78_28 word77_28 R_wl
Cwl_78_28 word78_28 gnd C_wl
Rw79_28 word79_28 word78_28 R_wl
Cwl_79_28 word79_28 gnd C_wl
Rw80_28 word80_28 word79_28 R_wl
Cwl_80_28 word80_28 gnd C_wl
Rw81_28 word81_28 word80_28 R_wl
Cwl_81_28 word81_28 gnd C_wl
Rw82_28 word82_28 word81_28 R_wl
Cwl_82_28 word82_28 gnd C_wl
Rw83_28 word83_28 word82_28 R_wl
Cwl_83_28 word83_28 gnd C_wl
Rw84_28 word84_28 word83_28 R_wl
Cwl_84_28 word84_28 gnd C_wl
Rw85_28 word85_28 word84_28 R_wl
Cwl_85_28 word85_28 gnd C_wl
Rw86_28 word86_28 word85_28 R_wl
Cwl_86_28 word86_28 gnd C_wl
Rw87_28 word87_28 word86_28 R_wl
Cwl_87_28 word87_28 gnd C_wl
Rw88_28 word88_28 word87_28 R_wl
Cwl_88_28 word88_28 gnd C_wl
Rw89_28 word89_28 word88_28 R_wl
Cwl_89_28 word89_28 gnd C_wl
Rw90_28 word90_28 word89_28 R_wl
Cwl_90_28 word90_28 gnd C_wl
Rw91_28 word91_28 word90_28 R_wl
Cwl_91_28 word91_28 gnd C_wl
Rw92_28 word92_28 word91_28 R_wl
Cwl_92_28 word92_28 gnd C_wl
Rw93_28 word93_28 word92_28 R_wl
Cwl_93_28 word93_28 gnd C_wl
Rw94_28 word94_28 word93_28 R_wl
Cwl_94_28 word94_28 gnd C_wl
Rw95_28 word95_28 word94_28 R_wl
Cwl_95_28 word95_28 gnd C_wl
Rw96_28 word96_28 word95_28 R_wl
Cwl_96_28 word96_28 gnd C_wl
Rw97_28 word97_28 word96_28 R_wl
Cwl_97_28 word97_28 gnd C_wl
Rw98_28 word98_28 word97_28 R_wl
Cwl_98_28 word98_28 gnd C_wl
Rw99_28 word99_28 word98_28 R_wl
Cwl_99_28 word99_28 gnd C_wl
Vwl_29 word_29 0 0
Rw0_29 word_29 word0_29 R_wl
Cwl_0_29 word0_29 gnd C_wl
Rw1_29 word1_29 word0_29 R_wl
Cwl_1_29 word1_29 gnd C_wl
Rw2_29 word2_29 word1_29 R_wl
Cwl_2_29 word2_29 gnd C_wl
Rw3_29 word3_29 word2_29 R_wl
Cwl_3_29 word3_29 gnd C_wl
Rw4_29 word4_29 word3_29 R_wl
Cwl_4_29 word4_29 gnd C_wl
Rw5_29 word5_29 word4_29 R_wl
Cwl_5_29 word5_29 gnd C_wl
Rw6_29 word6_29 word5_29 R_wl
Cwl_6_29 word6_29 gnd C_wl
Rw7_29 word7_29 word6_29 R_wl
Cwl_7_29 word7_29 gnd C_wl
Rw8_29 word8_29 word7_29 R_wl
Cwl_8_29 word8_29 gnd C_wl
Rw9_29 word9_29 word8_29 R_wl
Cwl_9_29 word9_29 gnd C_wl
Rw10_29 word10_29 word9_29 R_wl
Cwl_10_29 word10_29 gnd C_wl
Rw11_29 word11_29 word10_29 R_wl
Cwl_11_29 word11_29 gnd C_wl
Rw12_29 word12_29 word11_29 R_wl
Cwl_12_29 word12_29 gnd C_wl
Rw13_29 word13_29 word12_29 R_wl
Cwl_13_29 word13_29 gnd C_wl
Rw14_29 word14_29 word13_29 R_wl
Cwl_14_29 word14_29 gnd C_wl
Rw15_29 word15_29 word14_29 R_wl
Cwl_15_29 word15_29 gnd C_wl
Rw16_29 word16_29 word15_29 R_wl
Cwl_16_29 word16_29 gnd C_wl
Rw17_29 word17_29 word16_29 R_wl
Cwl_17_29 word17_29 gnd C_wl
Rw18_29 word18_29 word17_29 R_wl
Cwl_18_29 word18_29 gnd C_wl
Rw19_29 word19_29 word18_29 R_wl
Cwl_19_29 word19_29 gnd C_wl
Rw20_29 word20_29 word19_29 R_wl
Cwl_20_29 word20_29 gnd C_wl
Rw21_29 word21_29 word20_29 R_wl
Cwl_21_29 word21_29 gnd C_wl
Rw22_29 word22_29 word21_29 R_wl
Cwl_22_29 word22_29 gnd C_wl
Rw23_29 word23_29 word22_29 R_wl
Cwl_23_29 word23_29 gnd C_wl
Rw24_29 word24_29 word23_29 R_wl
Cwl_24_29 word24_29 gnd C_wl
Rw25_29 word25_29 word24_29 R_wl
Cwl_25_29 word25_29 gnd C_wl
Rw26_29 word26_29 word25_29 R_wl
Cwl_26_29 word26_29 gnd C_wl
Rw27_29 word27_29 word26_29 R_wl
Cwl_27_29 word27_29 gnd C_wl
Rw28_29 word28_29 word27_29 R_wl
Cwl_28_29 word28_29 gnd C_wl
Rw29_29 word29_29 word28_29 R_wl
Cwl_29_29 word29_29 gnd C_wl
Rw30_29 word30_29 word29_29 R_wl
Cwl_30_29 word30_29 gnd C_wl
Rw31_29 word31_29 word30_29 R_wl
Cwl_31_29 word31_29 gnd C_wl
Rw32_29 word32_29 word31_29 R_wl
Cwl_32_29 word32_29 gnd C_wl
Rw33_29 word33_29 word32_29 R_wl
Cwl_33_29 word33_29 gnd C_wl
Rw34_29 word34_29 word33_29 R_wl
Cwl_34_29 word34_29 gnd C_wl
Rw35_29 word35_29 word34_29 R_wl
Cwl_35_29 word35_29 gnd C_wl
Rw36_29 word36_29 word35_29 R_wl
Cwl_36_29 word36_29 gnd C_wl
Rw37_29 word37_29 word36_29 R_wl
Cwl_37_29 word37_29 gnd C_wl
Rw38_29 word38_29 word37_29 R_wl
Cwl_38_29 word38_29 gnd C_wl
Rw39_29 word39_29 word38_29 R_wl
Cwl_39_29 word39_29 gnd C_wl
Rw40_29 word40_29 word39_29 R_wl
Cwl_40_29 word40_29 gnd C_wl
Rw41_29 word41_29 word40_29 R_wl
Cwl_41_29 word41_29 gnd C_wl
Rw42_29 word42_29 word41_29 R_wl
Cwl_42_29 word42_29 gnd C_wl
Rw43_29 word43_29 word42_29 R_wl
Cwl_43_29 word43_29 gnd C_wl
Rw44_29 word44_29 word43_29 R_wl
Cwl_44_29 word44_29 gnd C_wl
Rw45_29 word45_29 word44_29 R_wl
Cwl_45_29 word45_29 gnd C_wl
Rw46_29 word46_29 word45_29 R_wl
Cwl_46_29 word46_29 gnd C_wl
Rw47_29 word47_29 word46_29 R_wl
Cwl_47_29 word47_29 gnd C_wl
Rw48_29 word48_29 word47_29 R_wl
Cwl_48_29 word48_29 gnd C_wl
Rw49_29 word49_29 word48_29 R_wl
Cwl_49_29 word49_29 gnd C_wl
Rw50_29 word50_29 word49_29 R_wl
Cwl_50_29 word50_29 gnd C_wl
Rw51_29 word51_29 word50_29 R_wl
Cwl_51_29 word51_29 gnd C_wl
Rw52_29 word52_29 word51_29 R_wl
Cwl_52_29 word52_29 gnd C_wl
Rw53_29 word53_29 word52_29 R_wl
Cwl_53_29 word53_29 gnd C_wl
Rw54_29 word54_29 word53_29 R_wl
Cwl_54_29 word54_29 gnd C_wl
Rw55_29 word55_29 word54_29 R_wl
Cwl_55_29 word55_29 gnd C_wl
Rw56_29 word56_29 word55_29 R_wl
Cwl_56_29 word56_29 gnd C_wl
Rw57_29 word57_29 word56_29 R_wl
Cwl_57_29 word57_29 gnd C_wl
Rw58_29 word58_29 word57_29 R_wl
Cwl_58_29 word58_29 gnd C_wl
Rw59_29 word59_29 word58_29 R_wl
Cwl_59_29 word59_29 gnd C_wl
Rw60_29 word60_29 word59_29 R_wl
Cwl_60_29 word60_29 gnd C_wl
Rw61_29 word61_29 word60_29 R_wl
Cwl_61_29 word61_29 gnd C_wl
Rw62_29 word62_29 word61_29 R_wl
Cwl_62_29 word62_29 gnd C_wl
Rw63_29 word63_29 word62_29 R_wl
Cwl_63_29 word63_29 gnd C_wl
Rw64_29 word64_29 word63_29 R_wl
Cwl_64_29 word64_29 gnd C_wl
Rw65_29 word65_29 word64_29 R_wl
Cwl_65_29 word65_29 gnd C_wl
Rw66_29 word66_29 word65_29 R_wl
Cwl_66_29 word66_29 gnd C_wl
Rw67_29 word67_29 word66_29 R_wl
Cwl_67_29 word67_29 gnd C_wl
Rw68_29 word68_29 word67_29 R_wl
Cwl_68_29 word68_29 gnd C_wl
Rw69_29 word69_29 word68_29 R_wl
Cwl_69_29 word69_29 gnd C_wl
Rw70_29 word70_29 word69_29 R_wl
Cwl_70_29 word70_29 gnd C_wl
Rw71_29 word71_29 word70_29 R_wl
Cwl_71_29 word71_29 gnd C_wl
Rw72_29 word72_29 word71_29 R_wl
Cwl_72_29 word72_29 gnd C_wl
Rw73_29 word73_29 word72_29 R_wl
Cwl_73_29 word73_29 gnd C_wl
Rw74_29 word74_29 word73_29 R_wl
Cwl_74_29 word74_29 gnd C_wl
Rw75_29 word75_29 word74_29 R_wl
Cwl_75_29 word75_29 gnd C_wl
Rw76_29 word76_29 word75_29 R_wl
Cwl_76_29 word76_29 gnd C_wl
Rw77_29 word77_29 word76_29 R_wl
Cwl_77_29 word77_29 gnd C_wl
Rw78_29 word78_29 word77_29 R_wl
Cwl_78_29 word78_29 gnd C_wl
Rw79_29 word79_29 word78_29 R_wl
Cwl_79_29 word79_29 gnd C_wl
Rw80_29 word80_29 word79_29 R_wl
Cwl_80_29 word80_29 gnd C_wl
Rw81_29 word81_29 word80_29 R_wl
Cwl_81_29 word81_29 gnd C_wl
Rw82_29 word82_29 word81_29 R_wl
Cwl_82_29 word82_29 gnd C_wl
Rw83_29 word83_29 word82_29 R_wl
Cwl_83_29 word83_29 gnd C_wl
Rw84_29 word84_29 word83_29 R_wl
Cwl_84_29 word84_29 gnd C_wl
Rw85_29 word85_29 word84_29 R_wl
Cwl_85_29 word85_29 gnd C_wl
Rw86_29 word86_29 word85_29 R_wl
Cwl_86_29 word86_29 gnd C_wl
Rw87_29 word87_29 word86_29 R_wl
Cwl_87_29 word87_29 gnd C_wl
Rw88_29 word88_29 word87_29 R_wl
Cwl_88_29 word88_29 gnd C_wl
Rw89_29 word89_29 word88_29 R_wl
Cwl_89_29 word89_29 gnd C_wl
Rw90_29 word90_29 word89_29 R_wl
Cwl_90_29 word90_29 gnd C_wl
Rw91_29 word91_29 word90_29 R_wl
Cwl_91_29 word91_29 gnd C_wl
Rw92_29 word92_29 word91_29 R_wl
Cwl_92_29 word92_29 gnd C_wl
Rw93_29 word93_29 word92_29 R_wl
Cwl_93_29 word93_29 gnd C_wl
Rw94_29 word94_29 word93_29 R_wl
Cwl_94_29 word94_29 gnd C_wl
Rw95_29 word95_29 word94_29 R_wl
Cwl_95_29 word95_29 gnd C_wl
Rw96_29 word96_29 word95_29 R_wl
Cwl_96_29 word96_29 gnd C_wl
Rw97_29 word97_29 word96_29 R_wl
Cwl_97_29 word97_29 gnd C_wl
Rw98_29 word98_29 word97_29 R_wl
Cwl_98_29 word98_29 gnd C_wl
Rw99_29 word99_29 word98_29 R_wl
Cwl_99_29 word99_29 gnd C_wl
Vwl_30 word_30 0 0
Rw0_30 word_30 word0_30 R_wl
Cwl_0_30 word0_30 gnd C_wl
Rw1_30 word1_30 word0_30 R_wl
Cwl_1_30 word1_30 gnd C_wl
Rw2_30 word2_30 word1_30 R_wl
Cwl_2_30 word2_30 gnd C_wl
Rw3_30 word3_30 word2_30 R_wl
Cwl_3_30 word3_30 gnd C_wl
Rw4_30 word4_30 word3_30 R_wl
Cwl_4_30 word4_30 gnd C_wl
Rw5_30 word5_30 word4_30 R_wl
Cwl_5_30 word5_30 gnd C_wl
Rw6_30 word6_30 word5_30 R_wl
Cwl_6_30 word6_30 gnd C_wl
Rw7_30 word7_30 word6_30 R_wl
Cwl_7_30 word7_30 gnd C_wl
Rw8_30 word8_30 word7_30 R_wl
Cwl_8_30 word8_30 gnd C_wl
Rw9_30 word9_30 word8_30 R_wl
Cwl_9_30 word9_30 gnd C_wl
Rw10_30 word10_30 word9_30 R_wl
Cwl_10_30 word10_30 gnd C_wl
Rw11_30 word11_30 word10_30 R_wl
Cwl_11_30 word11_30 gnd C_wl
Rw12_30 word12_30 word11_30 R_wl
Cwl_12_30 word12_30 gnd C_wl
Rw13_30 word13_30 word12_30 R_wl
Cwl_13_30 word13_30 gnd C_wl
Rw14_30 word14_30 word13_30 R_wl
Cwl_14_30 word14_30 gnd C_wl
Rw15_30 word15_30 word14_30 R_wl
Cwl_15_30 word15_30 gnd C_wl
Rw16_30 word16_30 word15_30 R_wl
Cwl_16_30 word16_30 gnd C_wl
Rw17_30 word17_30 word16_30 R_wl
Cwl_17_30 word17_30 gnd C_wl
Rw18_30 word18_30 word17_30 R_wl
Cwl_18_30 word18_30 gnd C_wl
Rw19_30 word19_30 word18_30 R_wl
Cwl_19_30 word19_30 gnd C_wl
Rw20_30 word20_30 word19_30 R_wl
Cwl_20_30 word20_30 gnd C_wl
Rw21_30 word21_30 word20_30 R_wl
Cwl_21_30 word21_30 gnd C_wl
Rw22_30 word22_30 word21_30 R_wl
Cwl_22_30 word22_30 gnd C_wl
Rw23_30 word23_30 word22_30 R_wl
Cwl_23_30 word23_30 gnd C_wl
Rw24_30 word24_30 word23_30 R_wl
Cwl_24_30 word24_30 gnd C_wl
Rw25_30 word25_30 word24_30 R_wl
Cwl_25_30 word25_30 gnd C_wl
Rw26_30 word26_30 word25_30 R_wl
Cwl_26_30 word26_30 gnd C_wl
Rw27_30 word27_30 word26_30 R_wl
Cwl_27_30 word27_30 gnd C_wl
Rw28_30 word28_30 word27_30 R_wl
Cwl_28_30 word28_30 gnd C_wl
Rw29_30 word29_30 word28_30 R_wl
Cwl_29_30 word29_30 gnd C_wl
Rw30_30 word30_30 word29_30 R_wl
Cwl_30_30 word30_30 gnd C_wl
Rw31_30 word31_30 word30_30 R_wl
Cwl_31_30 word31_30 gnd C_wl
Rw32_30 word32_30 word31_30 R_wl
Cwl_32_30 word32_30 gnd C_wl
Rw33_30 word33_30 word32_30 R_wl
Cwl_33_30 word33_30 gnd C_wl
Rw34_30 word34_30 word33_30 R_wl
Cwl_34_30 word34_30 gnd C_wl
Rw35_30 word35_30 word34_30 R_wl
Cwl_35_30 word35_30 gnd C_wl
Rw36_30 word36_30 word35_30 R_wl
Cwl_36_30 word36_30 gnd C_wl
Rw37_30 word37_30 word36_30 R_wl
Cwl_37_30 word37_30 gnd C_wl
Rw38_30 word38_30 word37_30 R_wl
Cwl_38_30 word38_30 gnd C_wl
Rw39_30 word39_30 word38_30 R_wl
Cwl_39_30 word39_30 gnd C_wl
Rw40_30 word40_30 word39_30 R_wl
Cwl_40_30 word40_30 gnd C_wl
Rw41_30 word41_30 word40_30 R_wl
Cwl_41_30 word41_30 gnd C_wl
Rw42_30 word42_30 word41_30 R_wl
Cwl_42_30 word42_30 gnd C_wl
Rw43_30 word43_30 word42_30 R_wl
Cwl_43_30 word43_30 gnd C_wl
Rw44_30 word44_30 word43_30 R_wl
Cwl_44_30 word44_30 gnd C_wl
Rw45_30 word45_30 word44_30 R_wl
Cwl_45_30 word45_30 gnd C_wl
Rw46_30 word46_30 word45_30 R_wl
Cwl_46_30 word46_30 gnd C_wl
Rw47_30 word47_30 word46_30 R_wl
Cwl_47_30 word47_30 gnd C_wl
Rw48_30 word48_30 word47_30 R_wl
Cwl_48_30 word48_30 gnd C_wl
Rw49_30 word49_30 word48_30 R_wl
Cwl_49_30 word49_30 gnd C_wl
Rw50_30 word50_30 word49_30 R_wl
Cwl_50_30 word50_30 gnd C_wl
Rw51_30 word51_30 word50_30 R_wl
Cwl_51_30 word51_30 gnd C_wl
Rw52_30 word52_30 word51_30 R_wl
Cwl_52_30 word52_30 gnd C_wl
Rw53_30 word53_30 word52_30 R_wl
Cwl_53_30 word53_30 gnd C_wl
Rw54_30 word54_30 word53_30 R_wl
Cwl_54_30 word54_30 gnd C_wl
Rw55_30 word55_30 word54_30 R_wl
Cwl_55_30 word55_30 gnd C_wl
Rw56_30 word56_30 word55_30 R_wl
Cwl_56_30 word56_30 gnd C_wl
Rw57_30 word57_30 word56_30 R_wl
Cwl_57_30 word57_30 gnd C_wl
Rw58_30 word58_30 word57_30 R_wl
Cwl_58_30 word58_30 gnd C_wl
Rw59_30 word59_30 word58_30 R_wl
Cwl_59_30 word59_30 gnd C_wl
Rw60_30 word60_30 word59_30 R_wl
Cwl_60_30 word60_30 gnd C_wl
Rw61_30 word61_30 word60_30 R_wl
Cwl_61_30 word61_30 gnd C_wl
Rw62_30 word62_30 word61_30 R_wl
Cwl_62_30 word62_30 gnd C_wl
Rw63_30 word63_30 word62_30 R_wl
Cwl_63_30 word63_30 gnd C_wl
Rw64_30 word64_30 word63_30 R_wl
Cwl_64_30 word64_30 gnd C_wl
Rw65_30 word65_30 word64_30 R_wl
Cwl_65_30 word65_30 gnd C_wl
Rw66_30 word66_30 word65_30 R_wl
Cwl_66_30 word66_30 gnd C_wl
Rw67_30 word67_30 word66_30 R_wl
Cwl_67_30 word67_30 gnd C_wl
Rw68_30 word68_30 word67_30 R_wl
Cwl_68_30 word68_30 gnd C_wl
Rw69_30 word69_30 word68_30 R_wl
Cwl_69_30 word69_30 gnd C_wl
Rw70_30 word70_30 word69_30 R_wl
Cwl_70_30 word70_30 gnd C_wl
Rw71_30 word71_30 word70_30 R_wl
Cwl_71_30 word71_30 gnd C_wl
Rw72_30 word72_30 word71_30 R_wl
Cwl_72_30 word72_30 gnd C_wl
Rw73_30 word73_30 word72_30 R_wl
Cwl_73_30 word73_30 gnd C_wl
Rw74_30 word74_30 word73_30 R_wl
Cwl_74_30 word74_30 gnd C_wl
Rw75_30 word75_30 word74_30 R_wl
Cwl_75_30 word75_30 gnd C_wl
Rw76_30 word76_30 word75_30 R_wl
Cwl_76_30 word76_30 gnd C_wl
Rw77_30 word77_30 word76_30 R_wl
Cwl_77_30 word77_30 gnd C_wl
Rw78_30 word78_30 word77_30 R_wl
Cwl_78_30 word78_30 gnd C_wl
Rw79_30 word79_30 word78_30 R_wl
Cwl_79_30 word79_30 gnd C_wl
Rw80_30 word80_30 word79_30 R_wl
Cwl_80_30 word80_30 gnd C_wl
Rw81_30 word81_30 word80_30 R_wl
Cwl_81_30 word81_30 gnd C_wl
Rw82_30 word82_30 word81_30 R_wl
Cwl_82_30 word82_30 gnd C_wl
Rw83_30 word83_30 word82_30 R_wl
Cwl_83_30 word83_30 gnd C_wl
Rw84_30 word84_30 word83_30 R_wl
Cwl_84_30 word84_30 gnd C_wl
Rw85_30 word85_30 word84_30 R_wl
Cwl_85_30 word85_30 gnd C_wl
Rw86_30 word86_30 word85_30 R_wl
Cwl_86_30 word86_30 gnd C_wl
Rw87_30 word87_30 word86_30 R_wl
Cwl_87_30 word87_30 gnd C_wl
Rw88_30 word88_30 word87_30 R_wl
Cwl_88_30 word88_30 gnd C_wl
Rw89_30 word89_30 word88_30 R_wl
Cwl_89_30 word89_30 gnd C_wl
Rw90_30 word90_30 word89_30 R_wl
Cwl_90_30 word90_30 gnd C_wl
Rw91_30 word91_30 word90_30 R_wl
Cwl_91_30 word91_30 gnd C_wl
Rw92_30 word92_30 word91_30 R_wl
Cwl_92_30 word92_30 gnd C_wl
Rw93_30 word93_30 word92_30 R_wl
Cwl_93_30 word93_30 gnd C_wl
Rw94_30 word94_30 word93_30 R_wl
Cwl_94_30 word94_30 gnd C_wl
Rw95_30 word95_30 word94_30 R_wl
Cwl_95_30 word95_30 gnd C_wl
Rw96_30 word96_30 word95_30 R_wl
Cwl_96_30 word96_30 gnd C_wl
Rw97_30 word97_30 word96_30 R_wl
Cwl_97_30 word97_30 gnd C_wl
Rw98_30 word98_30 word97_30 R_wl
Cwl_98_30 word98_30 gnd C_wl
Rw99_30 word99_30 word98_30 R_wl
Cwl_99_30 word99_30 gnd C_wl
Vwl_31 word_31 0 0
Rw0_31 word_31 word0_31 R_wl
Cwl_0_31 word0_31 gnd C_wl
Rw1_31 word1_31 word0_31 R_wl
Cwl_1_31 word1_31 gnd C_wl
Rw2_31 word2_31 word1_31 R_wl
Cwl_2_31 word2_31 gnd C_wl
Rw3_31 word3_31 word2_31 R_wl
Cwl_3_31 word3_31 gnd C_wl
Rw4_31 word4_31 word3_31 R_wl
Cwl_4_31 word4_31 gnd C_wl
Rw5_31 word5_31 word4_31 R_wl
Cwl_5_31 word5_31 gnd C_wl
Rw6_31 word6_31 word5_31 R_wl
Cwl_6_31 word6_31 gnd C_wl
Rw7_31 word7_31 word6_31 R_wl
Cwl_7_31 word7_31 gnd C_wl
Rw8_31 word8_31 word7_31 R_wl
Cwl_8_31 word8_31 gnd C_wl
Rw9_31 word9_31 word8_31 R_wl
Cwl_9_31 word9_31 gnd C_wl
Rw10_31 word10_31 word9_31 R_wl
Cwl_10_31 word10_31 gnd C_wl
Rw11_31 word11_31 word10_31 R_wl
Cwl_11_31 word11_31 gnd C_wl
Rw12_31 word12_31 word11_31 R_wl
Cwl_12_31 word12_31 gnd C_wl
Rw13_31 word13_31 word12_31 R_wl
Cwl_13_31 word13_31 gnd C_wl
Rw14_31 word14_31 word13_31 R_wl
Cwl_14_31 word14_31 gnd C_wl
Rw15_31 word15_31 word14_31 R_wl
Cwl_15_31 word15_31 gnd C_wl
Rw16_31 word16_31 word15_31 R_wl
Cwl_16_31 word16_31 gnd C_wl
Rw17_31 word17_31 word16_31 R_wl
Cwl_17_31 word17_31 gnd C_wl
Rw18_31 word18_31 word17_31 R_wl
Cwl_18_31 word18_31 gnd C_wl
Rw19_31 word19_31 word18_31 R_wl
Cwl_19_31 word19_31 gnd C_wl
Rw20_31 word20_31 word19_31 R_wl
Cwl_20_31 word20_31 gnd C_wl
Rw21_31 word21_31 word20_31 R_wl
Cwl_21_31 word21_31 gnd C_wl
Rw22_31 word22_31 word21_31 R_wl
Cwl_22_31 word22_31 gnd C_wl
Rw23_31 word23_31 word22_31 R_wl
Cwl_23_31 word23_31 gnd C_wl
Rw24_31 word24_31 word23_31 R_wl
Cwl_24_31 word24_31 gnd C_wl
Rw25_31 word25_31 word24_31 R_wl
Cwl_25_31 word25_31 gnd C_wl
Rw26_31 word26_31 word25_31 R_wl
Cwl_26_31 word26_31 gnd C_wl
Rw27_31 word27_31 word26_31 R_wl
Cwl_27_31 word27_31 gnd C_wl
Rw28_31 word28_31 word27_31 R_wl
Cwl_28_31 word28_31 gnd C_wl
Rw29_31 word29_31 word28_31 R_wl
Cwl_29_31 word29_31 gnd C_wl
Rw30_31 word30_31 word29_31 R_wl
Cwl_30_31 word30_31 gnd C_wl
Rw31_31 word31_31 word30_31 R_wl
Cwl_31_31 word31_31 gnd C_wl
Rw32_31 word32_31 word31_31 R_wl
Cwl_32_31 word32_31 gnd C_wl
Rw33_31 word33_31 word32_31 R_wl
Cwl_33_31 word33_31 gnd C_wl
Rw34_31 word34_31 word33_31 R_wl
Cwl_34_31 word34_31 gnd C_wl
Rw35_31 word35_31 word34_31 R_wl
Cwl_35_31 word35_31 gnd C_wl
Rw36_31 word36_31 word35_31 R_wl
Cwl_36_31 word36_31 gnd C_wl
Rw37_31 word37_31 word36_31 R_wl
Cwl_37_31 word37_31 gnd C_wl
Rw38_31 word38_31 word37_31 R_wl
Cwl_38_31 word38_31 gnd C_wl
Rw39_31 word39_31 word38_31 R_wl
Cwl_39_31 word39_31 gnd C_wl
Rw40_31 word40_31 word39_31 R_wl
Cwl_40_31 word40_31 gnd C_wl
Rw41_31 word41_31 word40_31 R_wl
Cwl_41_31 word41_31 gnd C_wl
Rw42_31 word42_31 word41_31 R_wl
Cwl_42_31 word42_31 gnd C_wl
Rw43_31 word43_31 word42_31 R_wl
Cwl_43_31 word43_31 gnd C_wl
Rw44_31 word44_31 word43_31 R_wl
Cwl_44_31 word44_31 gnd C_wl
Rw45_31 word45_31 word44_31 R_wl
Cwl_45_31 word45_31 gnd C_wl
Rw46_31 word46_31 word45_31 R_wl
Cwl_46_31 word46_31 gnd C_wl
Rw47_31 word47_31 word46_31 R_wl
Cwl_47_31 word47_31 gnd C_wl
Rw48_31 word48_31 word47_31 R_wl
Cwl_48_31 word48_31 gnd C_wl
Rw49_31 word49_31 word48_31 R_wl
Cwl_49_31 word49_31 gnd C_wl
Rw50_31 word50_31 word49_31 R_wl
Cwl_50_31 word50_31 gnd C_wl
Rw51_31 word51_31 word50_31 R_wl
Cwl_51_31 word51_31 gnd C_wl
Rw52_31 word52_31 word51_31 R_wl
Cwl_52_31 word52_31 gnd C_wl
Rw53_31 word53_31 word52_31 R_wl
Cwl_53_31 word53_31 gnd C_wl
Rw54_31 word54_31 word53_31 R_wl
Cwl_54_31 word54_31 gnd C_wl
Rw55_31 word55_31 word54_31 R_wl
Cwl_55_31 word55_31 gnd C_wl
Rw56_31 word56_31 word55_31 R_wl
Cwl_56_31 word56_31 gnd C_wl
Rw57_31 word57_31 word56_31 R_wl
Cwl_57_31 word57_31 gnd C_wl
Rw58_31 word58_31 word57_31 R_wl
Cwl_58_31 word58_31 gnd C_wl
Rw59_31 word59_31 word58_31 R_wl
Cwl_59_31 word59_31 gnd C_wl
Rw60_31 word60_31 word59_31 R_wl
Cwl_60_31 word60_31 gnd C_wl
Rw61_31 word61_31 word60_31 R_wl
Cwl_61_31 word61_31 gnd C_wl
Rw62_31 word62_31 word61_31 R_wl
Cwl_62_31 word62_31 gnd C_wl
Rw63_31 word63_31 word62_31 R_wl
Cwl_63_31 word63_31 gnd C_wl
Rw64_31 word64_31 word63_31 R_wl
Cwl_64_31 word64_31 gnd C_wl
Rw65_31 word65_31 word64_31 R_wl
Cwl_65_31 word65_31 gnd C_wl
Rw66_31 word66_31 word65_31 R_wl
Cwl_66_31 word66_31 gnd C_wl
Rw67_31 word67_31 word66_31 R_wl
Cwl_67_31 word67_31 gnd C_wl
Rw68_31 word68_31 word67_31 R_wl
Cwl_68_31 word68_31 gnd C_wl
Rw69_31 word69_31 word68_31 R_wl
Cwl_69_31 word69_31 gnd C_wl
Rw70_31 word70_31 word69_31 R_wl
Cwl_70_31 word70_31 gnd C_wl
Rw71_31 word71_31 word70_31 R_wl
Cwl_71_31 word71_31 gnd C_wl
Rw72_31 word72_31 word71_31 R_wl
Cwl_72_31 word72_31 gnd C_wl
Rw73_31 word73_31 word72_31 R_wl
Cwl_73_31 word73_31 gnd C_wl
Rw74_31 word74_31 word73_31 R_wl
Cwl_74_31 word74_31 gnd C_wl
Rw75_31 word75_31 word74_31 R_wl
Cwl_75_31 word75_31 gnd C_wl
Rw76_31 word76_31 word75_31 R_wl
Cwl_76_31 word76_31 gnd C_wl
Rw77_31 word77_31 word76_31 R_wl
Cwl_77_31 word77_31 gnd C_wl
Rw78_31 word78_31 word77_31 R_wl
Cwl_78_31 word78_31 gnd C_wl
Rw79_31 word79_31 word78_31 R_wl
Cwl_79_31 word79_31 gnd C_wl
Rw80_31 word80_31 word79_31 R_wl
Cwl_80_31 word80_31 gnd C_wl
Rw81_31 word81_31 word80_31 R_wl
Cwl_81_31 word81_31 gnd C_wl
Rw82_31 word82_31 word81_31 R_wl
Cwl_82_31 word82_31 gnd C_wl
Rw83_31 word83_31 word82_31 R_wl
Cwl_83_31 word83_31 gnd C_wl
Rw84_31 word84_31 word83_31 R_wl
Cwl_84_31 word84_31 gnd C_wl
Rw85_31 word85_31 word84_31 R_wl
Cwl_85_31 word85_31 gnd C_wl
Rw86_31 word86_31 word85_31 R_wl
Cwl_86_31 word86_31 gnd C_wl
Rw87_31 word87_31 word86_31 R_wl
Cwl_87_31 word87_31 gnd C_wl
Rw88_31 word88_31 word87_31 R_wl
Cwl_88_31 word88_31 gnd C_wl
Rw89_31 word89_31 word88_31 R_wl
Cwl_89_31 word89_31 gnd C_wl
Rw90_31 word90_31 word89_31 R_wl
Cwl_90_31 word90_31 gnd C_wl
Rw91_31 word91_31 word90_31 R_wl
Cwl_91_31 word91_31 gnd C_wl
Rw92_31 word92_31 word91_31 R_wl
Cwl_92_31 word92_31 gnd C_wl
Rw93_31 word93_31 word92_31 R_wl
Cwl_93_31 word93_31 gnd C_wl
Rw94_31 word94_31 word93_31 R_wl
Cwl_94_31 word94_31 gnd C_wl
Rw95_31 word95_31 word94_31 R_wl
Cwl_95_31 word95_31 gnd C_wl
Rw96_31 word96_31 word95_31 R_wl
Cwl_96_31 word96_31 gnd C_wl
Rw97_31 word97_31 word96_31 R_wl
Cwl_97_31 word97_31 gnd C_wl
Rw98_31 word98_31 word97_31 R_wl
Cwl_98_31 word98_31 gnd C_wl
Rw99_31 word99_31 word98_31 R_wl
Cwl_99_31 word99_31 gnd C_wl
Vwl_32 word_32 0 0
Rw0_32 word_32 word0_32 R_wl
Cwl_0_32 word0_32 gnd C_wl
Rw1_32 word1_32 word0_32 R_wl
Cwl_1_32 word1_32 gnd C_wl
Rw2_32 word2_32 word1_32 R_wl
Cwl_2_32 word2_32 gnd C_wl
Rw3_32 word3_32 word2_32 R_wl
Cwl_3_32 word3_32 gnd C_wl
Rw4_32 word4_32 word3_32 R_wl
Cwl_4_32 word4_32 gnd C_wl
Rw5_32 word5_32 word4_32 R_wl
Cwl_5_32 word5_32 gnd C_wl
Rw6_32 word6_32 word5_32 R_wl
Cwl_6_32 word6_32 gnd C_wl
Rw7_32 word7_32 word6_32 R_wl
Cwl_7_32 word7_32 gnd C_wl
Rw8_32 word8_32 word7_32 R_wl
Cwl_8_32 word8_32 gnd C_wl
Rw9_32 word9_32 word8_32 R_wl
Cwl_9_32 word9_32 gnd C_wl
Rw10_32 word10_32 word9_32 R_wl
Cwl_10_32 word10_32 gnd C_wl
Rw11_32 word11_32 word10_32 R_wl
Cwl_11_32 word11_32 gnd C_wl
Rw12_32 word12_32 word11_32 R_wl
Cwl_12_32 word12_32 gnd C_wl
Rw13_32 word13_32 word12_32 R_wl
Cwl_13_32 word13_32 gnd C_wl
Rw14_32 word14_32 word13_32 R_wl
Cwl_14_32 word14_32 gnd C_wl
Rw15_32 word15_32 word14_32 R_wl
Cwl_15_32 word15_32 gnd C_wl
Rw16_32 word16_32 word15_32 R_wl
Cwl_16_32 word16_32 gnd C_wl
Rw17_32 word17_32 word16_32 R_wl
Cwl_17_32 word17_32 gnd C_wl
Rw18_32 word18_32 word17_32 R_wl
Cwl_18_32 word18_32 gnd C_wl
Rw19_32 word19_32 word18_32 R_wl
Cwl_19_32 word19_32 gnd C_wl
Rw20_32 word20_32 word19_32 R_wl
Cwl_20_32 word20_32 gnd C_wl
Rw21_32 word21_32 word20_32 R_wl
Cwl_21_32 word21_32 gnd C_wl
Rw22_32 word22_32 word21_32 R_wl
Cwl_22_32 word22_32 gnd C_wl
Rw23_32 word23_32 word22_32 R_wl
Cwl_23_32 word23_32 gnd C_wl
Rw24_32 word24_32 word23_32 R_wl
Cwl_24_32 word24_32 gnd C_wl
Rw25_32 word25_32 word24_32 R_wl
Cwl_25_32 word25_32 gnd C_wl
Rw26_32 word26_32 word25_32 R_wl
Cwl_26_32 word26_32 gnd C_wl
Rw27_32 word27_32 word26_32 R_wl
Cwl_27_32 word27_32 gnd C_wl
Rw28_32 word28_32 word27_32 R_wl
Cwl_28_32 word28_32 gnd C_wl
Rw29_32 word29_32 word28_32 R_wl
Cwl_29_32 word29_32 gnd C_wl
Rw30_32 word30_32 word29_32 R_wl
Cwl_30_32 word30_32 gnd C_wl
Rw31_32 word31_32 word30_32 R_wl
Cwl_31_32 word31_32 gnd C_wl
Rw32_32 word32_32 word31_32 R_wl
Cwl_32_32 word32_32 gnd C_wl
Rw33_32 word33_32 word32_32 R_wl
Cwl_33_32 word33_32 gnd C_wl
Rw34_32 word34_32 word33_32 R_wl
Cwl_34_32 word34_32 gnd C_wl
Rw35_32 word35_32 word34_32 R_wl
Cwl_35_32 word35_32 gnd C_wl
Rw36_32 word36_32 word35_32 R_wl
Cwl_36_32 word36_32 gnd C_wl
Rw37_32 word37_32 word36_32 R_wl
Cwl_37_32 word37_32 gnd C_wl
Rw38_32 word38_32 word37_32 R_wl
Cwl_38_32 word38_32 gnd C_wl
Rw39_32 word39_32 word38_32 R_wl
Cwl_39_32 word39_32 gnd C_wl
Rw40_32 word40_32 word39_32 R_wl
Cwl_40_32 word40_32 gnd C_wl
Rw41_32 word41_32 word40_32 R_wl
Cwl_41_32 word41_32 gnd C_wl
Rw42_32 word42_32 word41_32 R_wl
Cwl_42_32 word42_32 gnd C_wl
Rw43_32 word43_32 word42_32 R_wl
Cwl_43_32 word43_32 gnd C_wl
Rw44_32 word44_32 word43_32 R_wl
Cwl_44_32 word44_32 gnd C_wl
Rw45_32 word45_32 word44_32 R_wl
Cwl_45_32 word45_32 gnd C_wl
Rw46_32 word46_32 word45_32 R_wl
Cwl_46_32 word46_32 gnd C_wl
Rw47_32 word47_32 word46_32 R_wl
Cwl_47_32 word47_32 gnd C_wl
Rw48_32 word48_32 word47_32 R_wl
Cwl_48_32 word48_32 gnd C_wl
Rw49_32 word49_32 word48_32 R_wl
Cwl_49_32 word49_32 gnd C_wl
Rw50_32 word50_32 word49_32 R_wl
Cwl_50_32 word50_32 gnd C_wl
Rw51_32 word51_32 word50_32 R_wl
Cwl_51_32 word51_32 gnd C_wl
Rw52_32 word52_32 word51_32 R_wl
Cwl_52_32 word52_32 gnd C_wl
Rw53_32 word53_32 word52_32 R_wl
Cwl_53_32 word53_32 gnd C_wl
Rw54_32 word54_32 word53_32 R_wl
Cwl_54_32 word54_32 gnd C_wl
Rw55_32 word55_32 word54_32 R_wl
Cwl_55_32 word55_32 gnd C_wl
Rw56_32 word56_32 word55_32 R_wl
Cwl_56_32 word56_32 gnd C_wl
Rw57_32 word57_32 word56_32 R_wl
Cwl_57_32 word57_32 gnd C_wl
Rw58_32 word58_32 word57_32 R_wl
Cwl_58_32 word58_32 gnd C_wl
Rw59_32 word59_32 word58_32 R_wl
Cwl_59_32 word59_32 gnd C_wl
Rw60_32 word60_32 word59_32 R_wl
Cwl_60_32 word60_32 gnd C_wl
Rw61_32 word61_32 word60_32 R_wl
Cwl_61_32 word61_32 gnd C_wl
Rw62_32 word62_32 word61_32 R_wl
Cwl_62_32 word62_32 gnd C_wl
Rw63_32 word63_32 word62_32 R_wl
Cwl_63_32 word63_32 gnd C_wl
Rw64_32 word64_32 word63_32 R_wl
Cwl_64_32 word64_32 gnd C_wl
Rw65_32 word65_32 word64_32 R_wl
Cwl_65_32 word65_32 gnd C_wl
Rw66_32 word66_32 word65_32 R_wl
Cwl_66_32 word66_32 gnd C_wl
Rw67_32 word67_32 word66_32 R_wl
Cwl_67_32 word67_32 gnd C_wl
Rw68_32 word68_32 word67_32 R_wl
Cwl_68_32 word68_32 gnd C_wl
Rw69_32 word69_32 word68_32 R_wl
Cwl_69_32 word69_32 gnd C_wl
Rw70_32 word70_32 word69_32 R_wl
Cwl_70_32 word70_32 gnd C_wl
Rw71_32 word71_32 word70_32 R_wl
Cwl_71_32 word71_32 gnd C_wl
Rw72_32 word72_32 word71_32 R_wl
Cwl_72_32 word72_32 gnd C_wl
Rw73_32 word73_32 word72_32 R_wl
Cwl_73_32 word73_32 gnd C_wl
Rw74_32 word74_32 word73_32 R_wl
Cwl_74_32 word74_32 gnd C_wl
Rw75_32 word75_32 word74_32 R_wl
Cwl_75_32 word75_32 gnd C_wl
Rw76_32 word76_32 word75_32 R_wl
Cwl_76_32 word76_32 gnd C_wl
Rw77_32 word77_32 word76_32 R_wl
Cwl_77_32 word77_32 gnd C_wl
Rw78_32 word78_32 word77_32 R_wl
Cwl_78_32 word78_32 gnd C_wl
Rw79_32 word79_32 word78_32 R_wl
Cwl_79_32 word79_32 gnd C_wl
Rw80_32 word80_32 word79_32 R_wl
Cwl_80_32 word80_32 gnd C_wl
Rw81_32 word81_32 word80_32 R_wl
Cwl_81_32 word81_32 gnd C_wl
Rw82_32 word82_32 word81_32 R_wl
Cwl_82_32 word82_32 gnd C_wl
Rw83_32 word83_32 word82_32 R_wl
Cwl_83_32 word83_32 gnd C_wl
Rw84_32 word84_32 word83_32 R_wl
Cwl_84_32 word84_32 gnd C_wl
Rw85_32 word85_32 word84_32 R_wl
Cwl_85_32 word85_32 gnd C_wl
Rw86_32 word86_32 word85_32 R_wl
Cwl_86_32 word86_32 gnd C_wl
Rw87_32 word87_32 word86_32 R_wl
Cwl_87_32 word87_32 gnd C_wl
Rw88_32 word88_32 word87_32 R_wl
Cwl_88_32 word88_32 gnd C_wl
Rw89_32 word89_32 word88_32 R_wl
Cwl_89_32 word89_32 gnd C_wl
Rw90_32 word90_32 word89_32 R_wl
Cwl_90_32 word90_32 gnd C_wl
Rw91_32 word91_32 word90_32 R_wl
Cwl_91_32 word91_32 gnd C_wl
Rw92_32 word92_32 word91_32 R_wl
Cwl_92_32 word92_32 gnd C_wl
Rw93_32 word93_32 word92_32 R_wl
Cwl_93_32 word93_32 gnd C_wl
Rw94_32 word94_32 word93_32 R_wl
Cwl_94_32 word94_32 gnd C_wl
Rw95_32 word95_32 word94_32 R_wl
Cwl_95_32 word95_32 gnd C_wl
Rw96_32 word96_32 word95_32 R_wl
Cwl_96_32 word96_32 gnd C_wl
Rw97_32 word97_32 word96_32 R_wl
Cwl_97_32 word97_32 gnd C_wl
Rw98_32 word98_32 word97_32 R_wl
Cwl_98_32 word98_32 gnd C_wl
Rw99_32 word99_32 word98_32 R_wl
Cwl_99_32 word99_32 gnd C_wl
Vwl_33 word_33 0 0
Rw0_33 word_33 word0_33 R_wl
Cwl_0_33 word0_33 gnd C_wl
Rw1_33 word1_33 word0_33 R_wl
Cwl_1_33 word1_33 gnd C_wl
Rw2_33 word2_33 word1_33 R_wl
Cwl_2_33 word2_33 gnd C_wl
Rw3_33 word3_33 word2_33 R_wl
Cwl_3_33 word3_33 gnd C_wl
Rw4_33 word4_33 word3_33 R_wl
Cwl_4_33 word4_33 gnd C_wl
Rw5_33 word5_33 word4_33 R_wl
Cwl_5_33 word5_33 gnd C_wl
Rw6_33 word6_33 word5_33 R_wl
Cwl_6_33 word6_33 gnd C_wl
Rw7_33 word7_33 word6_33 R_wl
Cwl_7_33 word7_33 gnd C_wl
Rw8_33 word8_33 word7_33 R_wl
Cwl_8_33 word8_33 gnd C_wl
Rw9_33 word9_33 word8_33 R_wl
Cwl_9_33 word9_33 gnd C_wl
Rw10_33 word10_33 word9_33 R_wl
Cwl_10_33 word10_33 gnd C_wl
Rw11_33 word11_33 word10_33 R_wl
Cwl_11_33 word11_33 gnd C_wl
Rw12_33 word12_33 word11_33 R_wl
Cwl_12_33 word12_33 gnd C_wl
Rw13_33 word13_33 word12_33 R_wl
Cwl_13_33 word13_33 gnd C_wl
Rw14_33 word14_33 word13_33 R_wl
Cwl_14_33 word14_33 gnd C_wl
Rw15_33 word15_33 word14_33 R_wl
Cwl_15_33 word15_33 gnd C_wl
Rw16_33 word16_33 word15_33 R_wl
Cwl_16_33 word16_33 gnd C_wl
Rw17_33 word17_33 word16_33 R_wl
Cwl_17_33 word17_33 gnd C_wl
Rw18_33 word18_33 word17_33 R_wl
Cwl_18_33 word18_33 gnd C_wl
Rw19_33 word19_33 word18_33 R_wl
Cwl_19_33 word19_33 gnd C_wl
Rw20_33 word20_33 word19_33 R_wl
Cwl_20_33 word20_33 gnd C_wl
Rw21_33 word21_33 word20_33 R_wl
Cwl_21_33 word21_33 gnd C_wl
Rw22_33 word22_33 word21_33 R_wl
Cwl_22_33 word22_33 gnd C_wl
Rw23_33 word23_33 word22_33 R_wl
Cwl_23_33 word23_33 gnd C_wl
Rw24_33 word24_33 word23_33 R_wl
Cwl_24_33 word24_33 gnd C_wl
Rw25_33 word25_33 word24_33 R_wl
Cwl_25_33 word25_33 gnd C_wl
Rw26_33 word26_33 word25_33 R_wl
Cwl_26_33 word26_33 gnd C_wl
Rw27_33 word27_33 word26_33 R_wl
Cwl_27_33 word27_33 gnd C_wl
Rw28_33 word28_33 word27_33 R_wl
Cwl_28_33 word28_33 gnd C_wl
Rw29_33 word29_33 word28_33 R_wl
Cwl_29_33 word29_33 gnd C_wl
Rw30_33 word30_33 word29_33 R_wl
Cwl_30_33 word30_33 gnd C_wl
Rw31_33 word31_33 word30_33 R_wl
Cwl_31_33 word31_33 gnd C_wl
Rw32_33 word32_33 word31_33 R_wl
Cwl_32_33 word32_33 gnd C_wl
Rw33_33 word33_33 word32_33 R_wl
Cwl_33_33 word33_33 gnd C_wl
Rw34_33 word34_33 word33_33 R_wl
Cwl_34_33 word34_33 gnd C_wl
Rw35_33 word35_33 word34_33 R_wl
Cwl_35_33 word35_33 gnd C_wl
Rw36_33 word36_33 word35_33 R_wl
Cwl_36_33 word36_33 gnd C_wl
Rw37_33 word37_33 word36_33 R_wl
Cwl_37_33 word37_33 gnd C_wl
Rw38_33 word38_33 word37_33 R_wl
Cwl_38_33 word38_33 gnd C_wl
Rw39_33 word39_33 word38_33 R_wl
Cwl_39_33 word39_33 gnd C_wl
Rw40_33 word40_33 word39_33 R_wl
Cwl_40_33 word40_33 gnd C_wl
Rw41_33 word41_33 word40_33 R_wl
Cwl_41_33 word41_33 gnd C_wl
Rw42_33 word42_33 word41_33 R_wl
Cwl_42_33 word42_33 gnd C_wl
Rw43_33 word43_33 word42_33 R_wl
Cwl_43_33 word43_33 gnd C_wl
Rw44_33 word44_33 word43_33 R_wl
Cwl_44_33 word44_33 gnd C_wl
Rw45_33 word45_33 word44_33 R_wl
Cwl_45_33 word45_33 gnd C_wl
Rw46_33 word46_33 word45_33 R_wl
Cwl_46_33 word46_33 gnd C_wl
Rw47_33 word47_33 word46_33 R_wl
Cwl_47_33 word47_33 gnd C_wl
Rw48_33 word48_33 word47_33 R_wl
Cwl_48_33 word48_33 gnd C_wl
Rw49_33 word49_33 word48_33 R_wl
Cwl_49_33 word49_33 gnd C_wl
Rw50_33 word50_33 word49_33 R_wl
Cwl_50_33 word50_33 gnd C_wl
Rw51_33 word51_33 word50_33 R_wl
Cwl_51_33 word51_33 gnd C_wl
Rw52_33 word52_33 word51_33 R_wl
Cwl_52_33 word52_33 gnd C_wl
Rw53_33 word53_33 word52_33 R_wl
Cwl_53_33 word53_33 gnd C_wl
Rw54_33 word54_33 word53_33 R_wl
Cwl_54_33 word54_33 gnd C_wl
Rw55_33 word55_33 word54_33 R_wl
Cwl_55_33 word55_33 gnd C_wl
Rw56_33 word56_33 word55_33 R_wl
Cwl_56_33 word56_33 gnd C_wl
Rw57_33 word57_33 word56_33 R_wl
Cwl_57_33 word57_33 gnd C_wl
Rw58_33 word58_33 word57_33 R_wl
Cwl_58_33 word58_33 gnd C_wl
Rw59_33 word59_33 word58_33 R_wl
Cwl_59_33 word59_33 gnd C_wl
Rw60_33 word60_33 word59_33 R_wl
Cwl_60_33 word60_33 gnd C_wl
Rw61_33 word61_33 word60_33 R_wl
Cwl_61_33 word61_33 gnd C_wl
Rw62_33 word62_33 word61_33 R_wl
Cwl_62_33 word62_33 gnd C_wl
Rw63_33 word63_33 word62_33 R_wl
Cwl_63_33 word63_33 gnd C_wl
Rw64_33 word64_33 word63_33 R_wl
Cwl_64_33 word64_33 gnd C_wl
Rw65_33 word65_33 word64_33 R_wl
Cwl_65_33 word65_33 gnd C_wl
Rw66_33 word66_33 word65_33 R_wl
Cwl_66_33 word66_33 gnd C_wl
Rw67_33 word67_33 word66_33 R_wl
Cwl_67_33 word67_33 gnd C_wl
Rw68_33 word68_33 word67_33 R_wl
Cwl_68_33 word68_33 gnd C_wl
Rw69_33 word69_33 word68_33 R_wl
Cwl_69_33 word69_33 gnd C_wl
Rw70_33 word70_33 word69_33 R_wl
Cwl_70_33 word70_33 gnd C_wl
Rw71_33 word71_33 word70_33 R_wl
Cwl_71_33 word71_33 gnd C_wl
Rw72_33 word72_33 word71_33 R_wl
Cwl_72_33 word72_33 gnd C_wl
Rw73_33 word73_33 word72_33 R_wl
Cwl_73_33 word73_33 gnd C_wl
Rw74_33 word74_33 word73_33 R_wl
Cwl_74_33 word74_33 gnd C_wl
Rw75_33 word75_33 word74_33 R_wl
Cwl_75_33 word75_33 gnd C_wl
Rw76_33 word76_33 word75_33 R_wl
Cwl_76_33 word76_33 gnd C_wl
Rw77_33 word77_33 word76_33 R_wl
Cwl_77_33 word77_33 gnd C_wl
Rw78_33 word78_33 word77_33 R_wl
Cwl_78_33 word78_33 gnd C_wl
Rw79_33 word79_33 word78_33 R_wl
Cwl_79_33 word79_33 gnd C_wl
Rw80_33 word80_33 word79_33 R_wl
Cwl_80_33 word80_33 gnd C_wl
Rw81_33 word81_33 word80_33 R_wl
Cwl_81_33 word81_33 gnd C_wl
Rw82_33 word82_33 word81_33 R_wl
Cwl_82_33 word82_33 gnd C_wl
Rw83_33 word83_33 word82_33 R_wl
Cwl_83_33 word83_33 gnd C_wl
Rw84_33 word84_33 word83_33 R_wl
Cwl_84_33 word84_33 gnd C_wl
Rw85_33 word85_33 word84_33 R_wl
Cwl_85_33 word85_33 gnd C_wl
Rw86_33 word86_33 word85_33 R_wl
Cwl_86_33 word86_33 gnd C_wl
Rw87_33 word87_33 word86_33 R_wl
Cwl_87_33 word87_33 gnd C_wl
Rw88_33 word88_33 word87_33 R_wl
Cwl_88_33 word88_33 gnd C_wl
Rw89_33 word89_33 word88_33 R_wl
Cwl_89_33 word89_33 gnd C_wl
Rw90_33 word90_33 word89_33 R_wl
Cwl_90_33 word90_33 gnd C_wl
Rw91_33 word91_33 word90_33 R_wl
Cwl_91_33 word91_33 gnd C_wl
Rw92_33 word92_33 word91_33 R_wl
Cwl_92_33 word92_33 gnd C_wl
Rw93_33 word93_33 word92_33 R_wl
Cwl_93_33 word93_33 gnd C_wl
Rw94_33 word94_33 word93_33 R_wl
Cwl_94_33 word94_33 gnd C_wl
Rw95_33 word95_33 word94_33 R_wl
Cwl_95_33 word95_33 gnd C_wl
Rw96_33 word96_33 word95_33 R_wl
Cwl_96_33 word96_33 gnd C_wl
Rw97_33 word97_33 word96_33 R_wl
Cwl_97_33 word97_33 gnd C_wl
Rw98_33 word98_33 word97_33 R_wl
Cwl_98_33 word98_33 gnd C_wl
Rw99_33 word99_33 word98_33 R_wl
Cwl_99_33 word99_33 gnd C_wl
Vwl_34 word_34 0 0
Rw0_34 word_34 word0_34 R_wl
Cwl_0_34 word0_34 gnd C_wl
Rw1_34 word1_34 word0_34 R_wl
Cwl_1_34 word1_34 gnd C_wl
Rw2_34 word2_34 word1_34 R_wl
Cwl_2_34 word2_34 gnd C_wl
Rw3_34 word3_34 word2_34 R_wl
Cwl_3_34 word3_34 gnd C_wl
Rw4_34 word4_34 word3_34 R_wl
Cwl_4_34 word4_34 gnd C_wl
Rw5_34 word5_34 word4_34 R_wl
Cwl_5_34 word5_34 gnd C_wl
Rw6_34 word6_34 word5_34 R_wl
Cwl_6_34 word6_34 gnd C_wl
Rw7_34 word7_34 word6_34 R_wl
Cwl_7_34 word7_34 gnd C_wl
Rw8_34 word8_34 word7_34 R_wl
Cwl_8_34 word8_34 gnd C_wl
Rw9_34 word9_34 word8_34 R_wl
Cwl_9_34 word9_34 gnd C_wl
Rw10_34 word10_34 word9_34 R_wl
Cwl_10_34 word10_34 gnd C_wl
Rw11_34 word11_34 word10_34 R_wl
Cwl_11_34 word11_34 gnd C_wl
Rw12_34 word12_34 word11_34 R_wl
Cwl_12_34 word12_34 gnd C_wl
Rw13_34 word13_34 word12_34 R_wl
Cwl_13_34 word13_34 gnd C_wl
Rw14_34 word14_34 word13_34 R_wl
Cwl_14_34 word14_34 gnd C_wl
Rw15_34 word15_34 word14_34 R_wl
Cwl_15_34 word15_34 gnd C_wl
Rw16_34 word16_34 word15_34 R_wl
Cwl_16_34 word16_34 gnd C_wl
Rw17_34 word17_34 word16_34 R_wl
Cwl_17_34 word17_34 gnd C_wl
Rw18_34 word18_34 word17_34 R_wl
Cwl_18_34 word18_34 gnd C_wl
Rw19_34 word19_34 word18_34 R_wl
Cwl_19_34 word19_34 gnd C_wl
Rw20_34 word20_34 word19_34 R_wl
Cwl_20_34 word20_34 gnd C_wl
Rw21_34 word21_34 word20_34 R_wl
Cwl_21_34 word21_34 gnd C_wl
Rw22_34 word22_34 word21_34 R_wl
Cwl_22_34 word22_34 gnd C_wl
Rw23_34 word23_34 word22_34 R_wl
Cwl_23_34 word23_34 gnd C_wl
Rw24_34 word24_34 word23_34 R_wl
Cwl_24_34 word24_34 gnd C_wl
Rw25_34 word25_34 word24_34 R_wl
Cwl_25_34 word25_34 gnd C_wl
Rw26_34 word26_34 word25_34 R_wl
Cwl_26_34 word26_34 gnd C_wl
Rw27_34 word27_34 word26_34 R_wl
Cwl_27_34 word27_34 gnd C_wl
Rw28_34 word28_34 word27_34 R_wl
Cwl_28_34 word28_34 gnd C_wl
Rw29_34 word29_34 word28_34 R_wl
Cwl_29_34 word29_34 gnd C_wl
Rw30_34 word30_34 word29_34 R_wl
Cwl_30_34 word30_34 gnd C_wl
Rw31_34 word31_34 word30_34 R_wl
Cwl_31_34 word31_34 gnd C_wl
Rw32_34 word32_34 word31_34 R_wl
Cwl_32_34 word32_34 gnd C_wl
Rw33_34 word33_34 word32_34 R_wl
Cwl_33_34 word33_34 gnd C_wl
Rw34_34 word34_34 word33_34 R_wl
Cwl_34_34 word34_34 gnd C_wl
Rw35_34 word35_34 word34_34 R_wl
Cwl_35_34 word35_34 gnd C_wl
Rw36_34 word36_34 word35_34 R_wl
Cwl_36_34 word36_34 gnd C_wl
Rw37_34 word37_34 word36_34 R_wl
Cwl_37_34 word37_34 gnd C_wl
Rw38_34 word38_34 word37_34 R_wl
Cwl_38_34 word38_34 gnd C_wl
Rw39_34 word39_34 word38_34 R_wl
Cwl_39_34 word39_34 gnd C_wl
Rw40_34 word40_34 word39_34 R_wl
Cwl_40_34 word40_34 gnd C_wl
Rw41_34 word41_34 word40_34 R_wl
Cwl_41_34 word41_34 gnd C_wl
Rw42_34 word42_34 word41_34 R_wl
Cwl_42_34 word42_34 gnd C_wl
Rw43_34 word43_34 word42_34 R_wl
Cwl_43_34 word43_34 gnd C_wl
Rw44_34 word44_34 word43_34 R_wl
Cwl_44_34 word44_34 gnd C_wl
Rw45_34 word45_34 word44_34 R_wl
Cwl_45_34 word45_34 gnd C_wl
Rw46_34 word46_34 word45_34 R_wl
Cwl_46_34 word46_34 gnd C_wl
Rw47_34 word47_34 word46_34 R_wl
Cwl_47_34 word47_34 gnd C_wl
Rw48_34 word48_34 word47_34 R_wl
Cwl_48_34 word48_34 gnd C_wl
Rw49_34 word49_34 word48_34 R_wl
Cwl_49_34 word49_34 gnd C_wl
Rw50_34 word50_34 word49_34 R_wl
Cwl_50_34 word50_34 gnd C_wl
Rw51_34 word51_34 word50_34 R_wl
Cwl_51_34 word51_34 gnd C_wl
Rw52_34 word52_34 word51_34 R_wl
Cwl_52_34 word52_34 gnd C_wl
Rw53_34 word53_34 word52_34 R_wl
Cwl_53_34 word53_34 gnd C_wl
Rw54_34 word54_34 word53_34 R_wl
Cwl_54_34 word54_34 gnd C_wl
Rw55_34 word55_34 word54_34 R_wl
Cwl_55_34 word55_34 gnd C_wl
Rw56_34 word56_34 word55_34 R_wl
Cwl_56_34 word56_34 gnd C_wl
Rw57_34 word57_34 word56_34 R_wl
Cwl_57_34 word57_34 gnd C_wl
Rw58_34 word58_34 word57_34 R_wl
Cwl_58_34 word58_34 gnd C_wl
Rw59_34 word59_34 word58_34 R_wl
Cwl_59_34 word59_34 gnd C_wl
Rw60_34 word60_34 word59_34 R_wl
Cwl_60_34 word60_34 gnd C_wl
Rw61_34 word61_34 word60_34 R_wl
Cwl_61_34 word61_34 gnd C_wl
Rw62_34 word62_34 word61_34 R_wl
Cwl_62_34 word62_34 gnd C_wl
Rw63_34 word63_34 word62_34 R_wl
Cwl_63_34 word63_34 gnd C_wl
Rw64_34 word64_34 word63_34 R_wl
Cwl_64_34 word64_34 gnd C_wl
Rw65_34 word65_34 word64_34 R_wl
Cwl_65_34 word65_34 gnd C_wl
Rw66_34 word66_34 word65_34 R_wl
Cwl_66_34 word66_34 gnd C_wl
Rw67_34 word67_34 word66_34 R_wl
Cwl_67_34 word67_34 gnd C_wl
Rw68_34 word68_34 word67_34 R_wl
Cwl_68_34 word68_34 gnd C_wl
Rw69_34 word69_34 word68_34 R_wl
Cwl_69_34 word69_34 gnd C_wl
Rw70_34 word70_34 word69_34 R_wl
Cwl_70_34 word70_34 gnd C_wl
Rw71_34 word71_34 word70_34 R_wl
Cwl_71_34 word71_34 gnd C_wl
Rw72_34 word72_34 word71_34 R_wl
Cwl_72_34 word72_34 gnd C_wl
Rw73_34 word73_34 word72_34 R_wl
Cwl_73_34 word73_34 gnd C_wl
Rw74_34 word74_34 word73_34 R_wl
Cwl_74_34 word74_34 gnd C_wl
Rw75_34 word75_34 word74_34 R_wl
Cwl_75_34 word75_34 gnd C_wl
Rw76_34 word76_34 word75_34 R_wl
Cwl_76_34 word76_34 gnd C_wl
Rw77_34 word77_34 word76_34 R_wl
Cwl_77_34 word77_34 gnd C_wl
Rw78_34 word78_34 word77_34 R_wl
Cwl_78_34 word78_34 gnd C_wl
Rw79_34 word79_34 word78_34 R_wl
Cwl_79_34 word79_34 gnd C_wl
Rw80_34 word80_34 word79_34 R_wl
Cwl_80_34 word80_34 gnd C_wl
Rw81_34 word81_34 word80_34 R_wl
Cwl_81_34 word81_34 gnd C_wl
Rw82_34 word82_34 word81_34 R_wl
Cwl_82_34 word82_34 gnd C_wl
Rw83_34 word83_34 word82_34 R_wl
Cwl_83_34 word83_34 gnd C_wl
Rw84_34 word84_34 word83_34 R_wl
Cwl_84_34 word84_34 gnd C_wl
Rw85_34 word85_34 word84_34 R_wl
Cwl_85_34 word85_34 gnd C_wl
Rw86_34 word86_34 word85_34 R_wl
Cwl_86_34 word86_34 gnd C_wl
Rw87_34 word87_34 word86_34 R_wl
Cwl_87_34 word87_34 gnd C_wl
Rw88_34 word88_34 word87_34 R_wl
Cwl_88_34 word88_34 gnd C_wl
Rw89_34 word89_34 word88_34 R_wl
Cwl_89_34 word89_34 gnd C_wl
Rw90_34 word90_34 word89_34 R_wl
Cwl_90_34 word90_34 gnd C_wl
Rw91_34 word91_34 word90_34 R_wl
Cwl_91_34 word91_34 gnd C_wl
Rw92_34 word92_34 word91_34 R_wl
Cwl_92_34 word92_34 gnd C_wl
Rw93_34 word93_34 word92_34 R_wl
Cwl_93_34 word93_34 gnd C_wl
Rw94_34 word94_34 word93_34 R_wl
Cwl_94_34 word94_34 gnd C_wl
Rw95_34 word95_34 word94_34 R_wl
Cwl_95_34 word95_34 gnd C_wl
Rw96_34 word96_34 word95_34 R_wl
Cwl_96_34 word96_34 gnd C_wl
Rw97_34 word97_34 word96_34 R_wl
Cwl_97_34 word97_34 gnd C_wl
Rw98_34 word98_34 word97_34 R_wl
Cwl_98_34 word98_34 gnd C_wl
Rw99_34 word99_34 word98_34 R_wl
Cwl_99_34 word99_34 gnd C_wl
Vwl_35 word_35 0 0
Rw0_35 word_35 word0_35 R_wl
Cwl_0_35 word0_35 gnd C_wl
Rw1_35 word1_35 word0_35 R_wl
Cwl_1_35 word1_35 gnd C_wl
Rw2_35 word2_35 word1_35 R_wl
Cwl_2_35 word2_35 gnd C_wl
Rw3_35 word3_35 word2_35 R_wl
Cwl_3_35 word3_35 gnd C_wl
Rw4_35 word4_35 word3_35 R_wl
Cwl_4_35 word4_35 gnd C_wl
Rw5_35 word5_35 word4_35 R_wl
Cwl_5_35 word5_35 gnd C_wl
Rw6_35 word6_35 word5_35 R_wl
Cwl_6_35 word6_35 gnd C_wl
Rw7_35 word7_35 word6_35 R_wl
Cwl_7_35 word7_35 gnd C_wl
Rw8_35 word8_35 word7_35 R_wl
Cwl_8_35 word8_35 gnd C_wl
Rw9_35 word9_35 word8_35 R_wl
Cwl_9_35 word9_35 gnd C_wl
Rw10_35 word10_35 word9_35 R_wl
Cwl_10_35 word10_35 gnd C_wl
Rw11_35 word11_35 word10_35 R_wl
Cwl_11_35 word11_35 gnd C_wl
Rw12_35 word12_35 word11_35 R_wl
Cwl_12_35 word12_35 gnd C_wl
Rw13_35 word13_35 word12_35 R_wl
Cwl_13_35 word13_35 gnd C_wl
Rw14_35 word14_35 word13_35 R_wl
Cwl_14_35 word14_35 gnd C_wl
Rw15_35 word15_35 word14_35 R_wl
Cwl_15_35 word15_35 gnd C_wl
Rw16_35 word16_35 word15_35 R_wl
Cwl_16_35 word16_35 gnd C_wl
Rw17_35 word17_35 word16_35 R_wl
Cwl_17_35 word17_35 gnd C_wl
Rw18_35 word18_35 word17_35 R_wl
Cwl_18_35 word18_35 gnd C_wl
Rw19_35 word19_35 word18_35 R_wl
Cwl_19_35 word19_35 gnd C_wl
Rw20_35 word20_35 word19_35 R_wl
Cwl_20_35 word20_35 gnd C_wl
Rw21_35 word21_35 word20_35 R_wl
Cwl_21_35 word21_35 gnd C_wl
Rw22_35 word22_35 word21_35 R_wl
Cwl_22_35 word22_35 gnd C_wl
Rw23_35 word23_35 word22_35 R_wl
Cwl_23_35 word23_35 gnd C_wl
Rw24_35 word24_35 word23_35 R_wl
Cwl_24_35 word24_35 gnd C_wl
Rw25_35 word25_35 word24_35 R_wl
Cwl_25_35 word25_35 gnd C_wl
Rw26_35 word26_35 word25_35 R_wl
Cwl_26_35 word26_35 gnd C_wl
Rw27_35 word27_35 word26_35 R_wl
Cwl_27_35 word27_35 gnd C_wl
Rw28_35 word28_35 word27_35 R_wl
Cwl_28_35 word28_35 gnd C_wl
Rw29_35 word29_35 word28_35 R_wl
Cwl_29_35 word29_35 gnd C_wl
Rw30_35 word30_35 word29_35 R_wl
Cwl_30_35 word30_35 gnd C_wl
Rw31_35 word31_35 word30_35 R_wl
Cwl_31_35 word31_35 gnd C_wl
Rw32_35 word32_35 word31_35 R_wl
Cwl_32_35 word32_35 gnd C_wl
Rw33_35 word33_35 word32_35 R_wl
Cwl_33_35 word33_35 gnd C_wl
Rw34_35 word34_35 word33_35 R_wl
Cwl_34_35 word34_35 gnd C_wl
Rw35_35 word35_35 word34_35 R_wl
Cwl_35_35 word35_35 gnd C_wl
Rw36_35 word36_35 word35_35 R_wl
Cwl_36_35 word36_35 gnd C_wl
Rw37_35 word37_35 word36_35 R_wl
Cwl_37_35 word37_35 gnd C_wl
Rw38_35 word38_35 word37_35 R_wl
Cwl_38_35 word38_35 gnd C_wl
Rw39_35 word39_35 word38_35 R_wl
Cwl_39_35 word39_35 gnd C_wl
Rw40_35 word40_35 word39_35 R_wl
Cwl_40_35 word40_35 gnd C_wl
Rw41_35 word41_35 word40_35 R_wl
Cwl_41_35 word41_35 gnd C_wl
Rw42_35 word42_35 word41_35 R_wl
Cwl_42_35 word42_35 gnd C_wl
Rw43_35 word43_35 word42_35 R_wl
Cwl_43_35 word43_35 gnd C_wl
Rw44_35 word44_35 word43_35 R_wl
Cwl_44_35 word44_35 gnd C_wl
Rw45_35 word45_35 word44_35 R_wl
Cwl_45_35 word45_35 gnd C_wl
Rw46_35 word46_35 word45_35 R_wl
Cwl_46_35 word46_35 gnd C_wl
Rw47_35 word47_35 word46_35 R_wl
Cwl_47_35 word47_35 gnd C_wl
Rw48_35 word48_35 word47_35 R_wl
Cwl_48_35 word48_35 gnd C_wl
Rw49_35 word49_35 word48_35 R_wl
Cwl_49_35 word49_35 gnd C_wl
Rw50_35 word50_35 word49_35 R_wl
Cwl_50_35 word50_35 gnd C_wl
Rw51_35 word51_35 word50_35 R_wl
Cwl_51_35 word51_35 gnd C_wl
Rw52_35 word52_35 word51_35 R_wl
Cwl_52_35 word52_35 gnd C_wl
Rw53_35 word53_35 word52_35 R_wl
Cwl_53_35 word53_35 gnd C_wl
Rw54_35 word54_35 word53_35 R_wl
Cwl_54_35 word54_35 gnd C_wl
Rw55_35 word55_35 word54_35 R_wl
Cwl_55_35 word55_35 gnd C_wl
Rw56_35 word56_35 word55_35 R_wl
Cwl_56_35 word56_35 gnd C_wl
Rw57_35 word57_35 word56_35 R_wl
Cwl_57_35 word57_35 gnd C_wl
Rw58_35 word58_35 word57_35 R_wl
Cwl_58_35 word58_35 gnd C_wl
Rw59_35 word59_35 word58_35 R_wl
Cwl_59_35 word59_35 gnd C_wl
Rw60_35 word60_35 word59_35 R_wl
Cwl_60_35 word60_35 gnd C_wl
Rw61_35 word61_35 word60_35 R_wl
Cwl_61_35 word61_35 gnd C_wl
Rw62_35 word62_35 word61_35 R_wl
Cwl_62_35 word62_35 gnd C_wl
Rw63_35 word63_35 word62_35 R_wl
Cwl_63_35 word63_35 gnd C_wl
Rw64_35 word64_35 word63_35 R_wl
Cwl_64_35 word64_35 gnd C_wl
Rw65_35 word65_35 word64_35 R_wl
Cwl_65_35 word65_35 gnd C_wl
Rw66_35 word66_35 word65_35 R_wl
Cwl_66_35 word66_35 gnd C_wl
Rw67_35 word67_35 word66_35 R_wl
Cwl_67_35 word67_35 gnd C_wl
Rw68_35 word68_35 word67_35 R_wl
Cwl_68_35 word68_35 gnd C_wl
Rw69_35 word69_35 word68_35 R_wl
Cwl_69_35 word69_35 gnd C_wl
Rw70_35 word70_35 word69_35 R_wl
Cwl_70_35 word70_35 gnd C_wl
Rw71_35 word71_35 word70_35 R_wl
Cwl_71_35 word71_35 gnd C_wl
Rw72_35 word72_35 word71_35 R_wl
Cwl_72_35 word72_35 gnd C_wl
Rw73_35 word73_35 word72_35 R_wl
Cwl_73_35 word73_35 gnd C_wl
Rw74_35 word74_35 word73_35 R_wl
Cwl_74_35 word74_35 gnd C_wl
Rw75_35 word75_35 word74_35 R_wl
Cwl_75_35 word75_35 gnd C_wl
Rw76_35 word76_35 word75_35 R_wl
Cwl_76_35 word76_35 gnd C_wl
Rw77_35 word77_35 word76_35 R_wl
Cwl_77_35 word77_35 gnd C_wl
Rw78_35 word78_35 word77_35 R_wl
Cwl_78_35 word78_35 gnd C_wl
Rw79_35 word79_35 word78_35 R_wl
Cwl_79_35 word79_35 gnd C_wl
Rw80_35 word80_35 word79_35 R_wl
Cwl_80_35 word80_35 gnd C_wl
Rw81_35 word81_35 word80_35 R_wl
Cwl_81_35 word81_35 gnd C_wl
Rw82_35 word82_35 word81_35 R_wl
Cwl_82_35 word82_35 gnd C_wl
Rw83_35 word83_35 word82_35 R_wl
Cwl_83_35 word83_35 gnd C_wl
Rw84_35 word84_35 word83_35 R_wl
Cwl_84_35 word84_35 gnd C_wl
Rw85_35 word85_35 word84_35 R_wl
Cwl_85_35 word85_35 gnd C_wl
Rw86_35 word86_35 word85_35 R_wl
Cwl_86_35 word86_35 gnd C_wl
Rw87_35 word87_35 word86_35 R_wl
Cwl_87_35 word87_35 gnd C_wl
Rw88_35 word88_35 word87_35 R_wl
Cwl_88_35 word88_35 gnd C_wl
Rw89_35 word89_35 word88_35 R_wl
Cwl_89_35 word89_35 gnd C_wl
Rw90_35 word90_35 word89_35 R_wl
Cwl_90_35 word90_35 gnd C_wl
Rw91_35 word91_35 word90_35 R_wl
Cwl_91_35 word91_35 gnd C_wl
Rw92_35 word92_35 word91_35 R_wl
Cwl_92_35 word92_35 gnd C_wl
Rw93_35 word93_35 word92_35 R_wl
Cwl_93_35 word93_35 gnd C_wl
Rw94_35 word94_35 word93_35 R_wl
Cwl_94_35 word94_35 gnd C_wl
Rw95_35 word95_35 word94_35 R_wl
Cwl_95_35 word95_35 gnd C_wl
Rw96_35 word96_35 word95_35 R_wl
Cwl_96_35 word96_35 gnd C_wl
Rw97_35 word97_35 word96_35 R_wl
Cwl_97_35 word97_35 gnd C_wl
Rw98_35 word98_35 word97_35 R_wl
Cwl_98_35 word98_35 gnd C_wl
Rw99_35 word99_35 word98_35 R_wl
Cwl_99_35 word99_35 gnd C_wl
Vwl_36 word_36 0 0
Rw0_36 word_36 word0_36 R_wl
Cwl_0_36 word0_36 gnd C_wl
Rw1_36 word1_36 word0_36 R_wl
Cwl_1_36 word1_36 gnd C_wl
Rw2_36 word2_36 word1_36 R_wl
Cwl_2_36 word2_36 gnd C_wl
Rw3_36 word3_36 word2_36 R_wl
Cwl_3_36 word3_36 gnd C_wl
Rw4_36 word4_36 word3_36 R_wl
Cwl_4_36 word4_36 gnd C_wl
Rw5_36 word5_36 word4_36 R_wl
Cwl_5_36 word5_36 gnd C_wl
Rw6_36 word6_36 word5_36 R_wl
Cwl_6_36 word6_36 gnd C_wl
Rw7_36 word7_36 word6_36 R_wl
Cwl_7_36 word7_36 gnd C_wl
Rw8_36 word8_36 word7_36 R_wl
Cwl_8_36 word8_36 gnd C_wl
Rw9_36 word9_36 word8_36 R_wl
Cwl_9_36 word9_36 gnd C_wl
Rw10_36 word10_36 word9_36 R_wl
Cwl_10_36 word10_36 gnd C_wl
Rw11_36 word11_36 word10_36 R_wl
Cwl_11_36 word11_36 gnd C_wl
Rw12_36 word12_36 word11_36 R_wl
Cwl_12_36 word12_36 gnd C_wl
Rw13_36 word13_36 word12_36 R_wl
Cwl_13_36 word13_36 gnd C_wl
Rw14_36 word14_36 word13_36 R_wl
Cwl_14_36 word14_36 gnd C_wl
Rw15_36 word15_36 word14_36 R_wl
Cwl_15_36 word15_36 gnd C_wl
Rw16_36 word16_36 word15_36 R_wl
Cwl_16_36 word16_36 gnd C_wl
Rw17_36 word17_36 word16_36 R_wl
Cwl_17_36 word17_36 gnd C_wl
Rw18_36 word18_36 word17_36 R_wl
Cwl_18_36 word18_36 gnd C_wl
Rw19_36 word19_36 word18_36 R_wl
Cwl_19_36 word19_36 gnd C_wl
Rw20_36 word20_36 word19_36 R_wl
Cwl_20_36 word20_36 gnd C_wl
Rw21_36 word21_36 word20_36 R_wl
Cwl_21_36 word21_36 gnd C_wl
Rw22_36 word22_36 word21_36 R_wl
Cwl_22_36 word22_36 gnd C_wl
Rw23_36 word23_36 word22_36 R_wl
Cwl_23_36 word23_36 gnd C_wl
Rw24_36 word24_36 word23_36 R_wl
Cwl_24_36 word24_36 gnd C_wl
Rw25_36 word25_36 word24_36 R_wl
Cwl_25_36 word25_36 gnd C_wl
Rw26_36 word26_36 word25_36 R_wl
Cwl_26_36 word26_36 gnd C_wl
Rw27_36 word27_36 word26_36 R_wl
Cwl_27_36 word27_36 gnd C_wl
Rw28_36 word28_36 word27_36 R_wl
Cwl_28_36 word28_36 gnd C_wl
Rw29_36 word29_36 word28_36 R_wl
Cwl_29_36 word29_36 gnd C_wl
Rw30_36 word30_36 word29_36 R_wl
Cwl_30_36 word30_36 gnd C_wl
Rw31_36 word31_36 word30_36 R_wl
Cwl_31_36 word31_36 gnd C_wl
Rw32_36 word32_36 word31_36 R_wl
Cwl_32_36 word32_36 gnd C_wl
Rw33_36 word33_36 word32_36 R_wl
Cwl_33_36 word33_36 gnd C_wl
Rw34_36 word34_36 word33_36 R_wl
Cwl_34_36 word34_36 gnd C_wl
Rw35_36 word35_36 word34_36 R_wl
Cwl_35_36 word35_36 gnd C_wl
Rw36_36 word36_36 word35_36 R_wl
Cwl_36_36 word36_36 gnd C_wl
Rw37_36 word37_36 word36_36 R_wl
Cwl_37_36 word37_36 gnd C_wl
Rw38_36 word38_36 word37_36 R_wl
Cwl_38_36 word38_36 gnd C_wl
Rw39_36 word39_36 word38_36 R_wl
Cwl_39_36 word39_36 gnd C_wl
Rw40_36 word40_36 word39_36 R_wl
Cwl_40_36 word40_36 gnd C_wl
Rw41_36 word41_36 word40_36 R_wl
Cwl_41_36 word41_36 gnd C_wl
Rw42_36 word42_36 word41_36 R_wl
Cwl_42_36 word42_36 gnd C_wl
Rw43_36 word43_36 word42_36 R_wl
Cwl_43_36 word43_36 gnd C_wl
Rw44_36 word44_36 word43_36 R_wl
Cwl_44_36 word44_36 gnd C_wl
Rw45_36 word45_36 word44_36 R_wl
Cwl_45_36 word45_36 gnd C_wl
Rw46_36 word46_36 word45_36 R_wl
Cwl_46_36 word46_36 gnd C_wl
Rw47_36 word47_36 word46_36 R_wl
Cwl_47_36 word47_36 gnd C_wl
Rw48_36 word48_36 word47_36 R_wl
Cwl_48_36 word48_36 gnd C_wl
Rw49_36 word49_36 word48_36 R_wl
Cwl_49_36 word49_36 gnd C_wl
Rw50_36 word50_36 word49_36 R_wl
Cwl_50_36 word50_36 gnd C_wl
Rw51_36 word51_36 word50_36 R_wl
Cwl_51_36 word51_36 gnd C_wl
Rw52_36 word52_36 word51_36 R_wl
Cwl_52_36 word52_36 gnd C_wl
Rw53_36 word53_36 word52_36 R_wl
Cwl_53_36 word53_36 gnd C_wl
Rw54_36 word54_36 word53_36 R_wl
Cwl_54_36 word54_36 gnd C_wl
Rw55_36 word55_36 word54_36 R_wl
Cwl_55_36 word55_36 gnd C_wl
Rw56_36 word56_36 word55_36 R_wl
Cwl_56_36 word56_36 gnd C_wl
Rw57_36 word57_36 word56_36 R_wl
Cwl_57_36 word57_36 gnd C_wl
Rw58_36 word58_36 word57_36 R_wl
Cwl_58_36 word58_36 gnd C_wl
Rw59_36 word59_36 word58_36 R_wl
Cwl_59_36 word59_36 gnd C_wl
Rw60_36 word60_36 word59_36 R_wl
Cwl_60_36 word60_36 gnd C_wl
Rw61_36 word61_36 word60_36 R_wl
Cwl_61_36 word61_36 gnd C_wl
Rw62_36 word62_36 word61_36 R_wl
Cwl_62_36 word62_36 gnd C_wl
Rw63_36 word63_36 word62_36 R_wl
Cwl_63_36 word63_36 gnd C_wl
Rw64_36 word64_36 word63_36 R_wl
Cwl_64_36 word64_36 gnd C_wl
Rw65_36 word65_36 word64_36 R_wl
Cwl_65_36 word65_36 gnd C_wl
Rw66_36 word66_36 word65_36 R_wl
Cwl_66_36 word66_36 gnd C_wl
Rw67_36 word67_36 word66_36 R_wl
Cwl_67_36 word67_36 gnd C_wl
Rw68_36 word68_36 word67_36 R_wl
Cwl_68_36 word68_36 gnd C_wl
Rw69_36 word69_36 word68_36 R_wl
Cwl_69_36 word69_36 gnd C_wl
Rw70_36 word70_36 word69_36 R_wl
Cwl_70_36 word70_36 gnd C_wl
Rw71_36 word71_36 word70_36 R_wl
Cwl_71_36 word71_36 gnd C_wl
Rw72_36 word72_36 word71_36 R_wl
Cwl_72_36 word72_36 gnd C_wl
Rw73_36 word73_36 word72_36 R_wl
Cwl_73_36 word73_36 gnd C_wl
Rw74_36 word74_36 word73_36 R_wl
Cwl_74_36 word74_36 gnd C_wl
Rw75_36 word75_36 word74_36 R_wl
Cwl_75_36 word75_36 gnd C_wl
Rw76_36 word76_36 word75_36 R_wl
Cwl_76_36 word76_36 gnd C_wl
Rw77_36 word77_36 word76_36 R_wl
Cwl_77_36 word77_36 gnd C_wl
Rw78_36 word78_36 word77_36 R_wl
Cwl_78_36 word78_36 gnd C_wl
Rw79_36 word79_36 word78_36 R_wl
Cwl_79_36 word79_36 gnd C_wl
Rw80_36 word80_36 word79_36 R_wl
Cwl_80_36 word80_36 gnd C_wl
Rw81_36 word81_36 word80_36 R_wl
Cwl_81_36 word81_36 gnd C_wl
Rw82_36 word82_36 word81_36 R_wl
Cwl_82_36 word82_36 gnd C_wl
Rw83_36 word83_36 word82_36 R_wl
Cwl_83_36 word83_36 gnd C_wl
Rw84_36 word84_36 word83_36 R_wl
Cwl_84_36 word84_36 gnd C_wl
Rw85_36 word85_36 word84_36 R_wl
Cwl_85_36 word85_36 gnd C_wl
Rw86_36 word86_36 word85_36 R_wl
Cwl_86_36 word86_36 gnd C_wl
Rw87_36 word87_36 word86_36 R_wl
Cwl_87_36 word87_36 gnd C_wl
Rw88_36 word88_36 word87_36 R_wl
Cwl_88_36 word88_36 gnd C_wl
Rw89_36 word89_36 word88_36 R_wl
Cwl_89_36 word89_36 gnd C_wl
Rw90_36 word90_36 word89_36 R_wl
Cwl_90_36 word90_36 gnd C_wl
Rw91_36 word91_36 word90_36 R_wl
Cwl_91_36 word91_36 gnd C_wl
Rw92_36 word92_36 word91_36 R_wl
Cwl_92_36 word92_36 gnd C_wl
Rw93_36 word93_36 word92_36 R_wl
Cwl_93_36 word93_36 gnd C_wl
Rw94_36 word94_36 word93_36 R_wl
Cwl_94_36 word94_36 gnd C_wl
Rw95_36 word95_36 word94_36 R_wl
Cwl_95_36 word95_36 gnd C_wl
Rw96_36 word96_36 word95_36 R_wl
Cwl_96_36 word96_36 gnd C_wl
Rw97_36 word97_36 word96_36 R_wl
Cwl_97_36 word97_36 gnd C_wl
Rw98_36 word98_36 word97_36 R_wl
Cwl_98_36 word98_36 gnd C_wl
Rw99_36 word99_36 word98_36 R_wl
Cwl_99_36 word99_36 gnd C_wl
Vwl_37 word_37 0 0
Rw0_37 word_37 word0_37 R_wl
Cwl_0_37 word0_37 gnd C_wl
Rw1_37 word1_37 word0_37 R_wl
Cwl_1_37 word1_37 gnd C_wl
Rw2_37 word2_37 word1_37 R_wl
Cwl_2_37 word2_37 gnd C_wl
Rw3_37 word3_37 word2_37 R_wl
Cwl_3_37 word3_37 gnd C_wl
Rw4_37 word4_37 word3_37 R_wl
Cwl_4_37 word4_37 gnd C_wl
Rw5_37 word5_37 word4_37 R_wl
Cwl_5_37 word5_37 gnd C_wl
Rw6_37 word6_37 word5_37 R_wl
Cwl_6_37 word6_37 gnd C_wl
Rw7_37 word7_37 word6_37 R_wl
Cwl_7_37 word7_37 gnd C_wl
Rw8_37 word8_37 word7_37 R_wl
Cwl_8_37 word8_37 gnd C_wl
Rw9_37 word9_37 word8_37 R_wl
Cwl_9_37 word9_37 gnd C_wl
Rw10_37 word10_37 word9_37 R_wl
Cwl_10_37 word10_37 gnd C_wl
Rw11_37 word11_37 word10_37 R_wl
Cwl_11_37 word11_37 gnd C_wl
Rw12_37 word12_37 word11_37 R_wl
Cwl_12_37 word12_37 gnd C_wl
Rw13_37 word13_37 word12_37 R_wl
Cwl_13_37 word13_37 gnd C_wl
Rw14_37 word14_37 word13_37 R_wl
Cwl_14_37 word14_37 gnd C_wl
Rw15_37 word15_37 word14_37 R_wl
Cwl_15_37 word15_37 gnd C_wl
Rw16_37 word16_37 word15_37 R_wl
Cwl_16_37 word16_37 gnd C_wl
Rw17_37 word17_37 word16_37 R_wl
Cwl_17_37 word17_37 gnd C_wl
Rw18_37 word18_37 word17_37 R_wl
Cwl_18_37 word18_37 gnd C_wl
Rw19_37 word19_37 word18_37 R_wl
Cwl_19_37 word19_37 gnd C_wl
Rw20_37 word20_37 word19_37 R_wl
Cwl_20_37 word20_37 gnd C_wl
Rw21_37 word21_37 word20_37 R_wl
Cwl_21_37 word21_37 gnd C_wl
Rw22_37 word22_37 word21_37 R_wl
Cwl_22_37 word22_37 gnd C_wl
Rw23_37 word23_37 word22_37 R_wl
Cwl_23_37 word23_37 gnd C_wl
Rw24_37 word24_37 word23_37 R_wl
Cwl_24_37 word24_37 gnd C_wl
Rw25_37 word25_37 word24_37 R_wl
Cwl_25_37 word25_37 gnd C_wl
Rw26_37 word26_37 word25_37 R_wl
Cwl_26_37 word26_37 gnd C_wl
Rw27_37 word27_37 word26_37 R_wl
Cwl_27_37 word27_37 gnd C_wl
Rw28_37 word28_37 word27_37 R_wl
Cwl_28_37 word28_37 gnd C_wl
Rw29_37 word29_37 word28_37 R_wl
Cwl_29_37 word29_37 gnd C_wl
Rw30_37 word30_37 word29_37 R_wl
Cwl_30_37 word30_37 gnd C_wl
Rw31_37 word31_37 word30_37 R_wl
Cwl_31_37 word31_37 gnd C_wl
Rw32_37 word32_37 word31_37 R_wl
Cwl_32_37 word32_37 gnd C_wl
Rw33_37 word33_37 word32_37 R_wl
Cwl_33_37 word33_37 gnd C_wl
Rw34_37 word34_37 word33_37 R_wl
Cwl_34_37 word34_37 gnd C_wl
Rw35_37 word35_37 word34_37 R_wl
Cwl_35_37 word35_37 gnd C_wl
Rw36_37 word36_37 word35_37 R_wl
Cwl_36_37 word36_37 gnd C_wl
Rw37_37 word37_37 word36_37 R_wl
Cwl_37_37 word37_37 gnd C_wl
Rw38_37 word38_37 word37_37 R_wl
Cwl_38_37 word38_37 gnd C_wl
Rw39_37 word39_37 word38_37 R_wl
Cwl_39_37 word39_37 gnd C_wl
Rw40_37 word40_37 word39_37 R_wl
Cwl_40_37 word40_37 gnd C_wl
Rw41_37 word41_37 word40_37 R_wl
Cwl_41_37 word41_37 gnd C_wl
Rw42_37 word42_37 word41_37 R_wl
Cwl_42_37 word42_37 gnd C_wl
Rw43_37 word43_37 word42_37 R_wl
Cwl_43_37 word43_37 gnd C_wl
Rw44_37 word44_37 word43_37 R_wl
Cwl_44_37 word44_37 gnd C_wl
Rw45_37 word45_37 word44_37 R_wl
Cwl_45_37 word45_37 gnd C_wl
Rw46_37 word46_37 word45_37 R_wl
Cwl_46_37 word46_37 gnd C_wl
Rw47_37 word47_37 word46_37 R_wl
Cwl_47_37 word47_37 gnd C_wl
Rw48_37 word48_37 word47_37 R_wl
Cwl_48_37 word48_37 gnd C_wl
Rw49_37 word49_37 word48_37 R_wl
Cwl_49_37 word49_37 gnd C_wl
Rw50_37 word50_37 word49_37 R_wl
Cwl_50_37 word50_37 gnd C_wl
Rw51_37 word51_37 word50_37 R_wl
Cwl_51_37 word51_37 gnd C_wl
Rw52_37 word52_37 word51_37 R_wl
Cwl_52_37 word52_37 gnd C_wl
Rw53_37 word53_37 word52_37 R_wl
Cwl_53_37 word53_37 gnd C_wl
Rw54_37 word54_37 word53_37 R_wl
Cwl_54_37 word54_37 gnd C_wl
Rw55_37 word55_37 word54_37 R_wl
Cwl_55_37 word55_37 gnd C_wl
Rw56_37 word56_37 word55_37 R_wl
Cwl_56_37 word56_37 gnd C_wl
Rw57_37 word57_37 word56_37 R_wl
Cwl_57_37 word57_37 gnd C_wl
Rw58_37 word58_37 word57_37 R_wl
Cwl_58_37 word58_37 gnd C_wl
Rw59_37 word59_37 word58_37 R_wl
Cwl_59_37 word59_37 gnd C_wl
Rw60_37 word60_37 word59_37 R_wl
Cwl_60_37 word60_37 gnd C_wl
Rw61_37 word61_37 word60_37 R_wl
Cwl_61_37 word61_37 gnd C_wl
Rw62_37 word62_37 word61_37 R_wl
Cwl_62_37 word62_37 gnd C_wl
Rw63_37 word63_37 word62_37 R_wl
Cwl_63_37 word63_37 gnd C_wl
Rw64_37 word64_37 word63_37 R_wl
Cwl_64_37 word64_37 gnd C_wl
Rw65_37 word65_37 word64_37 R_wl
Cwl_65_37 word65_37 gnd C_wl
Rw66_37 word66_37 word65_37 R_wl
Cwl_66_37 word66_37 gnd C_wl
Rw67_37 word67_37 word66_37 R_wl
Cwl_67_37 word67_37 gnd C_wl
Rw68_37 word68_37 word67_37 R_wl
Cwl_68_37 word68_37 gnd C_wl
Rw69_37 word69_37 word68_37 R_wl
Cwl_69_37 word69_37 gnd C_wl
Rw70_37 word70_37 word69_37 R_wl
Cwl_70_37 word70_37 gnd C_wl
Rw71_37 word71_37 word70_37 R_wl
Cwl_71_37 word71_37 gnd C_wl
Rw72_37 word72_37 word71_37 R_wl
Cwl_72_37 word72_37 gnd C_wl
Rw73_37 word73_37 word72_37 R_wl
Cwl_73_37 word73_37 gnd C_wl
Rw74_37 word74_37 word73_37 R_wl
Cwl_74_37 word74_37 gnd C_wl
Rw75_37 word75_37 word74_37 R_wl
Cwl_75_37 word75_37 gnd C_wl
Rw76_37 word76_37 word75_37 R_wl
Cwl_76_37 word76_37 gnd C_wl
Rw77_37 word77_37 word76_37 R_wl
Cwl_77_37 word77_37 gnd C_wl
Rw78_37 word78_37 word77_37 R_wl
Cwl_78_37 word78_37 gnd C_wl
Rw79_37 word79_37 word78_37 R_wl
Cwl_79_37 word79_37 gnd C_wl
Rw80_37 word80_37 word79_37 R_wl
Cwl_80_37 word80_37 gnd C_wl
Rw81_37 word81_37 word80_37 R_wl
Cwl_81_37 word81_37 gnd C_wl
Rw82_37 word82_37 word81_37 R_wl
Cwl_82_37 word82_37 gnd C_wl
Rw83_37 word83_37 word82_37 R_wl
Cwl_83_37 word83_37 gnd C_wl
Rw84_37 word84_37 word83_37 R_wl
Cwl_84_37 word84_37 gnd C_wl
Rw85_37 word85_37 word84_37 R_wl
Cwl_85_37 word85_37 gnd C_wl
Rw86_37 word86_37 word85_37 R_wl
Cwl_86_37 word86_37 gnd C_wl
Rw87_37 word87_37 word86_37 R_wl
Cwl_87_37 word87_37 gnd C_wl
Rw88_37 word88_37 word87_37 R_wl
Cwl_88_37 word88_37 gnd C_wl
Rw89_37 word89_37 word88_37 R_wl
Cwl_89_37 word89_37 gnd C_wl
Rw90_37 word90_37 word89_37 R_wl
Cwl_90_37 word90_37 gnd C_wl
Rw91_37 word91_37 word90_37 R_wl
Cwl_91_37 word91_37 gnd C_wl
Rw92_37 word92_37 word91_37 R_wl
Cwl_92_37 word92_37 gnd C_wl
Rw93_37 word93_37 word92_37 R_wl
Cwl_93_37 word93_37 gnd C_wl
Rw94_37 word94_37 word93_37 R_wl
Cwl_94_37 word94_37 gnd C_wl
Rw95_37 word95_37 word94_37 R_wl
Cwl_95_37 word95_37 gnd C_wl
Rw96_37 word96_37 word95_37 R_wl
Cwl_96_37 word96_37 gnd C_wl
Rw97_37 word97_37 word96_37 R_wl
Cwl_97_37 word97_37 gnd C_wl
Rw98_37 word98_37 word97_37 R_wl
Cwl_98_37 word98_37 gnd C_wl
Rw99_37 word99_37 word98_37 R_wl
Cwl_99_37 word99_37 gnd C_wl
Vwl_38 word_38 0 0
Rw0_38 word_38 word0_38 R_wl
Cwl_0_38 word0_38 gnd C_wl
Rw1_38 word1_38 word0_38 R_wl
Cwl_1_38 word1_38 gnd C_wl
Rw2_38 word2_38 word1_38 R_wl
Cwl_2_38 word2_38 gnd C_wl
Rw3_38 word3_38 word2_38 R_wl
Cwl_3_38 word3_38 gnd C_wl
Rw4_38 word4_38 word3_38 R_wl
Cwl_4_38 word4_38 gnd C_wl
Rw5_38 word5_38 word4_38 R_wl
Cwl_5_38 word5_38 gnd C_wl
Rw6_38 word6_38 word5_38 R_wl
Cwl_6_38 word6_38 gnd C_wl
Rw7_38 word7_38 word6_38 R_wl
Cwl_7_38 word7_38 gnd C_wl
Rw8_38 word8_38 word7_38 R_wl
Cwl_8_38 word8_38 gnd C_wl
Rw9_38 word9_38 word8_38 R_wl
Cwl_9_38 word9_38 gnd C_wl
Rw10_38 word10_38 word9_38 R_wl
Cwl_10_38 word10_38 gnd C_wl
Rw11_38 word11_38 word10_38 R_wl
Cwl_11_38 word11_38 gnd C_wl
Rw12_38 word12_38 word11_38 R_wl
Cwl_12_38 word12_38 gnd C_wl
Rw13_38 word13_38 word12_38 R_wl
Cwl_13_38 word13_38 gnd C_wl
Rw14_38 word14_38 word13_38 R_wl
Cwl_14_38 word14_38 gnd C_wl
Rw15_38 word15_38 word14_38 R_wl
Cwl_15_38 word15_38 gnd C_wl
Rw16_38 word16_38 word15_38 R_wl
Cwl_16_38 word16_38 gnd C_wl
Rw17_38 word17_38 word16_38 R_wl
Cwl_17_38 word17_38 gnd C_wl
Rw18_38 word18_38 word17_38 R_wl
Cwl_18_38 word18_38 gnd C_wl
Rw19_38 word19_38 word18_38 R_wl
Cwl_19_38 word19_38 gnd C_wl
Rw20_38 word20_38 word19_38 R_wl
Cwl_20_38 word20_38 gnd C_wl
Rw21_38 word21_38 word20_38 R_wl
Cwl_21_38 word21_38 gnd C_wl
Rw22_38 word22_38 word21_38 R_wl
Cwl_22_38 word22_38 gnd C_wl
Rw23_38 word23_38 word22_38 R_wl
Cwl_23_38 word23_38 gnd C_wl
Rw24_38 word24_38 word23_38 R_wl
Cwl_24_38 word24_38 gnd C_wl
Rw25_38 word25_38 word24_38 R_wl
Cwl_25_38 word25_38 gnd C_wl
Rw26_38 word26_38 word25_38 R_wl
Cwl_26_38 word26_38 gnd C_wl
Rw27_38 word27_38 word26_38 R_wl
Cwl_27_38 word27_38 gnd C_wl
Rw28_38 word28_38 word27_38 R_wl
Cwl_28_38 word28_38 gnd C_wl
Rw29_38 word29_38 word28_38 R_wl
Cwl_29_38 word29_38 gnd C_wl
Rw30_38 word30_38 word29_38 R_wl
Cwl_30_38 word30_38 gnd C_wl
Rw31_38 word31_38 word30_38 R_wl
Cwl_31_38 word31_38 gnd C_wl
Rw32_38 word32_38 word31_38 R_wl
Cwl_32_38 word32_38 gnd C_wl
Rw33_38 word33_38 word32_38 R_wl
Cwl_33_38 word33_38 gnd C_wl
Rw34_38 word34_38 word33_38 R_wl
Cwl_34_38 word34_38 gnd C_wl
Rw35_38 word35_38 word34_38 R_wl
Cwl_35_38 word35_38 gnd C_wl
Rw36_38 word36_38 word35_38 R_wl
Cwl_36_38 word36_38 gnd C_wl
Rw37_38 word37_38 word36_38 R_wl
Cwl_37_38 word37_38 gnd C_wl
Rw38_38 word38_38 word37_38 R_wl
Cwl_38_38 word38_38 gnd C_wl
Rw39_38 word39_38 word38_38 R_wl
Cwl_39_38 word39_38 gnd C_wl
Rw40_38 word40_38 word39_38 R_wl
Cwl_40_38 word40_38 gnd C_wl
Rw41_38 word41_38 word40_38 R_wl
Cwl_41_38 word41_38 gnd C_wl
Rw42_38 word42_38 word41_38 R_wl
Cwl_42_38 word42_38 gnd C_wl
Rw43_38 word43_38 word42_38 R_wl
Cwl_43_38 word43_38 gnd C_wl
Rw44_38 word44_38 word43_38 R_wl
Cwl_44_38 word44_38 gnd C_wl
Rw45_38 word45_38 word44_38 R_wl
Cwl_45_38 word45_38 gnd C_wl
Rw46_38 word46_38 word45_38 R_wl
Cwl_46_38 word46_38 gnd C_wl
Rw47_38 word47_38 word46_38 R_wl
Cwl_47_38 word47_38 gnd C_wl
Rw48_38 word48_38 word47_38 R_wl
Cwl_48_38 word48_38 gnd C_wl
Rw49_38 word49_38 word48_38 R_wl
Cwl_49_38 word49_38 gnd C_wl
Rw50_38 word50_38 word49_38 R_wl
Cwl_50_38 word50_38 gnd C_wl
Rw51_38 word51_38 word50_38 R_wl
Cwl_51_38 word51_38 gnd C_wl
Rw52_38 word52_38 word51_38 R_wl
Cwl_52_38 word52_38 gnd C_wl
Rw53_38 word53_38 word52_38 R_wl
Cwl_53_38 word53_38 gnd C_wl
Rw54_38 word54_38 word53_38 R_wl
Cwl_54_38 word54_38 gnd C_wl
Rw55_38 word55_38 word54_38 R_wl
Cwl_55_38 word55_38 gnd C_wl
Rw56_38 word56_38 word55_38 R_wl
Cwl_56_38 word56_38 gnd C_wl
Rw57_38 word57_38 word56_38 R_wl
Cwl_57_38 word57_38 gnd C_wl
Rw58_38 word58_38 word57_38 R_wl
Cwl_58_38 word58_38 gnd C_wl
Rw59_38 word59_38 word58_38 R_wl
Cwl_59_38 word59_38 gnd C_wl
Rw60_38 word60_38 word59_38 R_wl
Cwl_60_38 word60_38 gnd C_wl
Rw61_38 word61_38 word60_38 R_wl
Cwl_61_38 word61_38 gnd C_wl
Rw62_38 word62_38 word61_38 R_wl
Cwl_62_38 word62_38 gnd C_wl
Rw63_38 word63_38 word62_38 R_wl
Cwl_63_38 word63_38 gnd C_wl
Rw64_38 word64_38 word63_38 R_wl
Cwl_64_38 word64_38 gnd C_wl
Rw65_38 word65_38 word64_38 R_wl
Cwl_65_38 word65_38 gnd C_wl
Rw66_38 word66_38 word65_38 R_wl
Cwl_66_38 word66_38 gnd C_wl
Rw67_38 word67_38 word66_38 R_wl
Cwl_67_38 word67_38 gnd C_wl
Rw68_38 word68_38 word67_38 R_wl
Cwl_68_38 word68_38 gnd C_wl
Rw69_38 word69_38 word68_38 R_wl
Cwl_69_38 word69_38 gnd C_wl
Rw70_38 word70_38 word69_38 R_wl
Cwl_70_38 word70_38 gnd C_wl
Rw71_38 word71_38 word70_38 R_wl
Cwl_71_38 word71_38 gnd C_wl
Rw72_38 word72_38 word71_38 R_wl
Cwl_72_38 word72_38 gnd C_wl
Rw73_38 word73_38 word72_38 R_wl
Cwl_73_38 word73_38 gnd C_wl
Rw74_38 word74_38 word73_38 R_wl
Cwl_74_38 word74_38 gnd C_wl
Rw75_38 word75_38 word74_38 R_wl
Cwl_75_38 word75_38 gnd C_wl
Rw76_38 word76_38 word75_38 R_wl
Cwl_76_38 word76_38 gnd C_wl
Rw77_38 word77_38 word76_38 R_wl
Cwl_77_38 word77_38 gnd C_wl
Rw78_38 word78_38 word77_38 R_wl
Cwl_78_38 word78_38 gnd C_wl
Rw79_38 word79_38 word78_38 R_wl
Cwl_79_38 word79_38 gnd C_wl
Rw80_38 word80_38 word79_38 R_wl
Cwl_80_38 word80_38 gnd C_wl
Rw81_38 word81_38 word80_38 R_wl
Cwl_81_38 word81_38 gnd C_wl
Rw82_38 word82_38 word81_38 R_wl
Cwl_82_38 word82_38 gnd C_wl
Rw83_38 word83_38 word82_38 R_wl
Cwl_83_38 word83_38 gnd C_wl
Rw84_38 word84_38 word83_38 R_wl
Cwl_84_38 word84_38 gnd C_wl
Rw85_38 word85_38 word84_38 R_wl
Cwl_85_38 word85_38 gnd C_wl
Rw86_38 word86_38 word85_38 R_wl
Cwl_86_38 word86_38 gnd C_wl
Rw87_38 word87_38 word86_38 R_wl
Cwl_87_38 word87_38 gnd C_wl
Rw88_38 word88_38 word87_38 R_wl
Cwl_88_38 word88_38 gnd C_wl
Rw89_38 word89_38 word88_38 R_wl
Cwl_89_38 word89_38 gnd C_wl
Rw90_38 word90_38 word89_38 R_wl
Cwl_90_38 word90_38 gnd C_wl
Rw91_38 word91_38 word90_38 R_wl
Cwl_91_38 word91_38 gnd C_wl
Rw92_38 word92_38 word91_38 R_wl
Cwl_92_38 word92_38 gnd C_wl
Rw93_38 word93_38 word92_38 R_wl
Cwl_93_38 word93_38 gnd C_wl
Rw94_38 word94_38 word93_38 R_wl
Cwl_94_38 word94_38 gnd C_wl
Rw95_38 word95_38 word94_38 R_wl
Cwl_95_38 word95_38 gnd C_wl
Rw96_38 word96_38 word95_38 R_wl
Cwl_96_38 word96_38 gnd C_wl
Rw97_38 word97_38 word96_38 R_wl
Cwl_97_38 word97_38 gnd C_wl
Rw98_38 word98_38 word97_38 R_wl
Cwl_98_38 word98_38 gnd C_wl
Rw99_38 word99_38 word98_38 R_wl
Cwl_99_38 word99_38 gnd C_wl
Vwl_39 word_39 0 0
Rw0_39 word_39 word0_39 R_wl
Cwl_0_39 word0_39 gnd C_wl
Rw1_39 word1_39 word0_39 R_wl
Cwl_1_39 word1_39 gnd C_wl
Rw2_39 word2_39 word1_39 R_wl
Cwl_2_39 word2_39 gnd C_wl
Rw3_39 word3_39 word2_39 R_wl
Cwl_3_39 word3_39 gnd C_wl
Rw4_39 word4_39 word3_39 R_wl
Cwl_4_39 word4_39 gnd C_wl
Rw5_39 word5_39 word4_39 R_wl
Cwl_5_39 word5_39 gnd C_wl
Rw6_39 word6_39 word5_39 R_wl
Cwl_6_39 word6_39 gnd C_wl
Rw7_39 word7_39 word6_39 R_wl
Cwl_7_39 word7_39 gnd C_wl
Rw8_39 word8_39 word7_39 R_wl
Cwl_8_39 word8_39 gnd C_wl
Rw9_39 word9_39 word8_39 R_wl
Cwl_9_39 word9_39 gnd C_wl
Rw10_39 word10_39 word9_39 R_wl
Cwl_10_39 word10_39 gnd C_wl
Rw11_39 word11_39 word10_39 R_wl
Cwl_11_39 word11_39 gnd C_wl
Rw12_39 word12_39 word11_39 R_wl
Cwl_12_39 word12_39 gnd C_wl
Rw13_39 word13_39 word12_39 R_wl
Cwl_13_39 word13_39 gnd C_wl
Rw14_39 word14_39 word13_39 R_wl
Cwl_14_39 word14_39 gnd C_wl
Rw15_39 word15_39 word14_39 R_wl
Cwl_15_39 word15_39 gnd C_wl
Rw16_39 word16_39 word15_39 R_wl
Cwl_16_39 word16_39 gnd C_wl
Rw17_39 word17_39 word16_39 R_wl
Cwl_17_39 word17_39 gnd C_wl
Rw18_39 word18_39 word17_39 R_wl
Cwl_18_39 word18_39 gnd C_wl
Rw19_39 word19_39 word18_39 R_wl
Cwl_19_39 word19_39 gnd C_wl
Rw20_39 word20_39 word19_39 R_wl
Cwl_20_39 word20_39 gnd C_wl
Rw21_39 word21_39 word20_39 R_wl
Cwl_21_39 word21_39 gnd C_wl
Rw22_39 word22_39 word21_39 R_wl
Cwl_22_39 word22_39 gnd C_wl
Rw23_39 word23_39 word22_39 R_wl
Cwl_23_39 word23_39 gnd C_wl
Rw24_39 word24_39 word23_39 R_wl
Cwl_24_39 word24_39 gnd C_wl
Rw25_39 word25_39 word24_39 R_wl
Cwl_25_39 word25_39 gnd C_wl
Rw26_39 word26_39 word25_39 R_wl
Cwl_26_39 word26_39 gnd C_wl
Rw27_39 word27_39 word26_39 R_wl
Cwl_27_39 word27_39 gnd C_wl
Rw28_39 word28_39 word27_39 R_wl
Cwl_28_39 word28_39 gnd C_wl
Rw29_39 word29_39 word28_39 R_wl
Cwl_29_39 word29_39 gnd C_wl
Rw30_39 word30_39 word29_39 R_wl
Cwl_30_39 word30_39 gnd C_wl
Rw31_39 word31_39 word30_39 R_wl
Cwl_31_39 word31_39 gnd C_wl
Rw32_39 word32_39 word31_39 R_wl
Cwl_32_39 word32_39 gnd C_wl
Rw33_39 word33_39 word32_39 R_wl
Cwl_33_39 word33_39 gnd C_wl
Rw34_39 word34_39 word33_39 R_wl
Cwl_34_39 word34_39 gnd C_wl
Rw35_39 word35_39 word34_39 R_wl
Cwl_35_39 word35_39 gnd C_wl
Rw36_39 word36_39 word35_39 R_wl
Cwl_36_39 word36_39 gnd C_wl
Rw37_39 word37_39 word36_39 R_wl
Cwl_37_39 word37_39 gnd C_wl
Rw38_39 word38_39 word37_39 R_wl
Cwl_38_39 word38_39 gnd C_wl
Rw39_39 word39_39 word38_39 R_wl
Cwl_39_39 word39_39 gnd C_wl
Rw40_39 word40_39 word39_39 R_wl
Cwl_40_39 word40_39 gnd C_wl
Rw41_39 word41_39 word40_39 R_wl
Cwl_41_39 word41_39 gnd C_wl
Rw42_39 word42_39 word41_39 R_wl
Cwl_42_39 word42_39 gnd C_wl
Rw43_39 word43_39 word42_39 R_wl
Cwl_43_39 word43_39 gnd C_wl
Rw44_39 word44_39 word43_39 R_wl
Cwl_44_39 word44_39 gnd C_wl
Rw45_39 word45_39 word44_39 R_wl
Cwl_45_39 word45_39 gnd C_wl
Rw46_39 word46_39 word45_39 R_wl
Cwl_46_39 word46_39 gnd C_wl
Rw47_39 word47_39 word46_39 R_wl
Cwl_47_39 word47_39 gnd C_wl
Rw48_39 word48_39 word47_39 R_wl
Cwl_48_39 word48_39 gnd C_wl
Rw49_39 word49_39 word48_39 R_wl
Cwl_49_39 word49_39 gnd C_wl
Rw50_39 word50_39 word49_39 R_wl
Cwl_50_39 word50_39 gnd C_wl
Rw51_39 word51_39 word50_39 R_wl
Cwl_51_39 word51_39 gnd C_wl
Rw52_39 word52_39 word51_39 R_wl
Cwl_52_39 word52_39 gnd C_wl
Rw53_39 word53_39 word52_39 R_wl
Cwl_53_39 word53_39 gnd C_wl
Rw54_39 word54_39 word53_39 R_wl
Cwl_54_39 word54_39 gnd C_wl
Rw55_39 word55_39 word54_39 R_wl
Cwl_55_39 word55_39 gnd C_wl
Rw56_39 word56_39 word55_39 R_wl
Cwl_56_39 word56_39 gnd C_wl
Rw57_39 word57_39 word56_39 R_wl
Cwl_57_39 word57_39 gnd C_wl
Rw58_39 word58_39 word57_39 R_wl
Cwl_58_39 word58_39 gnd C_wl
Rw59_39 word59_39 word58_39 R_wl
Cwl_59_39 word59_39 gnd C_wl
Rw60_39 word60_39 word59_39 R_wl
Cwl_60_39 word60_39 gnd C_wl
Rw61_39 word61_39 word60_39 R_wl
Cwl_61_39 word61_39 gnd C_wl
Rw62_39 word62_39 word61_39 R_wl
Cwl_62_39 word62_39 gnd C_wl
Rw63_39 word63_39 word62_39 R_wl
Cwl_63_39 word63_39 gnd C_wl
Rw64_39 word64_39 word63_39 R_wl
Cwl_64_39 word64_39 gnd C_wl
Rw65_39 word65_39 word64_39 R_wl
Cwl_65_39 word65_39 gnd C_wl
Rw66_39 word66_39 word65_39 R_wl
Cwl_66_39 word66_39 gnd C_wl
Rw67_39 word67_39 word66_39 R_wl
Cwl_67_39 word67_39 gnd C_wl
Rw68_39 word68_39 word67_39 R_wl
Cwl_68_39 word68_39 gnd C_wl
Rw69_39 word69_39 word68_39 R_wl
Cwl_69_39 word69_39 gnd C_wl
Rw70_39 word70_39 word69_39 R_wl
Cwl_70_39 word70_39 gnd C_wl
Rw71_39 word71_39 word70_39 R_wl
Cwl_71_39 word71_39 gnd C_wl
Rw72_39 word72_39 word71_39 R_wl
Cwl_72_39 word72_39 gnd C_wl
Rw73_39 word73_39 word72_39 R_wl
Cwl_73_39 word73_39 gnd C_wl
Rw74_39 word74_39 word73_39 R_wl
Cwl_74_39 word74_39 gnd C_wl
Rw75_39 word75_39 word74_39 R_wl
Cwl_75_39 word75_39 gnd C_wl
Rw76_39 word76_39 word75_39 R_wl
Cwl_76_39 word76_39 gnd C_wl
Rw77_39 word77_39 word76_39 R_wl
Cwl_77_39 word77_39 gnd C_wl
Rw78_39 word78_39 word77_39 R_wl
Cwl_78_39 word78_39 gnd C_wl
Rw79_39 word79_39 word78_39 R_wl
Cwl_79_39 word79_39 gnd C_wl
Rw80_39 word80_39 word79_39 R_wl
Cwl_80_39 word80_39 gnd C_wl
Rw81_39 word81_39 word80_39 R_wl
Cwl_81_39 word81_39 gnd C_wl
Rw82_39 word82_39 word81_39 R_wl
Cwl_82_39 word82_39 gnd C_wl
Rw83_39 word83_39 word82_39 R_wl
Cwl_83_39 word83_39 gnd C_wl
Rw84_39 word84_39 word83_39 R_wl
Cwl_84_39 word84_39 gnd C_wl
Rw85_39 word85_39 word84_39 R_wl
Cwl_85_39 word85_39 gnd C_wl
Rw86_39 word86_39 word85_39 R_wl
Cwl_86_39 word86_39 gnd C_wl
Rw87_39 word87_39 word86_39 R_wl
Cwl_87_39 word87_39 gnd C_wl
Rw88_39 word88_39 word87_39 R_wl
Cwl_88_39 word88_39 gnd C_wl
Rw89_39 word89_39 word88_39 R_wl
Cwl_89_39 word89_39 gnd C_wl
Rw90_39 word90_39 word89_39 R_wl
Cwl_90_39 word90_39 gnd C_wl
Rw91_39 word91_39 word90_39 R_wl
Cwl_91_39 word91_39 gnd C_wl
Rw92_39 word92_39 word91_39 R_wl
Cwl_92_39 word92_39 gnd C_wl
Rw93_39 word93_39 word92_39 R_wl
Cwl_93_39 word93_39 gnd C_wl
Rw94_39 word94_39 word93_39 R_wl
Cwl_94_39 word94_39 gnd C_wl
Rw95_39 word95_39 word94_39 R_wl
Cwl_95_39 word95_39 gnd C_wl
Rw96_39 word96_39 word95_39 R_wl
Cwl_96_39 word96_39 gnd C_wl
Rw97_39 word97_39 word96_39 R_wl
Cwl_97_39 word97_39 gnd C_wl
Rw98_39 word98_39 word97_39 R_wl
Cwl_98_39 word98_39 gnd C_wl
Rw99_39 word99_39 word98_39 R_wl
Cwl_99_39 word99_39 gnd C_wl
Vwl_40 word_40 0 0
Rw0_40 word_40 word0_40 R_wl
Cwl_0_40 word0_40 gnd C_wl
Rw1_40 word1_40 word0_40 R_wl
Cwl_1_40 word1_40 gnd C_wl
Rw2_40 word2_40 word1_40 R_wl
Cwl_2_40 word2_40 gnd C_wl
Rw3_40 word3_40 word2_40 R_wl
Cwl_3_40 word3_40 gnd C_wl
Rw4_40 word4_40 word3_40 R_wl
Cwl_4_40 word4_40 gnd C_wl
Rw5_40 word5_40 word4_40 R_wl
Cwl_5_40 word5_40 gnd C_wl
Rw6_40 word6_40 word5_40 R_wl
Cwl_6_40 word6_40 gnd C_wl
Rw7_40 word7_40 word6_40 R_wl
Cwl_7_40 word7_40 gnd C_wl
Rw8_40 word8_40 word7_40 R_wl
Cwl_8_40 word8_40 gnd C_wl
Rw9_40 word9_40 word8_40 R_wl
Cwl_9_40 word9_40 gnd C_wl
Rw10_40 word10_40 word9_40 R_wl
Cwl_10_40 word10_40 gnd C_wl
Rw11_40 word11_40 word10_40 R_wl
Cwl_11_40 word11_40 gnd C_wl
Rw12_40 word12_40 word11_40 R_wl
Cwl_12_40 word12_40 gnd C_wl
Rw13_40 word13_40 word12_40 R_wl
Cwl_13_40 word13_40 gnd C_wl
Rw14_40 word14_40 word13_40 R_wl
Cwl_14_40 word14_40 gnd C_wl
Rw15_40 word15_40 word14_40 R_wl
Cwl_15_40 word15_40 gnd C_wl
Rw16_40 word16_40 word15_40 R_wl
Cwl_16_40 word16_40 gnd C_wl
Rw17_40 word17_40 word16_40 R_wl
Cwl_17_40 word17_40 gnd C_wl
Rw18_40 word18_40 word17_40 R_wl
Cwl_18_40 word18_40 gnd C_wl
Rw19_40 word19_40 word18_40 R_wl
Cwl_19_40 word19_40 gnd C_wl
Rw20_40 word20_40 word19_40 R_wl
Cwl_20_40 word20_40 gnd C_wl
Rw21_40 word21_40 word20_40 R_wl
Cwl_21_40 word21_40 gnd C_wl
Rw22_40 word22_40 word21_40 R_wl
Cwl_22_40 word22_40 gnd C_wl
Rw23_40 word23_40 word22_40 R_wl
Cwl_23_40 word23_40 gnd C_wl
Rw24_40 word24_40 word23_40 R_wl
Cwl_24_40 word24_40 gnd C_wl
Rw25_40 word25_40 word24_40 R_wl
Cwl_25_40 word25_40 gnd C_wl
Rw26_40 word26_40 word25_40 R_wl
Cwl_26_40 word26_40 gnd C_wl
Rw27_40 word27_40 word26_40 R_wl
Cwl_27_40 word27_40 gnd C_wl
Rw28_40 word28_40 word27_40 R_wl
Cwl_28_40 word28_40 gnd C_wl
Rw29_40 word29_40 word28_40 R_wl
Cwl_29_40 word29_40 gnd C_wl
Rw30_40 word30_40 word29_40 R_wl
Cwl_30_40 word30_40 gnd C_wl
Rw31_40 word31_40 word30_40 R_wl
Cwl_31_40 word31_40 gnd C_wl
Rw32_40 word32_40 word31_40 R_wl
Cwl_32_40 word32_40 gnd C_wl
Rw33_40 word33_40 word32_40 R_wl
Cwl_33_40 word33_40 gnd C_wl
Rw34_40 word34_40 word33_40 R_wl
Cwl_34_40 word34_40 gnd C_wl
Rw35_40 word35_40 word34_40 R_wl
Cwl_35_40 word35_40 gnd C_wl
Rw36_40 word36_40 word35_40 R_wl
Cwl_36_40 word36_40 gnd C_wl
Rw37_40 word37_40 word36_40 R_wl
Cwl_37_40 word37_40 gnd C_wl
Rw38_40 word38_40 word37_40 R_wl
Cwl_38_40 word38_40 gnd C_wl
Rw39_40 word39_40 word38_40 R_wl
Cwl_39_40 word39_40 gnd C_wl
Rw40_40 word40_40 word39_40 R_wl
Cwl_40_40 word40_40 gnd C_wl
Rw41_40 word41_40 word40_40 R_wl
Cwl_41_40 word41_40 gnd C_wl
Rw42_40 word42_40 word41_40 R_wl
Cwl_42_40 word42_40 gnd C_wl
Rw43_40 word43_40 word42_40 R_wl
Cwl_43_40 word43_40 gnd C_wl
Rw44_40 word44_40 word43_40 R_wl
Cwl_44_40 word44_40 gnd C_wl
Rw45_40 word45_40 word44_40 R_wl
Cwl_45_40 word45_40 gnd C_wl
Rw46_40 word46_40 word45_40 R_wl
Cwl_46_40 word46_40 gnd C_wl
Rw47_40 word47_40 word46_40 R_wl
Cwl_47_40 word47_40 gnd C_wl
Rw48_40 word48_40 word47_40 R_wl
Cwl_48_40 word48_40 gnd C_wl
Rw49_40 word49_40 word48_40 R_wl
Cwl_49_40 word49_40 gnd C_wl
Rw50_40 word50_40 word49_40 R_wl
Cwl_50_40 word50_40 gnd C_wl
Rw51_40 word51_40 word50_40 R_wl
Cwl_51_40 word51_40 gnd C_wl
Rw52_40 word52_40 word51_40 R_wl
Cwl_52_40 word52_40 gnd C_wl
Rw53_40 word53_40 word52_40 R_wl
Cwl_53_40 word53_40 gnd C_wl
Rw54_40 word54_40 word53_40 R_wl
Cwl_54_40 word54_40 gnd C_wl
Rw55_40 word55_40 word54_40 R_wl
Cwl_55_40 word55_40 gnd C_wl
Rw56_40 word56_40 word55_40 R_wl
Cwl_56_40 word56_40 gnd C_wl
Rw57_40 word57_40 word56_40 R_wl
Cwl_57_40 word57_40 gnd C_wl
Rw58_40 word58_40 word57_40 R_wl
Cwl_58_40 word58_40 gnd C_wl
Rw59_40 word59_40 word58_40 R_wl
Cwl_59_40 word59_40 gnd C_wl
Rw60_40 word60_40 word59_40 R_wl
Cwl_60_40 word60_40 gnd C_wl
Rw61_40 word61_40 word60_40 R_wl
Cwl_61_40 word61_40 gnd C_wl
Rw62_40 word62_40 word61_40 R_wl
Cwl_62_40 word62_40 gnd C_wl
Rw63_40 word63_40 word62_40 R_wl
Cwl_63_40 word63_40 gnd C_wl
Rw64_40 word64_40 word63_40 R_wl
Cwl_64_40 word64_40 gnd C_wl
Rw65_40 word65_40 word64_40 R_wl
Cwl_65_40 word65_40 gnd C_wl
Rw66_40 word66_40 word65_40 R_wl
Cwl_66_40 word66_40 gnd C_wl
Rw67_40 word67_40 word66_40 R_wl
Cwl_67_40 word67_40 gnd C_wl
Rw68_40 word68_40 word67_40 R_wl
Cwl_68_40 word68_40 gnd C_wl
Rw69_40 word69_40 word68_40 R_wl
Cwl_69_40 word69_40 gnd C_wl
Rw70_40 word70_40 word69_40 R_wl
Cwl_70_40 word70_40 gnd C_wl
Rw71_40 word71_40 word70_40 R_wl
Cwl_71_40 word71_40 gnd C_wl
Rw72_40 word72_40 word71_40 R_wl
Cwl_72_40 word72_40 gnd C_wl
Rw73_40 word73_40 word72_40 R_wl
Cwl_73_40 word73_40 gnd C_wl
Rw74_40 word74_40 word73_40 R_wl
Cwl_74_40 word74_40 gnd C_wl
Rw75_40 word75_40 word74_40 R_wl
Cwl_75_40 word75_40 gnd C_wl
Rw76_40 word76_40 word75_40 R_wl
Cwl_76_40 word76_40 gnd C_wl
Rw77_40 word77_40 word76_40 R_wl
Cwl_77_40 word77_40 gnd C_wl
Rw78_40 word78_40 word77_40 R_wl
Cwl_78_40 word78_40 gnd C_wl
Rw79_40 word79_40 word78_40 R_wl
Cwl_79_40 word79_40 gnd C_wl
Rw80_40 word80_40 word79_40 R_wl
Cwl_80_40 word80_40 gnd C_wl
Rw81_40 word81_40 word80_40 R_wl
Cwl_81_40 word81_40 gnd C_wl
Rw82_40 word82_40 word81_40 R_wl
Cwl_82_40 word82_40 gnd C_wl
Rw83_40 word83_40 word82_40 R_wl
Cwl_83_40 word83_40 gnd C_wl
Rw84_40 word84_40 word83_40 R_wl
Cwl_84_40 word84_40 gnd C_wl
Rw85_40 word85_40 word84_40 R_wl
Cwl_85_40 word85_40 gnd C_wl
Rw86_40 word86_40 word85_40 R_wl
Cwl_86_40 word86_40 gnd C_wl
Rw87_40 word87_40 word86_40 R_wl
Cwl_87_40 word87_40 gnd C_wl
Rw88_40 word88_40 word87_40 R_wl
Cwl_88_40 word88_40 gnd C_wl
Rw89_40 word89_40 word88_40 R_wl
Cwl_89_40 word89_40 gnd C_wl
Rw90_40 word90_40 word89_40 R_wl
Cwl_90_40 word90_40 gnd C_wl
Rw91_40 word91_40 word90_40 R_wl
Cwl_91_40 word91_40 gnd C_wl
Rw92_40 word92_40 word91_40 R_wl
Cwl_92_40 word92_40 gnd C_wl
Rw93_40 word93_40 word92_40 R_wl
Cwl_93_40 word93_40 gnd C_wl
Rw94_40 word94_40 word93_40 R_wl
Cwl_94_40 word94_40 gnd C_wl
Rw95_40 word95_40 word94_40 R_wl
Cwl_95_40 word95_40 gnd C_wl
Rw96_40 word96_40 word95_40 R_wl
Cwl_96_40 word96_40 gnd C_wl
Rw97_40 word97_40 word96_40 R_wl
Cwl_97_40 word97_40 gnd C_wl
Rw98_40 word98_40 word97_40 R_wl
Cwl_98_40 word98_40 gnd C_wl
Rw99_40 word99_40 word98_40 R_wl
Cwl_99_40 word99_40 gnd C_wl
Vwl_41 word_41 0 0
Rw0_41 word_41 word0_41 R_wl
Cwl_0_41 word0_41 gnd C_wl
Rw1_41 word1_41 word0_41 R_wl
Cwl_1_41 word1_41 gnd C_wl
Rw2_41 word2_41 word1_41 R_wl
Cwl_2_41 word2_41 gnd C_wl
Rw3_41 word3_41 word2_41 R_wl
Cwl_3_41 word3_41 gnd C_wl
Rw4_41 word4_41 word3_41 R_wl
Cwl_4_41 word4_41 gnd C_wl
Rw5_41 word5_41 word4_41 R_wl
Cwl_5_41 word5_41 gnd C_wl
Rw6_41 word6_41 word5_41 R_wl
Cwl_6_41 word6_41 gnd C_wl
Rw7_41 word7_41 word6_41 R_wl
Cwl_7_41 word7_41 gnd C_wl
Rw8_41 word8_41 word7_41 R_wl
Cwl_8_41 word8_41 gnd C_wl
Rw9_41 word9_41 word8_41 R_wl
Cwl_9_41 word9_41 gnd C_wl
Rw10_41 word10_41 word9_41 R_wl
Cwl_10_41 word10_41 gnd C_wl
Rw11_41 word11_41 word10_41 R_wl
Cwl_11_41 word11_41 gnd C_wl
Rw12_41 word12_41 word11_41 R_wl
Cwl_12_41 word12_41 gnd C_wl
Rw13_41 word13_41 word12_41 R_wl
Cwl_13_41 word13_41 gnd C_wl
Rw14_41 word14_41 word13_41 R_wl
Cwl_14_41 word14_41 gnd C_wl
Rw15_41 word15_41 word14_41 R_wl
Cwl_15_41 word15_41 gnd C_wl
Rw16_41 word16_41 word15_41 R_wl
Cwl_16_41 word16_41 gnd C_wl
Rw17_41 word17_41 word16_41 R_wl
Cwl_17_41 word17_41 gnd C_wl
Rw18_41 word18_41 word17_41 R_wl
Cwl_18_41 word18_41 gnd C_wl
Rw19_41 word19_41 word18_41 R_wl
Cwl_19_41 word19_41 gnd C_wl
Rw20_41 word20_41 word19_41 R_wl
Cwl_20_41 word20_41 gnd C_wl
Rw21_41 word21_41 word20_41 R_wl
Cwl_21_41 word21_41 gnd C_wl
Rw22_41 word22_41 word21_41 R_wl
Cwl_22_41 word22_41 gnd C_wl
Rw23_41 word23_41 word22_41 R_wl
Cwl_23_41 word23_41 gnd C_wl
Rw24_41 word24_41 word23_41 R_wl
Cwl_24_41 word24_41 gnd C_wl
Rw25_41 word25_41 word24_41 R_wl
Cwl_25_41 word25_41 gnd C_wl
Rw26_41 word26_41 word25_41 R_wl
Cwl_26_41 word26_41 gnd C_wl
Rw27_41 word27_41 word26_41 R_wl
Cwl_27_41 word27_41 gnd C_wl
Rw28_41 word28_41 word27_41 R_wl
Cwl_28_41 word28_41 gnd C_wl
Rw29_41 word29_41 word28_41 R_wl
Cwl_29_41 word29_41 gnd C_wl
Rw30_41 word30_41 word29_41 R_wl
Cwl_30_41 word30_41 gnd C_wl
Rw31_41 word31_41 word30_41 R_wl
Cwl_31_41 word31_41 gnd C_wl
Rw32_41 word32_41 word31_41 R_wl
Cwl_32_41 word32_41 gnd C_wl
Rw33_41 word33_41 word32_41 R_wl
Cwl_33_41 word33_41 gnd C_wl
Rw34_41 word34_41 word33_41 R_wl
Cwl_34_41 word34_41 gnd C_wl
Rw35_41 word35_41 word34_41 R_wl
Cwl_35_41 word35_41 gnd C_wl
Rw36_41 word36_41 word35_41 R_wl
Cwl_36_41 word36_41 gnd C_wl
Rw37_41 word37_41 word36_41 R_wl
Cwl_37_41 word37_41 gnd C_wl
Rw38_41 word38_41 word37_41 R_wl
Cwl_38_41 word38_41 gnd C_wl
Rw39_41 word39_41 word38_41 R_wl
Cwl_39_41 word39_41 gnd C_wl
Rw40_41 word40_41 word39_41 R_wl
Cwl_40_41 word40_41 gnd C_wl
Rw41_41 word41_41 word40_41 R_wl
Cwl_41_41 word41_41 gnd C_wl
Rw42_41 word42_41 word41_41 R_wl
Cwl_42_41 word42_41 gnd C_wl
Rw43_41 word43_41 word42_41 R_wl
Cwl_43_41 word43_41 gnd C_wl
Rw44_41 word44_41 word43_41 R_wl
Cwl_44_41 word44_41 gnd C_wl
Rw45_41 word45_41 word44_41 R_wl
Cwl_45_41 word45_41 gnd C_wl
Rw46_41 word46_41 word45_41 R_wl
Cwl_46_41 word46_41 gnd C_wl
Rw47_41 word47_41 word46_41 R_wl
Cwl_47_41 word47_41 gnd C_wl
Rw48_41 word48_41 word47_41 R_wl
Cwl_48_41 word48_41 gnd C_wl
Rw49_41 word49_41 word48_41 R_wl
Cwl_49_41 word49_41 gnd C_wl
Rw50_41 word50_41 word49_41 R_wl
Cwl_50_41 word50_41 gnd C_wl
Rw51_41 word51_41 word50_41 R_wl
Cwl_51_41 word51_41 gnd C_wl
Rw52_41 word52_41 word51_41 R_wl
Cwl_52_41 word52_41 gnd C_wl
Rw53_41 word53_41 word52_41 R_wl
Cwl_53_41 word53_41 gnd C_wl
Rw54_41 word54_41 word53_41 R_wl
Cwl_54_41 word54_41 gnd C_wl
Rw55_41 word55_41 word54_41 R_wl
Cwl_55_41 word55_41 gnd C_wl
Rw56_41 word56_41 word55_41 R_wl
Cwl_56_41 word56_41 gnd C_wl
Rw57_41 word57_41 word56_41 R_wl
Cwl_57_41 word57_41 gnd C_wl
Rw58_41 word58_41 word57_41 R_wl
Cwl_58_41 word58_41 gnd C_wl
Rw59_41 word59_41 word58_41 R_wl
Cwl_59_41 word59_41 gnd C_wl
Rw60_41 word60_41 word59_41 R_wl
Cwl_60_41 word60_41 gnd C_wl
Rw61_41 word61_41 word60_41 R_wl
Cwl_61_41 word61_41 gnd C_wl
Rw62_41 word62_41 word61_41 R_wl
Cwl_62_41 word62_41 gnd C_wl
Rw63_41 word63_41 word62_41 R_wl
Cwl_63_41 word63_41 gnd C_wl
Rw64_41 word64_41 word63_41 R_wl
Cwl_64_41 word64_41 gnd C_wl
Rw65_41 word65_41 word64_41 R_wl
Cwl_65_41 word65_41 gnd C_wl
Rw66_41 word66_41 word65_41 R_wl
Cwl_66_41 word66_41 gnd C_wl
Rw67_41 word67_41 word66_41 R_wl
Cwl_67_41 word67_41 gnd C_wl
Rw68_41 word68_41 word67_41 R_wl
Cwl_68_41 word68_41 gnd C_wl
Rw69_41 word69_41 word68_41 R_wl
Cwl_69_41 word69_41 gnd C_wl
Rw70_41 word70_41 word69_41 R_wl
Cwl_70_41 word70_41 gnd C_wl
Rw71_41 word71_41 word70_41 R_wl
Cwl_71_41 word71_41 gnd C_wl
Rw72_41 word72_41 word71_41 R_wl
Cwl_72_41 word72_41 gnd C_wl
Rw73_41 word73_41 word72_41 R_wl
Cwl_73_41 word73_41 gnd C_wl
Rw74_41 word74_41 word73_41 R_wl
Cwl_74_41 word74_41 gnd C_wl
Rw75_41 word75_41 word74_41 R_wl
Cwl_75_41 word75_41 gnd C_wl
Rw76_41 word76_41 word75_41 R_wl
Cwl_76_41 word76_41 gnd C_wl
Rw77_41 word77_41 word76_41 R_wl
Cwl_77_41 word77_41 gnd C_wl
Rw78_41 word78_41 word77_41 R_wl
Cwl_78_41 word78_41 gnd C_wl
Rw79_41 word79_41 word78_41 R_wl
Cwl_79_41 word79_41 gnd C_wl
Rw80_41 word80_41 word79_41 R_wl
Cwl_80_41 word80_41 gnd C_wl
Rw81_41 word81_41 word80_41 R_wl
Cwl_81_41 word81_41 gnd C_wl
Rw82_41 word82_41 word81_41 R_wl
Cwl_82_41 word82_41 gnd C_wl
Rw83_41 word83_41 word82_41 R_wl
Cwl_83_41 word83_41 gnd C_wl
Rw84_41 word84_41 word83_41 R_wl
Cwl_84_41 word84_41 gnd C_wl
Rw85_41 word85_41 word84_41 R_wl
Cwl_85_41 word85_41 gnd C_wl
Rw86_41 word86_41 word85_41 R_wl
Cwl_86_41 word86_41 gnd C_wl
Rw87_41 word87_41 word86_41 R_wl
Cwl_87_41 word87_41 gnd C_wl
Rw88_41 word88_41 word87_41 R_wl
Cwl_88_41 word88_41 gnd C_wl
Rw89_41 word89_41 word88_41 R_wl
Cwl_89_41 word89_41 gnd C_wl
Rw90_41 word90_41 word89_41 R_wl
Cwl_90_41 word90_41 gnd C_wl
Rw91_41 word91_41 word90_41 R_wl
Cwl_91_41 word91_41 gnd C_wl
Rw92_41 word92_41 word91_41 R_wl
Cwl_92_41 word92_41 gnd C_wl
Rw93_41 word93_41 word92_41 R_wl
Cwl_93_41 word93_41 gnd C_wl
Rw94_41 word94_41 word93_41 R_wl
Cwl_94_41 word94_41 gnd C_wl
Rw95_41 word95_41 word94_41 R_wl
Cwl_95_41 word95_41 gnd C_wl
Rw96_41 word96_41 word95_41 R_wl
Cwl_96_41 word96_41 gnd C_wl
Rw97_41 word97_41 word96_41 R_wl
Cwl_97_41 word97_41 gnd C_wl
Rw98_41 word98_41 word97_41 R_wl
Cwl_98_41 word98_41 gnd C_wl
Rw99_41 word99_41 word98_41 R_wl
Cwl_99_41 word99_41 gnd C_wl
Vwl_42 word_42 0 0
Rw0_42 word_42 word0_42 R_wl
Cwl_0_42 word0_42 gnd C_wl
Rw1_42 word1_42 word0_42 R_wl
Cwl_1_42 word1_42 gnd C_wl
Rw2_42 word2_42 word1_42 R_wl
Cwl_2_42 word2_42 gnd C_wl
Rw3_42 word3_42 word2_42 R_wl
Cwl_3_42 word3_42 gnd C_wl
Rw4_42 word4_42 word3_42 R_wl
Cwl_4_42 word4_42 gnd C_wl
Rw5_42 word5_42 word4_42 R_wl
Cwl_5_42 word5_42 gnd C_wl
Rw6_42 word6_42 word5_42 R_wl
Cwl_6_42 word6_42 gnd C_wl
Rw7_42 word7_42 word6_42 R_wl
Cwl_7_42 word7_42 gnd C_wl
Rw8_42 word8_42 word7_42 R_wl
Cwl_8_42 word8_42 gnd C_wl
Rw9_42 word9_42 word8_42 R_wl
Cwl_9_42 word9_42 gnd C_wl
Rw10_42 word10_42 word9_42 R_wl
Cwl_10_42 word10_42 gnd C_wl
Rw11_42 word11_42 word10_42 R_wl
Cwl_11_42 word11_42 gnd C_wl
Rw12_42 word12_42 word11_42 R_wl
Cwl_12_42 word12_42 gnd C_wl
Rw13_42 word13_42 word12_42 R_wl
Cwl_13_42 word13_42 gnd C_wl
Rw14_42 word14_42 word13_42 R_wl
Cwl_14_42 word14_42 gnd C_wl
Rw15_42 word15_42 word14_42 R_wl
Cwl_15_42 word15_42 gnd C_wl
Rw16_42 word16_42 word15_42 R_wl
Cwl_16_42 word16_42 gnd C_wl
Rw17_42 word17_42 word16_42 R_wl
Cwl_17_42 word17_42 gnd C_wl
Rw18_42 word18_42 word17_42 R_wl
Cwl_18_42 word18_42 gnd C_wl
Rw19_42 word19_42 word18_42 R_wl
Cwl_19_42 word19_42 gnd C_wl
Rw20_42 word20_42 word19_42 R_wl
Cwl_20_42 word20_42 gnd C_wl
Rw21_42 word21_42 word20_42 R_wl
Cwl_21_42 word21_42 gnd C_wl
Rw22_42 word22_42 word21_42 R_wl
Cwl_22_42 word22_42 gnd C_wl
Rw23_42 word23_42 word22_42 R_wl
Cwl_23_42 word23_42 gnd C_wl
Rw24_42 word24_42 word23_42 R_wl
Cwl_24_42 word24_42 gnd C_wl
Rw25_42 word25_42 word24_42 R_wl
Cwl_25_42 word25_42 gnd C_wl
Rw26_42 word26_42 word25_42 R_wl
Cwl_26_42 word26_42 gnd C_wl
Rw27_42 word27_42 word26_42 R_wl
Cwl_27_42 word27_42 gnd C_wl
Rw28_42 word28_42 word27_42 R_wl
Cwl_28_42 word28_42 gnd C_wl
Rw29_42 word29_42 word28_42 R_wl
Cwl_29_42 word29_42 gnd C_wl
Rw30_42 word30_42 word29_42 R_wl
Cwl_30_42 word30_42 gnd C_wl
Rw31_42 word31_42 word30_42 R_wl
Cwl_31_42 word31_42 gnd C_wl
Rw32_42 word32_42 word31_42 R_wl
Cwl_32_42 word32_42 gnd C_wl
Rw33_42 word33_42 word32_42 R_wl
Cwl_33_42 word33_42 gnd C_wl
Rw34_42 word34_42 word33_42 R_wl
Cwl_34_42 word34_42 gnd C_wl
Rw35_42 word35_42 word34_42 R_wl
Cwl_35_42 word35_42 gnd C_wl
Rw36_42 word36_42 word35_42 R_wl
Cwl_36_42 word36_42 gnd C_wl
Rw37_42 word37_42 word36_42 R_wl
Cwl_37_42 word37_42 gnd C_wl
Rw38_42 word38_42 word37_42 R_wl
Cwl_38_42 word38_42 gnd C_wl
Rw39_42 word39_42 word38_42 R_wl
Cwl_39_42 word39_42 gnd C_wl
Rw40_42 word40_42 word39_42 R_wl
Cwl_40_42 word40_42 gnd C_wl
Rw41_42 word41_42 word40_42 R_wl
Cwl_41_42 word41_42 gnd C_wl
Rw42_42 word42_42 word41_42 R_wl
Cwl_42_42 word42_42 gnd C_wl
Rw43_42 word43_42 word42_42 R_wl
Cwl_43_42 word43_42 gnd C_wl
Rw44_42 word44_42 word43_42 R_wl
Cwl_44_42 word44_42 gnd C_wl
Rw45_42 word45_42 word44_42 R_wl
Cwl_45_42 word45_42 gnd C_wl
Rw46_42 word46_42 word45_42 R_wl
Cwl_46_42 word46_42 gnd C_wl
Rw47_42 word47_42 word46_42 R_wl
Cwl_47_42 word47_42 gnd C_wl
Rw48_42 word48_42 word47_42 R_wl
Cwl_48_42 word48_42 gnd C_wl
Rw49_42 word49_42 word48_42 R_wl
Cwl_49_42 word49_42 gnd C_wl
Rw50_42 word50_42 word49_42 R_wl
Cwl_50_42 word50_42 gnd C_wl
Rw51_42 word51_42 word50_42 R_wl
Cwl_51_42 word51_42 gnd C_wl
Rw52_42 word52_42 word51_42 R_wl
Cwl_52_42 word52_42 gnd C_wl
Rw53_42 word53_42 word52_42 R_wl
Cwl_53_42 word53_42 gnd C_wl
Rw54_42 word54_42 word53_42 R_wl
Cwl_54_42 word54_42 gnd C_wl
Rw55_42 word55_42 word54_42 R_wl
Cwl_55_42 word55_42 gnd C_wl
Rw56_42 word56_42 word55_42 R_wl
Cwl_56_42 word56_42 gnd C_wl
Rw57_42 word57_42 word56_42 R_wl
Cwl_57_42 word57_42 gnd C_wl
Rw58_42 word58_42 word57_42 R_wl
Cwl_58_42 word58_42 gnd C_wl
Rw59_42 word59_42 word58_42 R_wl
Cwl_59_42 word59_42 gnd C_wl
Rw60_42 word60_42 word59_42 R_wl
Cwl_60_42 word60_42 gnd C_wl
Rw61_42 word61_42 word60_42 R_wl
Cwl_61_42 word61_42 gnd C_wl
Rw62_42 word62_42 word61_42 R_wl
Cwl_62_42 word62_42 gnd C_wl
Rw63_42 word63_42 word62_42 R_wl
Cwl_63_42 word63_42 gnd C_wl
Rw64_42 word64_42 word63_42 R_wl
Cwl_64_42 word64_42 gnd C_wl
Rw65_42 word65_42 word64_42 R_wl
Cwl_65_42 word65_42 gnd C_wl
Rw66_42 word66_42 word65_42 R_wl
Cwl_66_42 word66_42 gnd C_wl
Rw67_42 word67_42 word66_42 R_wl
Cwl_67_42 word67_42 gnd C_wl
Rw68_42 word68_42 word67_42 R_wl
Cwl_68_42 word68_42 gnd C_wl
Rw69_42 word69_42 word68_42 R_wl
Cwl_69_42 word69_42 gnd C_wl
Rw70_42 word70_42 word69_42 R_wl
Cwl_70_42 word70_42 gnd C_wl
Rw71_42 word71_42 word70_42 R_wl
Cwl_71_42 word71_42 gnd C_wl
Rw72_42 word72_42 word71_42 R_wl
Cwl_72_42 word72_42 gnd C_wl
Rw73_42 word73_42 word72_42 R_wl
Cwl_73_42 word73_42 gnd C_wl
Rw74_42 word74_42 word73_42 R_wl
Cwl_74_42 word74_42 gnd C_wl
Rw75_42 word75_42 word74_42 R_wl
Cwl_75_42 word75_42 gnd C_wl
Rw76_42 word76_42 word75_42 R_wl
Cwl_76_42 word76_42 gnd C_wl
Rw77_42 word77_42 word76_42 R_wl
Cwl_77_42 word77_42 gnd C_wl
Rw78_42 word78_42 word77_42 R_wl
Cwl_78_42 word78_42 gnd C_wl
Rw79_42 word79_42 word78_42 R_wl
Cwl_79_42 word79_42 gnd C_wl
Rw80_42 word80_42 word79_42 R_wl
Cwl_80_42 word80_42 gnd C_wl
Rw81_42 word81_42 word80_42 R_wl
Cwl_81_42 word81_42 gnd C_wl
Rw82_42 word82_42 word81_42 R_wl
Cwl_82_42 word82_42 gnd C_wl
Rw83_42 word83_42 word82_42 R_wl
Cwl_83_42 word83_42 gnd C_wl
Rw84_42 word84_42 word83_42 R_wl
Cwl_84_42 word84_42 gnd C_wl
Rw85_42 word85_42 word84_42 R_wl
Cwl_85_42 word85_42 gnd C_wl
Rw86_42 word86_42 word85_42 R_wl
Cwl_86_42 word86_42 gnd C_wl
Rw87_42 word87_42 word86_42 R_wl
Cwl_87_42 word87_42 gnd C_wl
Rw88_42 word88_42 word87_42 R_wl
Cwl_88_42 word88_42 gnd C_wl
Rw89_42 word89_42 word88_42 R_wl
Cwl_89_42 word89_42 gnd C_wl
Rw90_42 word90_42 word89_42 R_wl
Cwl_90_42 word90_42 gnd C_wl
Rw91_42 word91_42 word90_42 R_wl
Cwl_91_42 word91_42 gnd C_wl
Rw92_42 word92_42 word91_42 R_wl
Cwl_92_42 word92_42 gnd C_wl
Rw93_42 word93_42 word92_42 R_wl
Cwl_93_42 word93_42 gnd C_wl
Rw94_42 word94_42 word93_42 R_wl
Cwl_94_42 word94_42 gnd C_wl
Rw95_42 word95_42 word94_42 R_wl
Cwl_95_42 word95_42 gnd C_wl
Rw96_42 word96_42 word95_42 R_wl
Cwl_96_42 word96_42 gnd C_wl
Rw97_42 word97_42 word96_42 R_wl
Cwl_97_42 word97_42 gnd C_wl
Rw98_42 word98_42 word97_42 R_wl
Cwl_98_42 word98_42 gnd C_wl
Rw99_42 word99_42 word98_42 R_wl
Cwl_99_42 word99_42 gnd C_wl
Vwl_43 word_43 0 0
Rw0_43 word_43 word0_43 R_wl
Cwl_0_43 word0_43 gnd C_wl
Rw1_43 word1_43 word0_43 R_wl
Cwl_1_43 word1_43 gnd C_wl
Rw2_43 word2_43 word1_43 R_wl
Cwl_2_43 word2_43 gnd C_wl
Rw3_43 word3_43 word2_43 R_wl
Cwl_3_43 word3_43 gnd C_wl
Rw4_43 word4_43 word3_43 R_wl
Cwl_4_43 word4_43 gnd C_wl
Rw5_43 word5_43 word4_43 R_wl
Cwl_5_43 word5_43 gnd C_wl
Rw6_43 word6_43 word5_43 R_wl
Cwl_6_43 word6_43 gnd C_wl
Rw7_43 word7_43 word6_43 R_wl
Cwl_7_43 word7_43 gnd C_wl
Rw8_43 word8_43 word7_43 R_wl
Cwl_8_43 word8_43 gnd C_wl
Rw9_43 word9_43 word8_43 R_wl
Cwl_9_43 word9_43 gnd C_wl
Rw10_43 word10_43 word9_43 R_wl
Cwl_10_43 word10_43 gnd C_wl
Rw11_43 word11_43 word10_43 R_wl
Cwl_11_43 word11_43 gnd C_wl
Rw12_43 word12_43 word11_43 R_wl
Cwl_12_43 word12_43 gnd C_wl
Rw13_43 word13_43 word12_43 R_wl
Cwl_13_43 word13_43 gnd C_wl
Rw14_43 word14_43 word13_43 R_wl
Cwl_14_43 word14_43 gnd C_wl
Rw15_43 word15_43 word14_43 R_wl
Cwl_15_43 word15_43 gnd C_wl
Rw16_43 word16_43 word15_43 R_wl
Cwl_16_43 word16_43 gnd C_wl
Rw17_43 word17_43 word16_43 R_wl
Cwl_17_43 word17_43 gnd C_wl
Rw18_43 word18_43 word17_43 R_wl
Cwl_18_43 word18_43 gnd C_wl
Rw19_43 word19_43 word18_43 R_wl
Cwl_19_43 word19_43 gnd C_wl
Rw20_43 word20_43 word19_43 R_wl
Cwl_20_43 word20_43 gnd C_wl
Rw21_43 word21_43 word20_43 R_wl
Cwl_21_43 word21_43 gnd C_wl
Rw22_43 word22_43 word21_43 R_wl
Cwl_22_43 word22_43 gnd C_wl
Rw23_43 word23_43 word22_43 R_wl
Cwl_23_43 word23_43 gnd C_wl
Rw24_43 word24_43 word23_43 R_wl
Cwl_24_43 word24_43 gnd C_wl
Rw25_43 word25_43 word24_43 R_wl
Cwl_25_43 word25_43 gnd C_wl
Rw26_43 word26_43 word25_43 R_wl
Cwl_26_43 word26_43 gnd C_wl
Rw27_43 word27_43 word26_43 R_wl
Cwl_27_43 word27_43 gnd C_wl
Rw28_43 word28_43 word27_43 R_wl
Cwl_28_43 word28_43 gnd C_wl
Rw29_43 word29_43 word28_43 R_wl
Cwl_29_43 word29_43 gnd C_wl
Rw30_43 word30_43 word29_43 R_wl
Cwl_30_43 word30_43 gnd C_wl
Rw31_43 word31_43 word30_43 R_wl
Cwl_31_43 word31_43 gnd C_wl
Rw32_43 word32_43 word31_43 R_wl
Cwl_32_43 word32_43 gnd C_wl
Rw33_43 word33_43 word32_43 R_wl
Cwl_33_43 word33_43 gnd C_wl
Rw34_43 word34_43 word33_43 R_wl
Cwl_34_43 word34_43 gnd C_wl
Rw35_43 word35_43 word34_43 R_wl
Cwl_35_43 word35_43 gnd C_wl
Rw36_43 word36_43 word35_43 R_wl
Cwl_36_43 word36_43 gnd C_wl
Rw37_43 word37_43 word36_43 R_wl
Cwl_37_43 word37_43 gnd C_wl
Rw38_43 word38_43 word37_43 R_wl
Cwl_38_43 word38_43 gnd C_wl
Rw39_43 word39_43 word38_43 R_wl
Cwl_39_43 word39_43 gnd C_wl
Rw40_43 word40_43 word39_43 R_wl
Cwl_40_43 word40_43 gnd C_wl
Rw41_43 word41_43 word40_43 R_wl
Cwl_41_43 word41_43 gnd C_wl
Rw42_43 word42_43 word41_43 R_wl
Cwl_42_43 word42_43 gnd C_wl
Rw43_43 word43_43 word42_43 R_wl
Cwl_43_43 word43_43 gnd C_wl
Rw44_43 word44_43 word43_43 R_wl
Cwl_44_43 word44_43 gnd C_wl
Rw45_43 word45_43 word44_43 R_wl
Cwl_45_43 word45_43 gnd C_wl
Rw46_43 word46_43 word45_43 R_wl
Cwl_46_43 word46_43 gnd C_wl
Rw47_43 word47_43 word46_43 R_wl
Cwl_47_43 word47_43 gnd C_wl
Rw48_43 word48_43 word47_43 R_wl
Cwl_48_43 word48_43 gnd C_wl
Rw49_43 word49_43 word48_43 R_wl
Cwl_49_43 word49_43 gnd C_wl
Rw50_43 word50_43 word49_43 R_wl
Cwl_50_43 word50_43 gnd C_wl
Rw51_43 word51_43 word50_43 R_wl
Cwl_51_43 word51_43 gnd C_wl
Rw52_43 word52_43 word51_43 R_wl
Cwl_52_43 word52_43 gnd C_wl
Rw53_43 word53_43 word52_43 R_wl
Cwl_53_43 word53_43 gnd C_wl
Rw54_43 word54_43 word53_43 R_wl
Cwl_54_43 word54_43 gnd C_wl
Rw55_43 word55_43 word54_43 R_wl
Cwl_55_43 word55_43 gnd C_wl
Rw56_43 word56_43 word55_43 R_wl
Cwl_56_43 word56_43 gnd C_wl
Rw57_43 word57_43 word56_43 R_wl
Cwl_57_43 word57_43 gnd C_wl
Rw58_43 word58_43 word57_43 R_wl
Cwl_58_43 word58_43 gnd C_wl
Rw59_43 word59_43 word58_43 R_wl
Cwl_59_43 word59_43 gnd C_wl
Rw60_43 word60_43 word59_43 R_wl
Cwl_60_43 word60_43 gnd C_wl
Rw61_43 word61_43 word60_43 R_wl
Cwl_61_43 word61_43 gnd C_wl
Rw62_43 word62_43 word61_43 R_wl
Cwl_62_43 word62_43 gnd C_wl
Rw63_43 word63_43 word62_43 R_wl
Cwl_63_43 word63_43 gnd C_wl
Rw64_43 word64_43 word63_43 R_wl
Cwl_64_43 word64_43 gnd C_wl
Rw65_43 word65_43 word64_43 R_wl
Cwl_65_43 word65_43 gnd C_wl
Rw66_43 word66_43 word65_43 R_wl
Cwl_66_43 word66_43 gnd C_wl
Rw67_43 word67_43 word66_43 R_wl
Cwl_67_43 word67_43 gnd C_wl
Rw68_43 word68_43 word67_43 R_wl
Cwl_68_43 word68_43 gnd C_wl
Rw69_43 word69_43 word68_43 R_wl
Cwl_69_43 word69_43 gnd C_wl
Rw70_43 word70_43 word69_43 R_wl
Cwl_70_43 word70_43 gnd C_wl
Rw71_43 word71_43 word70_43 R_wl
Cwl_71_43 word71_43 gnd C_wl
Rw72_43 word72_43 word71_43 R_wl
Cwl_72_43 word72_43 gnd C_wl
Rw73_43 word73_43 word72_43 R_wl
Cwl_73_43 word73_43 gnd C_wl
Rw74_43 word74_43 word73_43 R_wl
Cwl_74_43 word74_43 gnd C_wl
Rw75_43 word75_43 word74_43 R_wl
Cwl_75_43 word75_43 gnd C_wl
Rw76_43 word76_43 word75_43 R_wl
Cwl_76_43 word76_43 gnd C_wl
Rw77_43 word77_43 word76_43 R_wl
Cwl_77_43 word77_43 gnd C_wl
Rw78_43 word78_43 word77_43 R_wl
Cwl_78_43 word78_43 gnd C_wl
Rw79_43 word79_43 word78_43 R_wl
Cwl_79_43 word79_43 gnd C_wl
Rw80_43 word80_43 word79_43 R_wl
Cwl_80_43 word80_43 gnd C_wl
Rw81_43 word81_43 word80_43 R_wl
Cwl_81_43 word81_43 gnd C_wl
Rw82_43 word82_43 word81_43 R_wl
Cwl_82_43 word82_43 gnd C_wl
Rw83_43 word83_43 word82_43 R_wl
Cwl_83_43 word83_43 gnd C_wl
Rw84_43 word84_43 word83_43 R_wl
Cwl_84_43 word84_43 gnd C_wl
Rw85_43 word85_43 word84_43 R_wl
Cwl_85_43 word85_43 gnd C_wl
Rw86_43 word86_43 word85_43 R_wl
Cwl_86_43 word86_43 gnd C_wl
Rw87_43 word87_43 word86_43 R_wl
Cwl_87_43 word87_43 gnd C_wl
Rw88_43 word88_43 word87_43 R_wl
Cwl_88_43 word88_43 gnd C_wl
Rw89_43 word89_43 word88_43 R_wl
Cwl_89_43 word89_43 gnd C_wl
Rw90_43 word90_43 word89_43 R_wl
Cwl_90_43 word90_43 gnd C_wl
Rw91_43 word91_43 word90_43 R_wl
Cwl_91_43 word91_43 gnd C_wl
Rw92_43 word92_43 word91_43 R_wl
Cwl_92_43 word92_43 gnd C_wl
Rw93_43 word93_43 word92_43 R_wl
Cwl_93_43 word93_43 gnd C_wl
Rw94_43 word94_43 word93_43 R_wl
Cwl_94_43 word94_43 gnd C_wl
Rw95_43 word95_43 word94_43 R_wl
Cwl_95_43 word95_43 gnd C_wl
Rw96_43 word96_43 word95_43 R_wl
Cwl_96_43 word96_43 gnd C_wl
Rw97_43 word97_43 word96_43 R_wl
Cwl_97_43 word97_43 gnd C_wl
Rw98_43 word98_43 word97_43 R_wl
Cwl_98_43 word98_43 gnd C_wl
Rw99_43 word99_43 word98_43 R_wl
Cwl_99_43 word99_43 gnd C_wl
Vwl_44 word_44 0 0
Rw0_44 word_44 word0_44 R_wl
Cwl_0_44 word0_44 gnd C_wl
Rw1_44 word1_44 word0_44 R_wl
Cwl_1_44 word1_44 gnd C_wl
Rw2_44 word2_44 word1_44 R_wl
Cwl_2_44 word2_44 gnd C_wl
Rw3_44 word3_44 word2_44 R_wl
Cwl_3_44 word3_44 gnd C_wl
Rw4_44 word4_44 word3_44 R_wl
Cwl_4_44 word4_44 gnd C_wl
Rw5_44 word5_44 word4_44 R_wl
Cwl_5_44 word5_44 gnd C_wl
Rw6_44 word6_44 word5_44 R_wl
Cwl_6_44 word6_44 gnd C_wl
Rw7_44 word7_44 word6_44 R_wl
Cwl_7_44 word7_44 gnd C_wl
Rw8_44 word8_44 word7_44 R_wl
Cwl_8_44 word8_44 gnd C_wl
Rw9_44 word9_44 word8_44 R_wl
Cwl_9_44 word9_44 gnd C_wl
Rw10_44 word10_44 word9_44 R_wl
Cwl_10_44 word10_44 gnd C_wl
Rw11_44 word11_44 word10_44 R_wl
Cwl_11_44 word11_44 gnd C_wl
Rw12_44 word12_44 word11_44 R_wl
Cwl_12_44 word12_44 gnd C_wl
Rw13_44 word13_44 word12_44 R_wl
Cwl_13_44 word13_44 gnd C_wl
Rw14_44 word14_44 word13_44 R_wl
Cwl_14_44 word14_44 gnd C_wl
Rw15_44 word15_44 word14_44 R_wl
Cwl_15_44 word15_44 gnd C_wl
Rw16_44 word16_44 word15_44 R_wl
Cwl_16_44 word16_44 gnd C_wl
Rw17_44 word17_44 word16_44 R_wl
Cwl_17_44 word17_44 gnd C_wl
Rw18_44 word18_44 word17_44 R_wl
Cwl_18_44 word18_44 gnd C_wl
Rw19_44 word19_44 word18_44 R_wl
Cwl_19_44 word19_44 gnd C_wl
Rw20_44 word20_44 word19_44 R_wl
Cwl_20_44 word20_44 gnd C_wl
Rw21_44 word21_44 word20_44 R_wl
Cwl_21_44 word21_44 gnd C_wl
Rw22_44 word22_44 word21_44 R_wl
Cwl_22_44 word22_44 gnd C_wl
Rw23_44 word23_44 word22_44 R_wl
Cwl_23_44 word23_44 gnd C_wl
Rw24_44 word24_44 word23_44 R_wl
Cwl_24_44 word24_44 gnd C_wl
Rw25_44 word25_44 word24_44 R_wl
Cwl_25_44 word25_44 gnd C_wl
Rw26_44 word26_44 word25_44 R_wl
Cwl_26_44 word26_44 gnd C_wl
Rw27_44 word27_44 word26_44 R_wl
Cwl_27_44 word27_44 gnd C_wl
Rw28_44 word28_44 word27_44 R_wl
Cwl_28_44 word28_44 gnd C_wl
Rw29_44 word29_44 word28_44 R_wl
Cwl_29_44 word29_44 gnd C_wl
Rw30_44 word30_44 word29_44 R_wl
Cwl_30_44 word30_44 gnd C_wl
Rw31_44 word31_44 word30_44 R_wl
Cwl_31_44 word31_44 gnd C_wl
Rw32_44 word32_44 word31_44 R_wl
Cwl_32_44 word32_44 gnd C_wl
Rw33_44 word33_44 word32_44 R_wl
Cwl_33_44 word33_44 gnd C_wl
Rw34_44 word34_44 word33_44 R_wl
Cwl_34_44 word34_44 gnd C_wl
Rw35_44 word35_44 word34_44 R_wl
Cwl_35_44 word35_44 gnd C_wl
Rw36_44 word36_44 word35_44 R_wl
Cwl_36_44 word36_44 gnd C_wl
Rw37_44 word37_44 word36_44 R_wl
Cwl_37_44 word37_44 gnd C_wl
Rw38_44 word38_44 word37_44 R_wl
Cwl_38_44 word38_44 gnd C_wl
Rw39_44 word39_44 word38_44 R_wl
Cwl_39_44 word39_44 gnd C_wl
Rw40_44 word40_44 word39_44 R_wl
Cwl_40_44 word40_44 gnd C_wl
Rw41_44 word41_44 word40_44 R_wl
Cwl_41_44 word41_44 gnd C_wl
Rw42_44 word42_44 word41_44 R_wl
Cwl_42_44 word42_44 gnd C_wl
Rw43_44 word43_44 word42_44 R_wl
Cwl_43_44 word43_44 gnd C_wl
Rw44_44 word44_44 word43_44 R_wl
Cwl_44_44 word44_44 gnd C_wl
Rw45_44 word45_44 word44_44 R_wl
Cwl_45_44 word45_44 gnd C_wl
Rw46_44 word46_44 word45_44 R_wl
Cwl_46_44 word46_44 gnd C_wl
Rw47_44 word47_44 word46_44 R_wl
Cwl_47_44 word47_44 gnd C_wl
Rw48_44 word48_44 word47_44 R_wl
Cwl_48_44 word48_44 gnd C_wl
Rw49_44 word49_44 word48_44 R_wl
Cwl_49_44 word49_44 gnd C_wl
Rw50_44 word50_44 word49_44 R_wl
Cwl_50_44 word50_44 gnd C_wl
Rw51_44 word51_44 word50_44 R_wl
Cwl_51_44 word51_44 gnd C_wl
Rw52_44 word52_44 word51_44 R_wl
Cwl_52_44 word52_44 gnd C_wl
Rw53_44 word53_44 word52_44 R_wl
Cwl_53_44 word53_44 gnd C_wl
Rw54_44 word54_44 word53_44 R_wl
Cwl_54_44 word54_44 gnd C_wl
Rw55_44 word55_44 word54_44 R_wl
Cwl_55_44 word55_44 gnd C_wl
Rw56_44 word56_44 word55_44 R_wl
Cwl_56_44 word56_44 gnd C_wl
Rw57_44 word57_44 word56_44 R_wl
Cwl_57_44 word57_44 gnd C_wl
Rw58_44 word58_44 word57_44 R_wl
Cwl_58_44 word58_44 gnd C_wl
Rw59_44 word59_44 word58_44 R_wl
Cwl_59_44 word59_44 gnd C_wl
Rw60_44 word60_44 word59_44 R_wl
Cwl_60_44 word60_44 gnd C_wl
Rw61_44 word61_44 word60_44 R_wl
Cwl_61_44 word61_44 gnd C_wl
Rw62_44 word62_44 word61_44 R_wl
Cwl_62_44 word62_44 gnd C_wl
Rw63_44 word63_44 word62_44 R_wl
Cwl_63_44 word63_44 gnd C_wl
Rw64_44 word64_44 word63_44 R_wl
Cwl_64_44 word64_44 gnd C_wl
Rw65_44 word65_44 word64_44 R_wl
Cwl_65_44 word65_44 gnd C_wl
Rw66_44 word66_44 word65_44 R_wl
Cwl_66_44 word66_44 gnd C_wl
Rw67_44 word67_44 word66_44 R_wl
Cwl_67_44 word67_44 gnd C_wl
Rw68_44 word68_44 word67_44 R_wl
Cwl_68_44 word68_44 gnd C_wl
Rw69_44 word69_44 word68_44 R_wl
Cwl_69_44 word69_44 gnd C_wl
Rw70_44 word70_44 word69_44 R_wl
Cwl_70_44 word70_44 gnd C_wl
Rw71_44 word71_44 word70_44 R_wl
Cwl_71_44 word71_44 gnd C_wl
Rw72_44 word72_44 word71_44 R_wl
Cwl_72_44 word72_44 gnd C_wl
Rw73_44 word73_44 word72_44 R_wl
Cwl_73_44 word73_44 gnd C_wl
Rw74_44 word74_44 word73_44 R_wl
Cwl_74_44 word74_44 gnd C_wl
Rw75_44 word75_44 word74_44 R_wl
Cwl_75_44 word75_44 gnd C_wl
Rw76_44 word76_44 word75_44 R_wl
Cwl_76_44 word76_44 gnd C_wl
Rw77_44 word77_44 word76_44 R_wl
Cwl_77_44 word77_44 gnd C_wl
Rw78_44 word78_44 word77_44 R_wl
Cwl_78_44 word78_44 gnd C_wl
Rw79_44 word79_44 word78_44 R_wl
Cwl_79_44 word79_44 gnd C_wl
Rw80_44 word80_44 word79_44 R_wl
Cwl_80_44 word80_44 gnd C_wl
Rw81_44 word81_44 word80_44 R_wl
Cwl_81_44 word81_44 gnd C_wl
Rw82_44 word82_44 word81_44 R_wl
Cwl_82_44 word82_44 gnd C_wl
Rw83_44 word83_44 word82_44 R_wl
Cwl_83_44 word83_44 gnd C_wl
Rw84_44 word84_44 word83_44 R_wl
Cwl_84_44 word84_44 gnd C_wl
Rw85_44 word85_44 word84_44 R_wl
Cwl_85_44 word85_44 gnd C_wl
Rw86_44 word86_44 word85_44 R_wl
Cwl_86_44 word86_44 gnd C_wl
Rw87_44 word87_44 word86_44 R_wl
Cwl_87_44 word87_44 gnd C_wl
Rw88_44 word88_44 word87_44 R_wl
Cwl_88_44 word88_44 gnd C_wl
Rw89_44 word89_44 word88_44 R_wl
Cwl_89_44 word89_44 gnd C_wl
Rw90_44 word90_44 word89_44 R_wl
Cwl_90_44 word90_44 gnd C_wl
Rw91_44 word91_44 word90_44 R_wl
Cwl_91_44 word91_44 gnd C_wl
Rw92_44 word92_44 word91_44 R_wl
Cwl_92_44 word92_44 gnd C_wl
Rw93_44 word93_44 word92_44 R_wl
Cwl_93_44 word93_44 gnd C_wl
Rw94_44 word94_44 word93_44 R_wl
Cwl_94_44 word94_44 gnd C_wl
Rw95_44 word95_44 word94_44 R_wl
Cwl_95_44 word95_44 gnd C_wl
Rw96_44 word96_44 word95_44 R_wl
Cwl_96_44 word96_44 gnd C_wl
Rw97_44 word97_44 word96_44 R_wl
Cwl_97_44 word97_44 gnd C_wl
Rw98_44 word98_44 word97_44 R_wl
Cwl_98_44 word98_44 gnd C_wl
Rw99_44 word99_44 word98_44 R_wl
Cwl_99_44 word99_44 gnd C_wl
Vwl_45 word_45 0 0
Rw0_45 word_45 word0_45 R_wl
Cwl_0_45 word0_45 gnd C_wl
Rw1_45 word1_45 word0_45 R_wl
Cwl_1_45 word1_45 gnd C_wl
Rw2_45 word2_45 word1_45 R_wl
Cwl_2_45 word2_45 gnd C_wl
Rw3_45 word3_45 word2_45 R_wl
Cwl_3_45 word3_45 gnd C_wl
Rw4_45 word4_45 word3_45 R_wl
Cwl_4_45 word4_45 gnd C_wl
Rw5_45 word5_45 word4_45 R_wl
Cwl_5_45 word5_45 gnd C_wl
Rw6_45 word6_45 word5_45 R_wl
Cwl_6_45 word6_45 gnd C_wl
Rw7_45 word7_45 word6_45 R_wl
Cwl_7_45 word7_45 gnd C_wl
Rw8_45 word8_45 word7_45 R_wl
Cwl_8_45 word8_45 gnd C_wl
Rw9_45 word9_45 word8_45 R_wl
Cwl_9_45 word9_45 gnd C_wl
Rw10_45 word10_45 word9_45 R_wl
Cwl_10_45 word10_45 gnd C_wl
Rw11_45 word11_45 word10_45 R_wl
Cwl_11_45 word11_45 gnd C_wl
Rw12_45 word12_45 word11_45 R_wl
Cwl_12_45 word12_45 gnd C_wl
Rw13_45 word13_45 word12_45 R_wl
Cwl_13_45 word13_45 gnd C_wl
Rw14_45 word14_45 word13_45 R_wl
Cwl_14_45 word14_45 gnd C_wl
Rw15_45 word15_45 word14_45 R_wl
Cwl_15_45 word15_45 gnd C_wl
Rw16_45 word16_45 word15_45 R_wl
Cwl_16_45 word16_45 gnd C_wl
Rw17_45 word17_45 word16_45 R_wl
Cwl_17_45 word17_45 gnd C_wl
Rw18_45 word18_45 word17_45 R_wl
Cwl_18_45 word18_45 gnd C_wl
Rw19_45 word19_45 word18_45 R_wl
Cwl_19_45 word19_45 gnd C_wl
Rw20_45 word20_45 word19_45 R_wl
Cwl_20_45 word20_45 gnd C_wl
Rw21_45 word21_45 word20_45 R_wl
Cwl_21_45 word21_45 gnd C_wl
Rw22_45 word22_45 word21_45 R_wl
Cwl_22_45 word22_45 gnd C_wl
Rw23_45 word23_45 word22_45 R_wl
Cwl_23_45 word23_45 gnd C_wl
Rw24_45 word24_45 word23_45 R_wl
Cwl_24_45 word24_45 gnd C_wl
Rw25_45 word25_45 word24_45 R_wl
Cwl_25_45 word25_45 gnd C_wl
Rw26_45 word26_45 word25_45 R_wl
Cwl_26_45 word26_45 gnd C_wl
Rw27_45 word27_45 word26_45 R_wl
Cwl_27_45 word27_45 gnd C_wl
Rw28_45 word28_45 word27_45 R_wl
Cwl_28_45 word28_45 gnd C_wl
Rw29_45 word29_45 word28_45 R_wl
Cwl_29_45 word29_45 gnd C_wl
Rw30_45 word30_45 word29_45 R_wl
Cwl_30_45 word30_45 gnd C_wl
Rw31_45 word31_45 word30_45 R_wl
Cwl_31_45 word31_45 gnd C_wl
Rw32_45 word32_45 word31_45 R_wl
Cwl_32_45 word32_45 gnd C_wl
Rw33_45 word33_45 word32_45 R_wl
Cwl_33_45 word33_45 gnd C_wl
Rw34_45 word34_45 word33_45 R_wl
Cwl_34_45 word34_45 gnd C_wl
Rw35_45 word35_45 word34_45 R_wl
Cwl_35_45 word35_45 gnd C_wl
Rw36_45 word36_45 word35_45 R_wl
Cwl_36_45 word36_45 gnd C_wl
Rw37_45 word37_45 word36_45 R_wl
Cwl_37_45 word37_45 gnd C_wl
Rw38_45 word38_45 word37_45 R_wl
Cwl_38_45 word38_45 gnd C_wl
Rw39_45 word39_45 word38_45 R_wl
Cwl_39_45 word39_45 gnd C_wl
Rw40_45 word40_45 word39_45 R_wl
Cwl_40_45 word40_45 gnd C_wl
Rw41_45 word41_45 word40_45 R_wl
Cwl_41_45 word41_45 gnd C_wl
Rw42_45 word42_45 word41_45 R_wl
Cwl_42_45 word42_45 gnd C_wl
Rw43_45 word43_45 word42_45 R_wl
Cwl_43_45 word43_45 gnd C_wl
Rw44_45 word44_45 word43_45 R_wl
Cwl_44_45 word44_45 gnd C_wl
Rw45_45 word45_45 word44_45 R_wl
Cwl_45_45 word45_45 gnd C_wl
Rw46_45 word46_45 word45_45 R_wl
Cwl_46_45 word46_45 gnd C_wl
Rw47_45 word47_45 word46_45 R_wl
Cwl_47_45 word47_45 gnd C_wl
Rw48_45 word48_45 word47_45 R_wl
Cwl_48_45 word48_45 gnd C_wl
Rw49_45 word49_45 word48_45 R_wl
Cwl_49_45 word49_45 gnd C_wl
Rw50_45 word50_45 word49_45 R_wl
Cwl_50_45 word50_45 gnd C_wl
Rw51_45 word51_45 word50_45 R_wl
Cwl_51_45 word51_45 gnd C_wl
Rw52_45 word52_45 word51_45 R_wl
Cwl_52_45 word52_45 gnd C_wl
Rw53_45 word53_45 word52_45 R_wl
Cwl_53_45 word53_45 gnd C_wl
Rw54_45 word54_45 word53_45 R_wl
Cwl_54_45 word54_45 gnd C_wl
Rw55_45 word55_45 word54_45 R_wl
Cwl_55_45 word55_45 gnd C_wl
Rw56_45 word56_45 word55_45 R_wl
Cwl_56_45 word56_45 gnd C_wl
Rw57_45 word57_45 word56_45 R_wl
Cwl_57_45 word57_45 gnd C_wl
Rw58_45 word58_45 word57_45 R_wl
Cwl_58_45 word58_45 gnd C_wl
Rw59_45 word59_45 word58_45 R_wl
Cwl_59_45 word59_45 gnd C_wl
Rw60_45 word60_45 word59_45 R_wl
Cwl_60_45 word60_45 gnd C_wl
Rw61_45 word61_45 word60_45 R_wl
Cwl_61_45 word61_45 gnd C_wl
Rw62_45 word62_45 word61_45 R_wl
Cwl_62_45 word62_45 gnd C_wl
Rw63_45 word63_45 word62_45 R_wl
Cwl_63_45 word63_45 gnd C_wl
Rw64_45 word64_45 word63_45 R_wl
Cwl_64_45 word64_45 gnd C_wl
Rw65_45 word65_45 word64_45 R_wl
Cwl_65_45 word65_45 gnd C_wl
Rw66_45 word66_45 word65_45 R_wl
Cwl_66_45 word66_45 gnd C_wl
Rw67_45 word67_45 word66_45 R_wl
Cwl_67_45 word67_45 gnd C_wl
Rw68_45 word68_45 word67_45 R_wl
Cwl_68_45 word68_45 gnd C_wl
Rw69_45 word69_45 word68_45 R_wl
Cwl_69_45 word69_45 gnd C_wl
Rw70_45 word70_45 word69_45 R_wl
Cwl_70_45 word70_45 gnd C_wl
Rw71_45 word71_45 word70_45 R_wl
Cwl_71_45 word71_45 gnd C_wl
Rw72_45 word72_45 word71_45 R_wl
Cwl_72_45 word72_45 gnd C_wl
Rw73_45 word73_45 word72_45 R_wl
Cwl_73_45 word73_45 gnd C_wl
Rw74_45 word74_45 word73_45 R_wl
Cwl_74_45 word74_45 gnd C_wl
Rw75_45 word75_45 word74_45 R_wl
Cwl_75_45 word75_45 gnd C_wl
Rw76_45 word76_45 word75_45 R_wl
Cwl_76_45 word76_45 gnd C_wl
Rw77_45 word77_45 word76_45 R_wl
Cwl_77_45 word77_45 gnd C_wl
Rw78_45 word78_45 word77_45 R_wl
Cwl_78_45 word78_45 gnd C_wl
Rw79_45 word79_45 word78_45 R_wl
Cwl_79_45 word79_45 gnd C_wl
Rw80_45 word80_45 word79_45 R_wl
Cwl_80_45 word80_45 gnd C_wl
Rw81_45 word81_45 word80_45 R_wl
Cwl_81_45 word81_45 gnd C_wl
Rw82_45 word82_45 word81_45 R_wl
Cwl_82_45 word82_45 gnd C_wl
Rw83_45 word83_45 word82_45 R_wl
Cwl_83_45 word83_45 gnd C_wl
Rw84_45 word84_45 word83_45 R_wl
Cwl_84_45 word84_45 gnd C_wl
Rw85_45 word85_45 word84_45 R_wl
Cwl_85_45 word85_45 gnd C_wl
Rw86_45 word86_45 word85_45 R_wl
Cwl_86_45 word86_45 gnd C_wl
Rw87_45 word87_45 word86_45 R_wl
Cwl_87_45 word87_45 gnd C_wl
Rw88_45 word88_45 word87_45 R_wl
Cwl_88_45 word88_45 gnd C_wl
Rw89_45 word89_45 word88_45 R_wl
Cwl_89_45 word89_45 gnd C_wl
Rw90_45 word90_45 word89_45 R_wl
Cwl_90_45 word90_45 gnd C_wl
Rw91_45 word91_45 word90_45 R_wl
Cwl_91_45 word91_45 gnd C_wl
Rw92_45 word92_45 word91_45 R_wl
Cwl_92_45 word92_45 gnd C_wl
Rw93_45 word93_45 word92_45 R_wl
Cwl_93_45 word93_45 gnd C_wl
Rw94_45 word94_45 word93_45 R_wl
Cwl_94_45 word94_45 gnd C_wl
Rw95_45 word95_45 word94_45 R_wl
Cwl_95_45 word95_45 gnd C_wl
Rw96_45 word96_45 word95_45 R_wl
Cwl_96_45 word96_45 gnd C_wl
Rw97_45 word97_45 word96_45 R_wl
Cwl_97_45 word97_45 gnd C_wl
Rw98_45 word98_45 word97_45 R_wl
Cwl_98_45 word98_45 gnd C_wl
Rw99_45 word99_45 word98_45 R_wl
Cwl_99_45 word99_45 gnd C_wl
Vwl_46 word_46 0 0
Rw0_46 word_46 word0_46 R_wl
Cwl_0_46 word0_46 gnd C_wl
Rw1_46 word1_46 word0_46 R_wl
Cwl_1_46 word1_46 gnd C_wl
Rw2_46 word2_46 word1_46 R_wl
Cwl_2_46 word2_46 gnd C_wl
Rw3_46 word3_46 word2_46 R_wl
Cwl_3_46 word3_46 gnd C_wl
Rw4_46 word4_46 word3_46 R_wl
Cwl_4_46 word4_46 gnd C_wl
Rw5_46 word5_46 word4_46 R_wl
Cwl_5_46 word5_46 gnd C_wl
Rw6_46 word6_46 word5_46 R_wl
Cwl_6_46 word6_46 gnd C_wl
Rw7_46 word7_46 word6_46 R_wl
Cwl_7_46 word7_46 gnd C_wl
Rw8_46 word8_46 word7_46 R_wl
Cwl_8_46 word8_46 gnd C_wl
Rw9_46 word9_46 word8_46 R_wl
Cwl_9_46 word9_46 gnd C_wl
Rw10_46 word10_46 word9_46 R_wl
Cwl_10_46 word10_46 gnd C_wl
Rw11_46 word11_46 word10_46 R_wl
Cwl_11_46 word11_46 gnd C_wl
Rw12_46 word12_46 word11_46 R_wl
Cwl_12_46 word12_46 gnd C_wl
Rw13_46 word13_46 word12_46 R_wl
Cwl_13_46 word13_46 gnd C_wl
Rw14_46 word14_46 word13_46 R_wl
Cwl_14_46 word14_46 gnd C_wl
Rw15_46 word15_46 word14_46 R_wl
Cwl_15_46 word15_46 gnd C_wl
Rw16_46 word16_46 word15_46 R_wl
Cwl_16_46 word16_46 gnd C_wl
Rw17_46 word17_46 word16_46 R_wl
Cwl_17_46 word17_46 gnd C_wl
Rw18_46 word18_46 word17_46 R_wl
Cwl_18_46 word18_46 gnd C_wl
Rw19_46 word19_46 word18_46 R_wl
Cwl_19_46 word19_46 gnd C_wl
Rw20_46 word20_46 word19_46 R_wl
Cwl_20_46 word20_46 gnd C_wl
Rw21_46 word21_46 word20_46 R_wl
Cwl_21_46 word21_46 gnd C_wl
Rw22_46 word22_46 word21_46 R_wl
Cwl_22_46 word22_46 gnd C_wl
Rw23_46 word23_46 word22_46 R_wl
Cwl_23_46 word23_46 gnd C_wl
Rw24_46 word24_46 word23_46 R_wl
Cwl_24_46 word24_46 gnd C_wl
Rw25_46 word25_46 word24_46 R_wl
Cwl_25_46 word25_46 gnd C_wl
Rw26_46 word26_46 word25_46 R_wl
Cwl_26_46 word26_46 gnd C_wl
Rw27_46 word27_46 word26_46 R_wl
Cwl_27_46 word27_46 gnd C_wl
Rw28_46 word28_46 word27_46 R_wl
Cwl_28_46 word28_46 gnd C_wl
Rw29_46 word29_46 word28_46 R_wl
Cwl_29_46 word29_46 gnd C_wl
Rw30_46 word30_46 word29_46 R_wl
Cwl_30_46 word30_46 gnd C_wl
Rw31_46 word31_46 word30_46 R_wl
Cwl_31_46 word31_46 gnd C_wl
Rw32_46 word32_46 word31_46 R_wl
Cwl_32_46 word32_46 gnd C_wl
Rw33_46 word33_46 word32_46 R_wl
Cwl_33_46 word33_46 gnd C_wl
Rw34_46 word34_46 word33_46 R_wl
Cwl_34_46 word34_46 gnd C_wl
Rw35_46 word35_46 word34_46 R_wl
Cwl_35_46 word35_46 gnd C_wl
Rw36_46 word36_46 word35_46 R_wl
Cwl_36_46 word36_46 gnd C_wl
Rw37_46 word37_46 word36_46 R_wl
Cwl_37_46 word37_46 gnd C_wl
Rw38_46 word38_46 word37_46 R_wl
Cwl_38_46 word38_46 gnd C_wl
Rw39_46 word39_46 word38_46 R_wl
Cwl_39_46 word39_46 gnd C_wl
Rw40_46 word40_46 word39_46 R_wl
Cwl_40_46 word40_46 gnd C_wl
Rw41_46 word41_46 word40_46 R_wl
Cwl_41_46 word41_46 gnd C_wl
Rw42_46 word42_46 word41_46 R_wl
Cwl_42_46 word42_46 gnd C_wl
Rw43_46 word43_46 word42_46 R_wl
Cwl_43_46 word43_46 gnd C_wl
Rw44_46 word44_46 word43_46 R_wl
Cwl_44_46 word44_46 gnd C_wl
Rw45_46 word45_46 word44_46 R_wl
Cwl_45_46 word45_46 gnd C_wl
Rw46_46 word46_46 word45_46 R_wl
Cwl_46_46 word46_46 gnd C_wl
Rw47_46 word47_46 word46_46 R_wl
Cwl_47_46 word47_46 gnd C_wl
Rw48_46 word48_46 word47_46 R_wl
Cwl_48_46 word48_46 gnd C_wl
Rw49_46 word49_46 word48_46 R_wl
Cwl_49_46 word49_46 gnd C_wl
Rw50_46 word50_46 word49_46 R_wl
Cwl_50_46 word50_46 gnd C_wl
Rw51_46 word51_46 word50_46 R_wl
Cwl_51_46 word51_46 gnd C_wl
Rw52_46 word52_46 word51_46 R_wl
Cwl_52_46 word52_46 gnd C_wl
Rw53_46 word53_46 word52_46 R_wl
Cwl_53_46 word53_46 gnd C_wl
Rw54_46 word54_46 word53_46 R_wl
Cwl_54_46 word54_46 gnd C_wl
Rw55_46 word55_46 word54_46 R_wl
Cwl_55_46 word55_46 gnd C_wl
Rw56_46 word56_46 word55_46 R_wl
Cwl_56_46 word56_46 gnd C_wl
Rw57_46 word57_46 word56_46 R_wl
Cwl_57_46 word57_46 gnd C_wl
Rw58_46 word58_46 word57_46 R_wl
Cwl_58_46 word58_46 gnd C_wl
Rw59_46 word59_46 word58_46 R_wl
Cwl_59_46 word59_46 gnd C_wl
Rw60_46 word60_46 word59_46 R_wl
Cwl_60_46 word60_46 gnd C_wl
Rw61_46 word61_46 word60_46 R_wl
Cwl_61_46 word61_46 gnd C_wl
Rw62_46 word62_46 word61_46 R_wl
Cwl_62_46 word62_46 gnd C_wl
Rw63_46 word63_46 word62_46 R_wl
Cwl_63_46 word63_46 gnd C_wl
Rw64_46 word64_46 word63_46 R_wl
Cwl_64_46 word64_46 gnd C_wl
Rw65_46 word65_46 word64_46 R_wl
Cwl_65_46 word65_46 gnd C_wl
Rw66_46 word66_46 word65_46 R_wl
Cwl_66_46 word66_46 gnd C_wl
Rw67_46 word67_46 word66_46 R_wl
Cwl_67_46 word67_46 gnd C_wl
Rw68_46 word68_46 word67_46 R_wl
Cwl_68_46 word68_46 gnd C_wl
Rw69_46 word69_46 word68_46 R_wl
Cwl_69_46 word69_46 gnd C_wl
Rw70_46 word70_46 word69_46 R_wl
Cwl_70_46 word70_46 gnd C_wl
Rw71_46 word71_46 word70_46 R_wl
Cwl_71_46 word71_46 gnd C_wl
Rw72_46 word72_46 word71_46 R_wl
Cwl_72_46 word72_46 gnd C_wl
Rw73_46 word73_46 word72_46 R_wl
Cwl_73_46 word73_46 gnd C_wl
Rw74_46 word74_46 word73_46 R_wl
Cwl_74_46 word74_46 gnd C_wl
Rw75_46 word75_46 word74_46 R_wl
Cwl_75_46 word75_46 gnd C_wl
Rw76_46 word76_46 word75_46 R_wl
Cwl_76_46 word76_46 gnd C_wl
Rw77_46 word77_46 word76_46 R_wl
Cwl_77_46 word77_46 gnd C_wl
Rw78_46 word78_46 word77_46 R_wl
Cwl_78_46 word78_46 gnd C_wl
Rw79_46 word79_46 word78_46 R_wl
Cwl_79_46 word79_46 gnd C_wl
Rw80_46 word80_46 word79_46 R_wl
Cwl_80_46 word80_46 gnd C_wl
Rw81_46 word81_46 word80_46 R_wl
Cwl_81_46 word81_46 gnd C_wl
Rw82_46 word82_46 word81_46 R_wl
Cwl_82_46 word82_46 gnd C_wl
Rw83_46 word83_46 word82_46 R_wl
Cwl_83_46 word83_46 gnd C_wl
Rw84_46 word84_46 word83_46 R_wl
Cwl_84_46 word84_46 gnd C_wl
Rw85_46 word85_46 word84_46 R_wl
Cwl_85_46 word85_46 gnd C_wl
Rw86_46 word86_46 word85_46 R_wl
Cwl_86_46 word86_46 gnd C_wl
Rw87_46 word87_46 word86_46 R_wl
Cwl_87_46 word87_46 gnd C_wl
Rw88_46 word88_46 word87_46 R_wl
Cwl_88_46 word88_46 gnd C_wl
Rw89_46 word89_46 word88_46 R_wl
Cwl_89_46 word89_46 gnd C_wl
Rw90_46 word90_46 word89_46 R_wl
Cwl_90_46 word90_46 gnd C_wl
Rw91_46 word91_46 word90_46 R_wl
Cwl_91_46 word91_46 gnd C_wl
Rw92_46 word92_46 word91_46 R_wl
Cwl_92_46 word92_46 gnd C_wl
Rw93_46 word93_46 word92_46 R_wl
Cwl_93_46 word93_46 gnd C_wl
Rw94_46 word94_46 word93_46 R_wl
Cwl_94_46 word94_46 gnd C_wl
Rw95_46 word95_46 word94_46 R_wl
Cwl_95_46 word95_46 gnd C_wl
Rw96_46 word96_46 word95_46 R_wl
Cwl_96_46 word96_46 gnd C_wl
Rw97_46 word97_46 word96_46 R_wl
Cwl_97_46 word97_46 gnd C_wl
Rw98_46 word98_46 word97_46 R_wl
Cwl_98_46 word98_46 gnd C_wl
Rw99_46 word99_46 word98_46 R_wl
Cwl_99_46 word99_46 gnd C_wl
Vwl_47 word_47 0 0
Rw0_47 word_47 word0_47 R_wl
Cwl_0_47 word0_47 gnd C_wl
Rw1_47 word1_47 word0_47 R_wl
Cwl_1_47 word1_47 gnd C_wl
Rw2_47 word2_47 word1_47 R_wl
Cwl_2_47 word2_47 gnd C_wl
Rw3_47 word3_47 word2_47 R_wl
Cwl_3_47 word3_47 gnd C_wl
Rw4_47 word4_47 word3_47 R_wl
Cwl_4_47 word4_47 gnd C_wl
Rw5_47 word5_47 word4_47 R_wl
Cwl_5_47 word5_47 gnd C_wl
Rw6_47 word6_47 word5_47 R_wl
Cwl_6_47 word6_47 gnd C_wl
Rw7_47 word7_47 word6_47 R_wl
Cwl_7_47 word7_47 gnd C_wl
Rw8_47 word8_47 word7_47 R_wl
Cwl_8_47 word8_47 gnd C_wl
Rw9_47 word9_47 word8_47 R_wl
Cwl_9_47 word9_47 gnd C_wl
Rw10_47 word10_47 word9_47 R_wl
Cwl_10_47 word10_47 gnd C_wl
Rw11_47 word11_47 word10_47 R_wl
Cwl_11_47 word11_47 gnd C_wl
Rw12_47 word12_47 word11_47 R_wl
Cwl_12_47 word12_47 gnd C_wl
Rw13_47 word13_47 word12_47 R_wl
Cwl_13_47 word13_47 gnd C_wl
Rw14_47 word14_47 word13_47 R_wl
Cwl_14_47 word14_47 gnd C_wl
Rw15_47 word15_47 word14_47 R_wl
Cwl_15_47 word15_47 gnd C_wl
Rw16_47 word16_47 word15_47 R_wl
Cwl_16_47 word16_47 gnd C_wl
Rw17_47 word17_47 word16_47 R_wl
Cwl_17_47 word17_47 gnd C_wl
Rw18_47 word18_47 word17_47 R_wl
Cwl_18_47 word18_47 gnd C_wl
Rw19_47 word19_47 word18_47 R_wl
Cwl_19_47 word19_47 gnd C_wl
Rw20_47 word20_47 word19_47 R_wl
Cwl_20_47 word20_47 gnd C_wl
Rw21_47 word21_47 word20_47 R_wl
Cwl_21_47 word21_47 gnd C_wl
Rw22_47 word22_47 word21_47 R_wl
Cwl_22_47 word22_47 gnd C_wl
Rw23_47 word23_47 word22_47 R_wl
Cwl_23_47 word23_47 gnd C_wl
Rw24_47 word24_47 word23_47 R_wl
Cwl_24_47 word24_47 gnd C_wl
Rw25_47 word25_47 word24_47 R_wl
Cwl_25_47 word25_47 gnd C_wl
Rw26_47 word26_47 word25_47 R_wl
Cwl_26_47 word26_47 gnd C_wl
Rw27_47 word27_47 word26_47 R_wl
Cwl_27_47 word27_47 gnd C_wl
Rw28_47 word28_47 word27_47 R_wl
Cwl_28_47 word28_47 gnd C_wl
Rw29_47 word29_47 word28_47 R_wl
Cwl_29_47 word29_47 gnd C_wl
Rw30_47 word30_47 word29_47 R_wl
Cwl_30_47 word30_47 gnd C_wl
Rw31_47 word31_47 word30_47 R_wl
Cwl_31_47 word31_47 gnd C_wl
Rw32_47 word32_47 word31_47 R_wl
Cwl_32_47 word32_47 gnd C_wl
Rw33_47 word33_47 word32_47 R_wl
Cwl_33_47 word33_47 gnd C_wl
Rw34_47 word34_47 word33_47 R_wl
Cwl_34_47 word34_47 gnd C_wl
Rw35_47 word35_47 word34_47 R_wl
Cwl_35_47 word35_47 gnd C_wl
Rw36_47 word36_47 word35_47 R_wl
Cwl_36_47 word36_47 gnd C_wl
Rw37_47 word37_47 word36_47 R_wl
Cwl_37_47 word37_47 gnd C_wl
Rw38_47 word38_47 word37_47 R_wl
Cwl_38_47 word38_47 gnd C_wl
Rw39_47 word39_47 word38_47 R_wl
Cwl_39_47 word39_47 gnd C_wl
Rw40_47 word40_47 word39_47 R_wl
Cwl_40_47 word40_47 gnd C_wl
Rw41_47 word41_47 word40_47 R_wl
Cwl_41_47 word41_47 gnd C_wl
Rw42_47 word42_47 word41_47 R_wl
Cwl_42_47 word42_47 gnd C_wl
Rw43_47 word43_47 word42_47 R_wl
Cwl_43_47 word43_47 gnd C_wl
Rw44_47 word44_47 word43_47 R_wl
Cwl_44_47 word44_47 gnd C_wl
Rw45_47 word45_47 word44_47 R_wl
Cwl_45_47 word45_47 gnd C_wl
Rw46_47 word46_47 word45_47 R_wl
Cwl_46_47 word46_47 gnd C_wl
Rw47_47 word47_47 word46_47 R_wl
Cwl_47_47 word47_47 gnd C_wl
Rw48_47 word48_47 word47_47 R_wl
Cwl_48_47 word48_47 gnd C_wl
Rw49_47 word49_47 word48_47 R_wl
Cwl_49_47 word49_47 gnd C_wl
Rw50_47 word50_47 word49_47 R_wl
Cwl_50_47 word50_47 gnd C_wl
Rw51_47 word51_47 word50_47 R_wl
Cwl_51_47 word51_47 gnd C_wl
Rw52_47 word52_47 word51_47 R_wl
Cwl_52_47 word52_47 gnd C_wl
Rw53_47 word53_47 word52_47 R_wl
Cwl_53_47 word53_47 gnd C_wl
Rw54_47 word54_47 word53_47 R_wl
Cwl_54_47 word54_47 gnd C_wl
Rw55_47 word55_47 word54_47 R_wl
Cwl_55_47 word55_47 gnd C_wl
Rw56_47 word56_47 word55_47 R_wl
Cwl_56_47 word56_47 gnd C_wl
Rw57_47 word57_47 word56_47 R_wl
Cwl_57_47 word57_47 gnd C_wl
Rw58_47 word58_47 word57_47 R_wl
Cwl_58_47 word58_47 gnd C_wl
Rw59_47 word59_47 word58_47 R_wl
Cwl_59_47 word59_47 gnd C_wl
Rw60_47 word60_47 word59_47 R_wl
Cwl_60_47 word60_47 gnd C_wl
Rw61_47 word61_47 word60_47 R_wl
Cwl_61_47 word61_47 gnd C_wl
Rw62_47 word62_47 word61_47 R_wl
Cwl_62_47 word62_47 gnd C_wl
Rw63_47 word63_47 word62_47 R_wl
Cwl_63_47 word63_47 gnd C_wl
Rw64_47 word64_47 word63_47 R_wl
Cwl_64_47 word64_47 gnd C_wl
Rw65_47 word65_47 word64_47 R_wl
Cwl_65_47 word65_47 gnd C_wl
Rw66_47 word66_47 word65_47 R_wl
Cwl_66_47 word66_47 gnd C_wl
Rw67_47 word67_47 word66_47 R_wl
Cwl_67_47 word67_47 gnd C_wl
Rw68_47 word68_47 word67_47 R_wl
Cwl_68_47 word68_47 gnd C_wl
Rw69_47 word69_47 word68_47 R_wl
Cwl_69_47 word69_47 gnd C_wl
Rw70_47 word70_47 word69_47 R_wl
Cwl_70_47 word70_47 gnd C_wl
Rw71_47 word71_47 word70_47 R_wl
Cwl_71_47 word71_47 gnd C_wl
Rw72_47 word72_47 word71_47 R_wl
Cwl_72_47 word72_47 gnd C_wl
Rw73_47 word73_47 word72_47 R_wl
Cwl_73_47 word73_47 gnd C_wl
Rw74_47 word74_47 word73_47 R_wl
Cwl_74_47 word74_47 gnd C_wl
Rw75_47 word75_47 word74_47 R_wl
Cwl_75_47 word75_47 gnd C_wl
Rw76_47 word76_47 word75_47 R_wl
Cwl_76_47 word76_47 gnd C_wl
Rw77_47 word77_47 word76_47 R_wl
Cwl_77_47 word77_47 gnd C_wl
Rw78_47 word78_47 word77_47 R_wl
Cwl_78_47 word78_47 gnd C_wl
Rw79_47 word79_47 word78_47 R_wl
Cwl_79_47 word79_47 gnd C_wl
Rw80_47 word80_47 word79_47 R_wl
Cwl_80_47 word80_47 gnd C_wl
Rw81_47 word81_47 word80_47 R_wl
Cwl_81_47 word81_47 gnd C_wl
Rw82_47 word82_47 word81_47 R_wl
Cwl_82_47 word82_47 gnd C_wl
Rw83_47 word83_47 word82_47 R_wl
Cwl_83_47 word83_47 gnd C_wl
Rw84_47 word84_47 word83_47 R_wl
Cwl_84_47 word84_47 gnd C_wl
Rw85_47 word85_47 word84_47 R_wl
Cwl_85_47 word85_47 gnd C_wl
Rw86_47 word86_47 word85_47 R_wl
Cwl_86_47 word86_47 gnd C_wl
Rw87_47 word87_47 word86_47 R_wl
Cwl_87_47 word87_47 gnd C_wl
Rw88_47 word88_47 word87_47 R_wl
Cwl_88_47 word88_47 gnd C_wl
Rw89_47 word89_47 word88_47 R_wl
Cwl_89_47 word89_47 gnd C_wl
Rw90_47 word90_47 word89_47 R_wl
Cwl_90_47 word90_47 gnd C_wl
Rw91_47 word91_47 word90_47 R_wl
Cwl_91_47 word91_47 gnd C_wl
Rw92_47 word92_47 word91_47 R_wl
Cwl_92_47 word92_47 gnd C_wl
Rw93_47 word93_47 word92_47 R_wl
Cwl_93_47 word93_47 gnd C_wl
Rw94_47 word94_47 word93_47 R_wl
Cwl_94_47 word94_47 gnd C_wl
Rw95_47 word95_47 word94_47 R_wl
Cwl_95_47 word95_47 gnd C_wl
Rw96_47 word96_47 word95_47 R_wl
Cwl_96_47 word96_47 gnd C_wl
Rw97_47 word97_47 word96_47 R_wl
Cwl_97_47 word97_47 gnd C_wl
Rw98_47 word98_47 word97_47 R_wl
Cwl_98_47 word98_47 gnd C_wl
Rw99_47 word99_47 word98_47 R_wl
Cwl_99_47 word99_47 gnd C_wl
Vwl_48 word_48 0 0
Rw0_48 word_48 word0_48 R_wl
Cwl_0_48 word0_48 gnd C_wl
Rw1_48 word1_48 word0_48 R_wl
Cwl_1_48 word1_48 gnd C_wl
Rw2_48 word2_48 word1_48 R_wl
Cwl_2_48 word2_48 gnd C_wl
Rw3_48 word3_48 word2_48 R_wl
Cwl_3_48 word3_48 gnd C_wl
Rw4_48 word4_48 word3_48 R_wl
Cwl_4_48 word4_48 gnd C_wl
Rw5_48 word5_48 word4_48 R_wl
Cwl_5_48 word5_48 gnd C_wl
Rw6_48 word6_48 word5_48 R_wl
Cwl_6_48 word6_48 gnd C_wl
Rw7_48 word7_48 word6_48 R_wl
Cwl_7_48 word7_48 gnd C_wl
Rw8_48 word8_48 word7_48 R_wl
Cwl_8_48 word8_48 gnd C_wl
Rw9_48 word9_48 word8_48 R_wl
Cwl_9_48 word9_48 gnd C_wl
Rw10_48 word10_48 word9_48 R_wl
Cwl_10_48 word10_48 gnd C_wl
Rw11_48 word11_48 word10_48 R_wl
Cwl_11_48 word11_48 gnd C_wl
Rw12_48 word12_48 word11_48 R_wl
Cwl_12_48 word12_48 gnd C_wl
Rw13_48 word13_48 word12_48 R_wl
Cwl_13_48 word13_48 gnd C_wl
Rw14_48 word14_48 word13_48 R_wl
Cwl_14_48 word14_48 gnd C_wl
Rw15_48 word15_48 word14_48 R_wl
Cwl_15_48 word15_48 gnd C_wl
Rw16_48 word16_48 word15_48 R_wl
Cwl_16_48 word16_48 gnd C_wl
Rw17_48 word17_48 word16_48 R_wl
Cwl_17_48 word17_48 gnd C_wl
Rw18_48 word18_48 word17_48 R_wl
Cwl_18_48 word18_48 gnd C_wl
Rw19_48 word19_48 word18_48 R_wl
Cwl_19_48 word19_48 gnd C_wl
Rw20_48 word20_48 word19_48 R_wl
Cwl_20_48 word20_48 gnd C_wl
Rw21_48 word21_48 word20_48 R_wl
Cwl_21_48 word21_48 gnd C_wl
Rw22_48 word22_48 word21_48 R_wl
Cwl_22_48 word22_48 gnd C_wl
Rw23_48 word23_48 word22_48 R_wl
Cwl_23_48 word23_48 gnd C_wl
Rw24_48 word24_48 word23_48 R_wl
Cwl_24_48 word24_48 gnd C_wl
Rw25_48 word25_48 word24_48 R_wl
Cwl_25_48 word25_48 gnd C_wl
Rw26_48 word26_48 word25_48 R_wl
Cwl_26_48 word26_48 gnd C_wl
Rw27_48 word27_48 word26_48 R_wl
Cwl_27_48 word27_48 gnd C_wl
Rw28_48 word28_48 word27_48 R_wl
Cwl_28_48 word28_48 gnd C_wl
Rw29_48 word29_48 word28_48 R_wl
Cwl_29_48 word29_48 gnd C_wl
Rw30_48 word30_48 word29_48 R_wl
Cwl_30_48 word30_48 gnd C_wl
Rw31_48 word31_48 word30_48 R_wl
Cwl_31_48 word31_48 gnd C_wl
Rw32_48 word32_48 word31_48 R_wl
Cwl_32_48 word32_48 gnd C_wl
Rw33_48 word33_48 word32_48 R_wl
Cwl_33_48 word33_48 gnd C_wl
Rw34_48 word34_48 word33_48 R_wl
Cwl_34_48 word34_48 gnd C_wl
Rw35_48 word35_48 word34_48 R_wl
Cwl_35_48 word35_48 gnd C_wl
Rw36_48 word36_48 word35_48 R_wl
Cwl_36_48 word36_48 gnd C_wl
Rw37_48 word37_48 word36_48 R_wl
Cwl_37_48 word37_48 gnd C_wl
Rw38_48 word38_48 word37_48 R_wl
Cwl_38_48 word38_48 gnd C_wl
Rw39_48 word39_48 word38_48 R_wl
Cwl_39_48 word39_48 gnd C_wl
Rw40_48 word40_48 word39_48 R_wl
Cwl_40_48 word40_48 gnd C_wl
Rw41_48 word41_48 word40_48 R_wl
Cwl_41_48 word41_48 gnd C_wl
Rw42_48 word42_48 word41_48 R_wl
Cwl_42_48 word42_48 gnd C_wl
Rw43_48 word43_48 word42_48 R_wl
Cwl_43_48 word43_48 gnd C_wl
Rw44_48 word44_48 word43_48 R_wl
Cwl_44_48 word44_48 gnd C_wl
Rw45_48 word45_48 word44_48 R_wl
Cwl_45_48 word45_48 gnd C_wl
Rw46_48 word46_48 word45_48 R_wl
Cwl_46_48 word46_48 gnd C_wl
Rw47_48 word47_48 word46_48 R_wl
Cwl_47_48 word47_48 gnd C_wl
Rw48_48 word48_48 word47_48 R_wl
Cwl_48_48 word48_48 gnd C_wl
Rw49_48 word49_48 word48_48 R_wl
Cwl_49_48 word49_48 gnd C_wl
Rw50_48 word50_48 word49_48 R_wl
Cwl_50_48 word50_48 gnd C_wl
Rw51_48 word51_48 word50_48 R_wl
Cwl_51_48 word51_48 gnd C_wl
Rw52_48 word52_48 word51_48 R_wl
Cwl_52_48 word52_48 gnd C_wl
Rw53_48 word53_48 word52_48 R_wl
Cwl_53_48 word53_48 gnd C_wl
Rw54_48 word54_48 word53_48 R_wl
Cwl_54_48 word54_48 gnd C_wl
Rw55_48 word55_48 word54_48 R_wl
Cwl_55_48 word55_48 gnd C_wl
Rw56_48 word56_48 word55_48 R_wl
Cwl_56_48 word56_48 gnd C_wl
Rw57_48 word57_48 word56_48 R_wl
Cwl_57_48 word57_48 gnd C_wl
Rw58_48 word58_48 word57_48 R_wl
Cwl_58_48 word58_48 gnd C_wl
Rw59_48 word59_48 word58_48 R_wl
Cwl_59_48 word59_48 gnd C_wl
Rw60_48 word60_48 word59_48 R_wl
Cwl_60_48 word60_48 gnd C_wl
Rw61_48 word61_48 word60_48 R_wl
Cwl_61_48 word61_48 gnd C_wl
Rw62_48 word62_48 word61_48 R_wl
Cwl_62_48 word62_48 gnd C_wl
Rw63_48 word63_48 word62_48 R_wl
Cwl_63_48 word63_48 gnd C_wl
Rw64_48 word64_48 word63_48 R_wl
Cwl_64_48 word64_48 gnd C_wl
Rw65_48 word65_48 word64_48 R_wl
Cwl_65_48 word65_48 gnd C_wl
Rw66_48 word66_48 word65_48 R_wl
Cwl_66_48 word66_48 gnd C_wl
Rw67_48 word67_48 word66_48 R_wl
Cwl_67_48 word67_48 gnd C_wl
Rw68_48 word68_48 word67_48 R_wl
Cwl_68_48 word68_48 gnd C_wl
Rw69_48 word69_48 word68_48 R_wl
Cwl_69_48 word69_48 gnd C_wl
Rw70_48 word70_48 word69_48 R_wl
Cwl_70_48 word70_48 gnd C_wl
Rw71_48 word71_48 word70_48 R_wl
Cwl_71_48 word71_48 gnd C_wl
Rw72_48 word72_48 word71_48 R_wl
Cwl_72_48 word72_48 gnd C_wl
Rw73_48 word73_48 word72_48 R_wl
Cwl_73_48 word73_48 gnd C_wl
Rw74_48 word74_48 word73_48 R_wl
Cwl_74_48 word74_48 gnd C_wl
Rw75_48 word75_48 word74_48 R_wl
Cwl_75_48 word75_48 gnd C_wl
Rw76_48 word76_48 word75_48 R_wl
Cwl_76_48 word76_48 gnd C_wl
Rw77_48 word77_48 word76_48 R_wl
Cwl_77_48 word77_48 gnd C_wl
Rw78_48 word78_48 word77_48 R_wl
Cwl_78_48 word78_48 gnd C_wl
Rw79_48 word79_48 word78_48 R_wl
Cwl_79_48 word79_48 gnd C_wl
Rw80_48 word80_48 word79_48 R_wl
Cwl_80_48 word80_48 gnd C_wl
Rw81_48 word81_48 word80_48 R_wl
Cwl_81_48 word81_48 gnd C_wl
Rw82_48 word82_48 word81_48 R_wl
Cwl_82_48 word82_48 gnd C_wl
Rw83_48 word83_48 word82_48 R_wl
Cwl_83_48 word83_48 gnd C_wl
Rw84_48 word84_48 word83_48 R_wl
Cwl_84_48 word84_48 gnd C_wl
Rw85_48 word85_48 word84_48 R_wl
Cwl_85_48 word85_48 gnd C_wl
Rw86_48 word86_48 word85_48 R_wl
Cwl_86_48 word86_48 gnd C_wl
Rw87_48 word87_48 word86_48 R_wl
Cwl_87_48 word87_48 gnd C_wl
Rw88_48 word88_48 word87_48 R_wl
Cwl_88_48 word88_48 gnd C_wl
Rw89_48 word89_48 word88_48 R_wl
Cwl_89_48 word89_48 gnd C_wl
Rw90_48 word90_48 word89_48 R_wl
Cwl_90_48 word90_48 gnd C_wl
Rw91_48 word91_48 word90_48 R_wl
Cwl_91_48 word91_48 gnd C_wl
Rw92_48 word92_48 word91_48 R_wl
Cwl_92_48 word92_48 gnd C_wl
Rw93_48 word93_48 word92_48 R_wl
Cwl_93_48 word93_48 gnd C_wl
Rw94_48 word94_48 word93_48 R_wl
Cwl_94_48 word94_48 gnd C_wl
Rw95_48 word95_48 word94_48 R_wl
Cwl_95_48 word95_48 gnd C_wl
Rw96_48 word96_48 word95_48 R_wl
Cwl_96_48 word96_48 gnd C_wl
Rw97_48 word97_48 word96_48 R_wl
Cwl_97_48 word97_48 gnd C_wl
Rw98_48 word98_48 word97_48 R_wl
Cwl_98_48 word98_48 gnd C_wl
Rw99_48 word99_48 word98_48 R_wl
Cwl_99_48 word99_48 gnd C_wl
Vwl_49 word_49 0 0
Rw0_49 word_49 word0_49 R_wl
Cwl_0_49 word0_49 gnd C_wl
Rw1_49 word1_49 word0_49 R_wl
Cwl_1_49 word1_49 gnd C_wl
Rw2_49 word2_49 word1_49 R_wl
Cwl_2_49 word2_49 gnd C_wl
Rw3_49 word3_49 word2_49 R_wl
Cwl_3_49 word3_49 gnd C_wl
Rw4_49 word4_49 word3_49 R_wl
Cwl_4_49 word4_49 gnd C_wl
Rw5_49 word5_49 word4_49 R_wl
Cwl_5_49 word5_49 gnd C_wl
Rw6_49 word6_49 word5_49 R_wl
Cwl_6_49 word6_49 gnd C_wl
Rw7_49 word7_49 word6_49 R_wl
Cwl_7_49 word7_49 gnd C_wl
Rw8_49 word8_49 word7_49 R_wl
Cwl_8_49 word8_49 gnd C_wl
Rw9_49 word9_49 word8_49 R_wl
Cwl_9_49 word9_49 gnd C_wl
Rw10_49 word10_49 word9_49 R_wl
Cwl_10_49 word10_49 gnd C_wl
Rw11_49 word11_49 word10_49 R_wl
Cwl_11_49 word11_49 gnd C_wl
Rw12_49 word12_49 word11_49 R_wl
Cwl_12_49 word12_49 gnd C_wl
Rw13_49 word13_49 word12_49 R_wl
Cwl_13_49 word13_49 gnd C_wl
Rw14_49 word14_49 word13_49 R_wl
Cwl_14_49 word14_49 gnd C_wl
Rw15_49 word15_49 word14_49 R_wl
Cwl_15_49 word15_49 gnd C_wl
Rw16_49 word16_49 word15_49 R_wl
Cwl_16_49 word16_49 gnd C_wl
Rw17_49 word17_49 word16_49 R_wl
Cwl_17_49 word17_49 gnd C_wl
Rw18_49 word18_49 word17_49 R_wl
Cwl_18_49 word18_49 gnd C_wl
Rw19_49 word19_49 word18_49 R_wl
Cwl_19_49 word19_49 gnd C_wl
Rw20_49 word20_49 word19_49 R_wl
Cwl_20_49 word20_49 gnd C_wl
Rw21_49 word21_49 word20_49 R_wl
Cwl_21_49 word21_49 gnd C_wl
Rw22_49 word22_49 word21_49 R_wl
Cwl_22_49 word22_49 gnd C_wl
Rw23_49 word23_49 word22_49 R_wl
Cwl_23_49 word23_49 gnd C_wl
Rw24_49 word24_49 word23_49 R_wl
Cwl_24_49 word24_49 gnd C_wl
Rw25_49 word25_49 word24_49 R_wl
Cwl_25_49 word25_49 gnd C_wl
Rw26_49 word26_49 word25_49 R_wl
Cwl_26_49 word26_49 gnd C_wl
Rw27_49 word27_49 word26_49 R_wl
Cwl_27_49 word27_49 gnd C_wl
Rw28_49 word28_49 word27_49 R_wl
Cwl_28_49 word28_49 gnd C_wl
Rw29_49 word29_49 word28_49 R_wl
Cwl_29_49 word29_49 gnd C_wl
Rw30_49 word30_49 word29_49 R_wl
Cwl_30_49 word30_49 gnd C_wl
Rw31_49 word31_49 word30_49 R_wl
Cwl_31_49 word31_49 gnd C_wl
Rw32_49 word32_49 word31_49 R_wl
Cwl_32_49 word32_49 gnd C_wl
Rw33_49 word33_49 word32_49 R_wl
Cwl_33_49 word33_49 gnd C_wl
Rw34_49 word34_49 word33_49 R_wl
Cwl_34_49 word34_49 gnd C_wl
Rw35_49 word35_49 word34_49 R_wl
Cwl_35_49 word35_49 gnd C_wl
Rw36_49 word36_49 word35_49 R_wl
Cwl_36_49 word36_49 gnd C_wl
Rw37_49 word37_49 word36_49 R_wl
Cwl_37_49 word37_49 gnd C_wl
Rw38_49 word38_49 word37_49 R_wl
Cwl_38_49 word38_49 gnd C_wl
Rw39_49 word39_49 word38_49 R_wl
Cwl_39_49 word39_49 gnd C_wl
Rw40_49 word40_49 word39_49 R_wl
Cwl_40_49 word40_49 gnd C_wl
Rw41_49 word41_49 word40_49 R_wl
Cwl_41_49 word41_49 gnd C_wl
Rw42_49 word42_49 word41_49 R_wl
Cwl_42_49 word42_49 gnd C_wl
Rw43_49 word43_49 word42_49 R_wl
Cwl_43_49 word43_49 gnd C_wl
Rw44_49 word44_49 word43_49 R_wl
Cwl_44_49 word44_49 gnd C_wl
Rw45_49 word45_49 word44_49 R_wl
Cwl_45_49 word45_49 gnd C_wl
Rw46_49 word46_49 word45_49 R_wl
Cwl_46_49 word46_49 gnd C_wl
Rw47_49 word47_49 word46_49 R_wl
Cwl_47_49 word47_49 gnd C_wl
Rw48_49 word48_49 word47_49 R_wl
Cwl_48_49 word48_49 gnd C_wl
Rw49_49 word49_49 word48_49 R_wl
Cwl_49_49 word49_49 gnd C_wl
Rw50_49 word50_49 word49_49 R_wl
Cwl_50_49 word50_49 gnd C_wl
Rw51_49 word51_49 word50_49 R_wl
Cwl_51_49 word51_49 gnd C_wl
Rw52_49 word52_49 word51_49 R_wl
Cwl_52_49 word52_49 gnd C_wl
Rw53_49 word53_49 word52_49 R_wl
Cwl_53_49 word53_49 gnd C_wl
Rw54_49 word54_49 word53_49 R_wl
Cwl_54_49 word54_49 gnd C_wl
Rw55_49 word55_49 word54_49 R_wl
Cwl_55_49 word55_49 gnd C_wl
Rw56_49 word56_49 word55_49 R_wl
Cwl_56_49 word56_49 gnd C_wl
Rw57_49 word57_49 word56_49 R_wl
Cwl_57_49 word57_49 gnd C_wl
Rw58_49 word58_49 word57_49 R_wl
Cwl_58_49 word58_49 gnd C_wl
Rw59_49 word59_49 word58_49 R_wl
Cwl_59_49 word59_49 gnd C_wl
Rw60_49 word60_49 word59_49 R_wl
Cwl_60_49 word60_49 gnd C_wl
Rw61_49 word61_49 word60_49 R_wl
Cwl_61_49 word61_49 gnd C_wl
Rw62_49 word62_49 word61_49 R_wl
Cwl_62_49 word62_49 gnd C_wl
Rw63_49 word63_49 word62_49 R_wl
Cwl_63_49 word63_49 gnd C_wl
Rw64_49 word64_49 word63_49 R_wl
Cwl_64_49 word64_49 gnd C_wl
Rw65_49 word65_49 word64_49 R_wl
Cwl_65_49 word65_49 gnd C_wl
Rw66_49 word66_49 word65_49 R_wl
Cwl_66_49 word66_49 gnd C_wl
Rw67_49 word67_49 word66_49 R_wl
Cwl_67_49 word67_49 gnd C_wl
Rw68_49 word68_49 word67_49 R_wl
Cwl_68_49 word68_49 gnd C_wl
Rw69_49 word69_49 word68_49 R_wl
Cwl_69_49 word69_49 gnd C_wl
Rw70_49 word70_49 word69_49 R_wl
Cwl_70_49 word70_49 gnd C_wl
Rw71_49 word71_49 word70_49 R_wl
Cwl_71_49 word71_49 gnd C_wl
Rw72_49 word72_49 word71_49 R_wl
Cwl_72_49 word72_49 gnd C_wl
Rw73_49 word73_49 word72_49 R_wl
Cwl_73_49 word73_49 gnd C_wl
Rw74_49 word74_49 word73_49 R_wl
Cwl_74_49 word74_49 gnd C_wl
Rw75_49 word75_49 word74_49 R_wl
Cwl_75_49 word75_49 gnd C_wl
Rw76_49 word76_49 word75_49 R_wl
Cwl_76_49 word76_49 gnd C_wl
Rw77_49 word77_49 word76_49 R_wl
Cwl_77_49 word77_49 gnd C_wl
Rw78_49 word78_49 word77_49 R_wl
Cwl_78_49 word78_49 gnd C_wl
Rw79_49 word79_49 word78_49 R_wl
Cwl_79_49 word79_49 gnd C_wl
Rw80_49 word80_49 word79_49 R_wl
Cwl_80_49 word80_49 gnd C_wl
Rw81_49 word81_49 word80_49 R_wl
Cwl_81_49 word81_49 gnd C_wl
Rw82_49 word82_49 word81_49 R_wl
Cwl_82_49 word82_49 gnd C_wl
Rw83_49 word83_49 word82_49 R_wl
Cwl_83_49 word83_49 gnd C_wl
Rw84_49 word84_49 word83_49 R_wl
Cwl_84_49 word84_49 gnd C_wl
Rw85_49 word85_49 word84_49 R_wl
Cwl_85_49 word85_49 gnd C_wl
Rw86_49 word86_49 word85_49 R_wl
Cwl_86_49 word86_49 gnd C_wl
Rw87_49 word87_49 word86_49 R_wl
Cwl_87_49 word87_49 gnd C_wl
Rw88_49 word88_49 word87_49 R_wl
Cwl_88_49 word88_49 gnd C_wl
Rw89_49 word89_49 word88_49 R_wl
Cwl_89_49 word89_49 gnd C_wl
Rw90_49 word90_49 word89_49 R_wl
Cwl_90_49 word90_49 gnd C_wl
Rw91_49 word91_49 word90_49 R_wl
Cwl_91_49 word91_49 gnd C_wl
Rw92_49 word92_49 word91_49 R_wl
Cwl_92_49 word92_49 gnd C_wl
Rw93_49 word93_49 word92_49 R_wl
Cwl_93_49 word93_49 gnd C_wl
Rw94_49 word94_49 word93_49 R_wl
Cwl_94_49 word94_49 gnd C_wl
Rw95_49 word95_49 word94_49 R_wl
Cwl_95_49 word95_49 gnd C_wl
Rw96_49 word96_49 word95_49 R_wl
Cwl_96_49 word96_49 gnd C_wl
Rw97_49 word97_49 word96_49 R_wl
Cwl_97_49 word97_49 gnd C_wl
Rw98_49 word98_49 word97_49 R_wl
Cwl_98_49 word98_49 gnd C_wl
Rw99_49 word99_49 word98_49 R_wl
Cwl_99_49 word99_49 gnd C_wl
Vwl_50 word_50 0 0
Rw0_50 word_50 word0_50 R_wl
Cwl_0_50 word0_50 gnd C_wl
Rw1_50 word1_50 word0_50 R_wl
Cwl_1_50 word1_50 gnd C_wl
Rw2_50 word2_50 word1_50 R_wl
Cwl_2_50 word2_50 gnd C_wl
Rw3_50 word3_50 word2_50 R_wl
Cwl_3_50 word3_50 gnd C_wl
Rw4_50 word4_50 word3_50 R_wl
Cwl_4_50 word4_50 gnd C_wl
Rw5_50 word5_50 word4_50 R_wl
Cwl_5_50 word5_50 gnd C_wl
Rw6_50 word6_50 word5_50 R_wl
Cwl_6_50 word6_50 gnd C_wl
Rw7_50 word7_50 word6_50 R_wl
Cwl_7_50 word7_50 gnd C_wl
Rw8_50 word8_50 word7_50 R_wl
Cwl_8_50 word8_50 gnd C_wl
Rw9_50 word9_50 word8_50 R_wl
Cwl_9_50 word9_50 gnd C_wl
Rw10_50 word10_50 word9_50 R_wl
Cwl_10_50 word10_50 gnd C_wl
Rw11_50 word11_50 word10_50 R_wl
Cwl_11_50 word11_50 gnd C_wl
Rw12_50 word12_50 word11_50 R_wl
Cwl_12_50 word12_50 gnd C_wl
Rw13_50 word13_50 word12_50 R_wl
Cwl_13_50 word13_50 gnd C_wl
Rw14_50 word14_50 word13_50 R_wl
Cwl_14_50 word14_50 gnd C_wl
Rw15_50 word15_50 word14_50 R_wl
Cwl_15_50 word15_50 gnd C_wl
Rw16_50 word16_50 word15_50 R_wl
Cwl_16_50 word16_50 gnd C_wl
Rw17_50 word17_50 word16_50 R_wl
Cwl_17_50 word17_50 gnd C_wl
Rw18_50 word18_50 word17_50 R_wl
Cwl_18_50 word18_50 gnd C_wl
Rw19_50 word19_50 word18_50 R_wl
Cwl_19_50 word19_50 gnd C_wl
Rw20_50 word20_50 word19_50 R_wl
Cwl_20_50 word20_50 gnd C_wl
Rw21_50 word21_50 word20_50 R_wl
Cwl_21_50 word21_50 gnd C_wl
Rw22_50 word22_50 word21_50 R_wl
Cwl_22_50 word22_50 gnd C_wl
Rw23_50 word23_50 word22_50 R_wl
Cwl_23_50 word23_50 gnd C_wl
Rw24_50 word24_50 word23_50 R_wl
Cwl_24_50 word24_50 gnd C_wl
Rw25_50 word25_50 word24_50 R_wl
Cwl_25_50 word25_50 gnd C_wl
Rw26_50 word26_50 word25_50 R_wl
Cwl_26_50 word26_50 gnd C_wl
Rw27_50 word27_50 word26_50 R_wl
Cwl_27_50 word27_50 gnd C_wl
Rw28_50 word28_50 word27_50 R_wl
Cwl_28_50 word28_50 gnd C_wl
Rw29_50 word29_50 word28_50 R_wl
Cwl_29_50 word29_50 gnd C_wl
Rw30_50 word30_50 word29_50 R_wl
Cwl_30_50 word30_50 gnd C_wl
Rw31_50 word31_50 word30_50 R_wl
Cwl_31_50 word31_50 gnd C_wl
Rw32_50 word32_50 word31_50 R_wl
Cwl_32_50 word32_50 gnd C_wl
Rw33_50 word33_50 word32_50 R_wl
Cwl_33_50 word33_50 gnd C_wl
Rw34_50 word34_50 word33_50 R_wl
Cwl_34_50 word34_50 gnd C_wl
Rw35_50 word35_50 word34_50 R_wl
Cwl_35_50 word35_50 gnd C_wl
Rw36_50 word36_50 word35_50 R_wl
Cwl_36_50 word36_50 gnd C_wl
Rw37_50 word37_50 word36_50 R_wl
Cwl_37_50 word37_50 gnd C_wl
Rw38_50 word38_50 word37_50 R_wl
Cwl_38_50 word38_50 gnd C_wl
Rw39_50 word39_50 word38_50 R_wl
Cwl_39_50 word39_50 gnd C_wl
Rw40_50 word40_50 word39_50 R_wl
Cwl_40_50 word40_50 gnd C_wl
Rw41_50 word41_50 word40_50 R_wl
Cwl_41_50 word41_50 gnd C_wl
Rw42_50 word42_50 word41_50 R_wl
Cwl_42_50 word42_50 gnd C_wl
Rw43_50 word43_50 word42_50 R_wl
Cwl_43_50 word43_50 gnd C_wl
Rw44_50 word44_50 word43_50 R_wl
Cwl_44_50 word44_50 gnd C_wl
Rw45_50 word45_50 word44_50 R_wl
Cwl_45_50 word45_50 gnd C_wl
Rw46_50 word46_50 word45_50 R_wl
Cwl_46_50 word46_50 gnd C_wl
Rw47_50 word47_50 word46_50 R_wl
Cwl_47_50 word47_50 gnd C_wl
Rw48_50 word48_50 word47_50 R_wl
Cwl_48_50 word48_50 gnd C_wl
Rw49_50 word49_50 word48_50 R_wl
Cwl_49_50 word49_50 gnd C_wl
Rw50_50 word50_50 word49_50 R_wl
Cwl_50_50 word50_50 gnd C_wl
Rw51_50 word51_50 word50_50 R_wl
Cwl_51_50 word51_50 gnd C_wl
Rw52_50 word52_50 word51_50 R_wl
Cwl_52_50 word52_50 gnd C_wl
Rw53_50 word53_50 word52_50 R_wl
Cwl_53_50 word53_50 gnd C_wl
Rw54_50 word54_50 word53_50 R_wl
Cwl_54_50 word54_50 gnd C_wl
Rw55_50 word55_50 word54_50 R_wl
Cwl_55_50 word55_50 gnd C_wl
Rw56_50 word56_50 word55_50 R_wl
Cwl_56_50 word56_50 gnd C_wl
Rw57_50 word57_50 word56_50 R_wl
Cwl_57_50 word57_50 gnd C_wl
Rw58_50 word58_50 word57_50 R_wl
Cwl_58_50 word58_50 gnd C_wl
Rw59_50 word59_50 word58_50 R_wl
Cwl_59_50 word59_50 gnd C_wl
Rw60_50 word60_50 word59_50 R_wl
Cwl_60_50 word60_50 gnd C_wl
Rw61_50 word61_50 word60_50 R_wl
Cwl_61_50 word61_50 gnd C_wl
Rw62_50 word62_50 word61_50 R_wl
Cwl_62_50 word62_50 gnd C_wl
Rw63_50 word63_50 word62_50 R_wl
Cwl_63_50 word63_50 gnd C_wl
Rw64_50 word64_50 word63_50 R_wl
Cwl_64_50 word64_50 gnd C_wl
Rw65_50 word65_50 word64_50 R_wl
Cwl_65_50 word65_50 gnd C_wl
Rw66_50 word66_50 word65_50 R_wl
Cwl_66_50 word66_50 gnd C_wl
Rw67_50 word67_50 word66_50 R_wl
Cwl_67_50 word67_50 gnd C_wl
Rw68_50 word68_50 word67_50 R_wl
Cwl_68_50 word68_50 gnd C_wl
Rw69_50 word69_50 word68_50 R_wl
Cwl_69_50 word69_50 gnd C_wl
Rw70_50 word70_50 word69_50 R_wl
Cwl_70_50 word70_50 gnd C_wl
Rw71_50 word71_50 word70_50 R_wl
Cwl_71_50 word71_50 gnd C_wl
Rw72_50 word72_50 word71_50 R_wl
Cwl_72_50 word72_50 gnd C_wl
Rw73_50 word73_50 word72_50 R_wl
Cwl_73_50 word73_50 gnd C_wl
Rw74_50 word74_50 word73_50 R_wl
Cwl_74_50 word74_50 gnd C_wl
Rw75_50 word75_50 word74_50 R_wl
Cwl_75_50 word75_50 gnd C_wl
Rw76_50 word76_50 word75_50 R_wl
Cwl_76_50 word76_50 gnd C_wl
Rw77_50 word77_50 word76_50 R_wl
Cwl_77_50 word77_50 gnd C_wl
Rw78_50 word78_50 word77_50 R_wl
Cwl_78_50 word78_50 gnd C_wl
Rw79_50 word79_50 word78_50 R_wl
Cwl_79_50 word79_50 gnd C_wl
Rw80_50 word80_50 word79_50 R_wl
Cwl_80_50 word80_50 gnd C_wl
Rw81_50 word81_50 word80_50 R_wl
Cwl_81_50 word81_50 gnd C_wl
Rw82_50 word82_50 word81_50 R_wl
Cwl_82_50 word82_50 gnd C_wl
Rw83_50 word83_50 word82_50 R_wl
Cwl_83_50 word83_50 gnd C_wl
Rw84_50 word84_50 word83_50 R_wl
Cwl_84_50 word84_50 gnd C_wl
Rw85_50 word85_50 word84_50 R_wl
Cwl_85_50 word85_50 gnd C_wl
Rw86_50 word86_50 word85_50 R_wl
Cwl_86_50 word86_50 gnd C_wl
Rw87_50 word87_50 word86_50 R_wl
Cwl_87_50 word87_50 gnd C_wl
Rw88_50 word88_50 word87_50 R_wl
Cwl_88_50 word88_50 gnd C_wl
Rw89_50 word89_50 word88_50 R_wl
Cwl_89_50 word89_50 gnd C_wl
Rw90_50 word90_50 word89_50 R_wl
Cwl_90_50 word90_50 gnd C_wl
Rw91_50 word91_50 word90_50 R_wl
Cwl_91_50 word91_50 gnd C_wl
Rw92_50 word92_50 word91_50 R_wl
Cwl_92_50 word92_50 gnd C_wl
Rw93_50 word93_50 word92_50 R_wl
Cwl_93_50 word93_50 gnd C_wl
Rw94_50 word94_50 word93_50 R_wl
Cwl_94_50 word94_50 gnd C_wl
Rw95_50 word95_50 word94_50 R_wl
Cwl_95_50 word95_50 gnd C_wl
Rw96_50 word96_50 word95_50 R_wl
Cwl_96_50 word96_50 gnd C_wl
Rw97_50 word97_50 word96_50 R_wl
Cwl_97_50 word97_50 gnd C_wl
Rw98_50 word98_50 word97_50 R_wl
Cwl_98_50 word98_50 gnd C_wl
Rw99_50 word99_50 word98_50 R_wl
Cwl_99_50 word99_50 gnd C_wl
Vwl_51 word_51 0 0
Rw0_51 word_51 word0_51 R_wl
Cwl_0_51 word0_51 gnd C_wl
Rw1_51 word1_51 word0_51 R_wl
Cwl_1_51 word1_51 gnd C_wl
Rw2_51 word2_51 word1_51 R_wl
Cwl_2_51 word2_51 gnd C_wl
Rw3_51 word3_51 word2_51 R_wl
Cwl_3_51 word3_51 gnd C_wl
Rw4_51 word4_51 word3_51 R_wl
Cwl_4_51 word4_51 gnd C_wl
Rw5_51 word5_51 word4_51 R_wl
Cwl_5_51 word5_51 gnd C_wl
Rw6_51 word6_51 word5_51 R_wl
Cwl_6_51 word6_51 gnd C_wl
Rw7_51 word7_51 word6_51 R_wl
Cwl_7_51 word7_51 gnd C_wl
Rw8_51 word8_51 word7_51 R_wl
Cwl_8_51 word8_51 gnd C_wl
Rw9_51 word9_51 word8_51 R_wl
Cwl_9_51 word9_51 gnd C_wl
Rw10_51 word10_51 word9_51 R_wl
Cwl_10_51 word10_51 gnd C_wl
Rw11_51 word11_51 word10_51 R_wl
Cwl_11_51 word11_51 gnd C_wl
Rw12_51 word12_51 word11_51 R_wl
Cwl_12_51 word12_51 gnd C_wl
Rw13_51 word13_51 word12_51 R_wl
Cwl_13_51 word13_51 gnd C_wl
Rw14_51 word14_51 word13_51 R_wl
Cwl_14_51 word14_51 gnd C_wl
Rw15_51 word15_51 word14_51 R_wl
Cwl_15_51 word15_51 gnd C_wl
Rw16_51 word16_51 word15_51 R_wl
Cwl_16_51 word16_51 gnd C_wl
Rw17_51 word17_51 word16_51 R_wl
Cwl_17_51 word17_51 gnd C_wl
Rw18_51 word18_51 word17_51 R_wl
Cwl_18_51 word18_51 gnd C_wl
Rw19_51 word19_51 word18_51 R_wl
Cwl_19_51 word19_51 gnd C_wl
Rw20_51 word20_51 word19_51 R_wl
Cwl_20_51 word20_51 gnd C_wl
Rw21_51 word21_51 word20_51 R_wl
Cwl_21_51 word21_51 gnd C_wl
Rw22_51 word22_51 word21_51 R_wl
Cwl_22_51 word22_51 gnd C_wl
Rw23_51 word23_51 word22_51 R_wl
Cwl_23_51 word23_51 gnd C_wl
Rw24_51 word24_51 word23_51 R_wl
Cwl_24_51 word24_51 gnd C_wl
Rw25_51 word25_51 word24_51 R_wl
Cwl_25_51 word25_51 gnd C_wl
Rw26_51 word26_51 word25_51 R_wl
Cwl_26_51 word26_51 gnd C_wl
Rw27_51 word27_51 word26_51 R_wl
Cwl_27_51 word27_51 gnd C_wl
Rw28_51 word28_51 word27_51 R_wl
Cwl_28_51 word28_51 gnd C_wl
Rw29_51 word29_51 word28_51 R_wl
Cwl_29_51 word29_51 gnd C_wl
Rw30_51 word30_51 word29_51 R_wl
Cwl_30_51 word30_51 gnd C_wl
Rw31_51 word31_51 word30_51 R_wl
Cwl_31_51 word31_51 gnd C_wl
Rw32_51 word32_51 word31_51 R_wl
Cwl_32_51 word32_51 gnd C_wl
Rw33_51 word33_51 word32_51 R_wl
Cwl_33_51 word33_51 gnd C_wl
Rw34_51 word34_51 word33_51 R_wl
Cwl_34_51 word34_51 gnd C_wl
Rw35_51 word35_51 word34_51 R_wl
Cwl_35_51 word35_51 gnd C_wl
Rw36_51 word36_51 word35_51 R_wl
Cwl_36_51 word36_51 gnd C_wl
Rw37_51 word37_51 word36_51 R_wl
Cwl_37_51 word37_51 gnd C_wl
Rw38_51 word38_51 word37_51 R_wl
Cwl_38_51 word38_51 gnd C_wl
Rw39_51 word39_51 word38_51 R_wl
Cwl_39_51 word39_51 gnd C_wl
Rw40_51 word40_51 word39_51 R_wl
Cwl_40_51 word40_51 gnd C_wl
Rw41_51 word41_51 word40_51 R_wl
Cwl_41_51 word41_51 gnd C_wl
Rw42_51 word42_51 word41_51 R_wl
Cwl_42_51 word42_51 gnd C_wl
Rw43_51 word43_51 word42_51 R_wl
Cwl_43_51 word43_51 gnd C_wl
Rw44_51 word44_51 word43_51 R_wl
Cwl_44_51 word44_51 gnd C_wl
Rw45_51 word45_51 word44_51 R_wl
Cwl_45_51 word45_51 gnd C_wl
Rw46_51 word46_51 word45_51 R_wl
Cwl_46_51 word46_51 gnd C_wl
Rw47_51 word47_51 word46_51 R_wl
Cwl_47_51 word47_51 gnd C_wl
Rw48_51 word48_51 word47_51 R_wl
Cwl_48_51 word48_51 gnd C_wl
Rw49_51 word49_51 word48_51 R_wl
Cwl_49_51 word49_51 gnd C_wl
Rw50_51 word50_51 word49_51 R_wl
Cwl_50_51 word50_51 gnd C_wl
Rw51_51 word51_51 word50_51 R_wl
Cwl_51_51 word51_51 gnd C_wl
Rw52_51 word52_51 word51_51 R_wl
Cwl_52_51 word52_51 gnd C_wl
Rw53_51 word53_51 word52_51 R_wl
Cwl_53_51 word53_51 gnd C_wl
Rw54_51 word54_51 word53_51 R_wl
Cwl_54_51 word54_51 gnd C_wl
Rw55_51 word55_51 word54_51 R_wl
Cwl_55_51 word55_51 gnd C_wl
Rw56_51 word56_51 word55_51 R_wl
Cwl_56_51 word56_51 gnd C_wl
Rw57_51 word57_51 word56_51 R_wl
Cwl_57_51 word57_51 gnd C_wl
Rw58_51 word58_51 word57_51 R_wl
Cwl_58_51 word58_51 gnd C_wl
Rw59_51 word59_51 word58_51 R_wl
Cwl_59_51 word59_51 gnd C_wl
Rw60_51 word60_51 word59_51 R_wl
Cwl_60_51 word60_51 gnd C_wl
Rw61_51 word61_51 word60_51 R_wl
Cwl_61_51 word61_51 gnd C_wl
Rw62_51 word62_51 word61_51 R_wl
Cwl_62_51 word62_51 gnd C_wl
Rw63_51 word63_51 word62_51 R_wl
Cwl_63_51 word63_51 gnd C_wl
Rw64_51 word64_51 word63_51 R_wl
Cwl_64_51 word64_51 gnd C_wl
Rw65_51 word65_51 word64_51 R_wl
Cwl_65_51 word65_51 gnd C_wl
Rw66_51 word66_51 word65_51 R_wl
Cwl_66_51 word66_51 gnd C_wl
Rw67_51 word67_51 word66_51 R_wl
Cwl_67_51 word67_51 gnd C_wl
Rw68_51 word68_51 word67_51 R_wl
Cwl_68_51 word68_51 gnd C_wl
Rw69_51 word69_51 word68_51 R_wl
Cwl_69_51 word69_51 gnd C_wl
Rw70_51 word70_51 word69_51 R_wl
Cwl_70_51 word70_51 gnd C_wl
Rw71_51 word71_51 word70_51 R_wl
Cwl_71_51 word71_51 gnd C_wl
Rw72_51 word72_51 word71_51 R_wl
Cwl_72_51 word72_51 gnd C_wl
Rw73_51 word73_51 word72_51 R_wl
Cwl_73_51 word73_51 gnd C_wl
Rw74_51 word74_51 word73_51 R_wl
Cwl_74_51 word74_51 gnd C_wl
Rw75_51 word75_51 word74_51 R_wl
Cwl_75_51 word75_51 gnd C_wl
Rw76_51 word76_51 word75_51 R_wl
Cwl_76_51 word76_51 gnd C_wl
Rw77_51 word77_51 word76_51 R_wl
Cwl_77_51 word77_51 gnd C_wl
Rw78_51 word78_51 word77_51 R_wl
Cwl_78_51 word78_51 gnd C_wl
Rw79_51 word79_51 word78_51 R_wl
Cwl_79_51 word79_51 gnd C_wl
Rw80_51 word80_51 word79_51 R_wl
Cwl_80_51 word80_51 gnd C_wl
Rw81_51 word81_51 word80_51 R_wl
Cwl_81_51 word81_51 gnd C_wl
Rw82_51 word82_51 word81_51 R_wl
Cwl_82_51 word82_51 gnd C_wl
Rw83_51 word83_51 word82_51 R_wl
Cwl_83_51 word83_51 gnd C_wl
Rw84_51 word84_51 word83_51 R_wl
Cwl_84_51 word84_51 gnd C_wl
Rw85_51 word85_51 word84_51 R_wl
Cwl_85_51 word85_51 gnd C_wl
Rw86_51 word86_51 word85_51 R_wl
Cwl_86_51 word86_51 gnd C_wl
Rw87_51 word87_51 word86_51 R_wl
Cwl_87_51 word87_51 gnd C_wl
Rw88_51 word88_51 word87_51 R_wl
Cwl_88_51 word88_51 gnd C_wl
Rw89_51 word89_51 word88_51 R_wl
Cwl_89_51 word89_51 gnd C_wl
Rw90_51 word90_51 word89_51 R_wl
Cwl_90_51 word90_51 gnd C_wl
Rw91_51 word91_51 word90_51 R_wl
Cwl_91_51 word91_51 gnd C_wl
Rw92_51 word92_51 word91_51 R_wl
Cwl_92_51 word92_51 gnd C_wl
Rw93_51 word93_51 word92_51 R_wl
Cwl_93_51 word93_51 gnd C_wl
Rw94_51 word94_51 word93_51 R_wl
Cwl_94_51 word94_51 gnd C_wl
Rw95_51 word95_51 word94_51 R_wl
Cwl_95_51 word95_51 gnd C_wl
Rw96_51 word96_51 word95_51 R_wl
Cwl_96_51 word96_51 gnd C_wl
Rw97_51 word97_51 word96_51 R_wl
Cwl_97_51 word97_51 gnd C_wl
Rw98_51 word98_51 word97_51 R_wl
Cwl_98_51 word98_51 gnd C_wl
Rw99_51 word99_51 word98_51 R_wl
Cwl_99_51 word99_51 gnd C_wl
Vwl_52 word_52 0 0
Rw0_52 word_52 word0_52 R_wl
Cwl_0_52 word0_52 gnd C_wl
Rw1_52 word1_52 word0_52 R_wl
Cwl_1_52 word1_52 gnd C_wl
Rw2_52 word2_52 word1_52 R_wl
Cwl_2_52 word2_52 gnd C_wl
Rw3_52 word3_52 word2_52 R_wl
Cwl_3_52 word3_52 gnd C_wl
Rw4_52 word4_52 word3_52 R_wl
Cwl_4_52 word4_52 gnd C_wl
Rw5_52 word5_52 word4_52 R_wl
Cwl_5_52 word5_52 gnd C_wl
Rw6_52 word6_52 word5_52 R_wl
Cwl_6_52 word6_52 gnd C_wl
Rw7_52 word7_52 word6_52 R_wl
Cwl_7_52 word7_52 gnd C_wl
Rw8_52 word8_52 word7_52 R_wl
Cwl_8_52 word8_52 gnd C_wl
Rw9_52 word9_52 word8_52 R_wl
Cwl_9_52 word9_52 gnd C_wl
Rw10_52 word10_52 word9_52 R_wl
Cwl_10_52 word10_52 gnd C_wl
Rw11_52 word11_52 word10_52 R_wl
Cwl_11_52 word11_52 gnd C_wl
Rw12_52 word12_52 word11_52 R_wl
Cwl_12_52 word12_52 gnd C_wl
Rw13_52 word13_52 word12_52 R_wl
Cwl_13_52 word13_52 gnd C_wl
Rw14_52 word14_52 word13_52 R_wl
Cwl_14_52 word14_52 gnd C_wl
Rw15_52 word15_52 word14_52 R_wl
Cwl_15_52 word15_52 gnd C_wl
Rw16_52 word16_52 word15_52 R_wl
Cwl_16_52 word16_52 gnd C_wl
Rw17_52 word17_52 word16_52 R_wl
Cwl_17_52 word17_52 gnd C_wl
Rw18_52 word18_52 word17_52 R_wl
Cwl_18_52 word18_52 gnd C_wl
Rw19_52 word19_52 word18_52 R_wl
Cwl_19_52 word19_52 gnd C_wl
Rw20_52 word20_52 word19_52 R_wl
Cwl_20_52 word20_52 gnd C_wl
Rw21_52 word21_52 word20_52 R_wl
Cwl_21_52 word21_52 gnd C_wl
Rw22_52 word22_52 word21_52 R_wl
Cwl_22_52 word22_52 gnd C_wl
Rw23_52 word23_52 word22_52 R_wl
Cwl_23_52 word23_52 gnd C_wl
Rw24_52 word24_52 word23_52 R_wl
Cwl_24_52 word24_52 gnd C_wl
Rw25_52 word25_52 word24_52 R_wl
Cwl_25_52 word25_52 gnd C_wl
Rw26_52 word26_52 word25_52 R_wl
Cwl_26_52 word26_52 gnd C_wl
Rw27_52 word27_52 word26_52 R_wl
Cwl_27_52 word27_52 gnd C_wl
Rw28_52 word28_52 word27_52 R_wl
Cwl_28_52 word28_52 gnd C_wl
Rw29_52 word29_52 word28_52 R_wl
Cwl_29_52 word29_52 gnd C_wl
Rw30_52 word30_52 word29_52 R_wl
Cwl_30_52 word30_52 gnd C_wl
Rw31_52 word31_52 word30_52 R_wl
Cwl_31_52 word31_52 gnd C_wl
Rw32_52 word32_52 word31_52 R_wl
Cwl_32_52 word32_52 gnd C_wl
Rw33_52 word33_52 word32_52 R_wl
Cwl_33_52 word33_52 gnd C_wl
Rw34_52 word34_52 word33_52 R_wl
Cwl_34_52 word34_52 gnd C_wl
Rw35_52 word35_52 word34_52 R_wl
Cwl_35_52 word35_52 gnd C_wl
Rw36_52 word36_52 word35_52 R_wl
Cwl_36_52 word36_52 gnd C_wl
Rw37_52 word37_52 word36_52 R_wl
Cwl_37_52 word37_52 gnd C_wl
Rw38_52 word38_52 word37_52 R_wl
Cwl_38_52 word38_52 gnd C_wl
Rw39_52 word39_52 word38_52 R_wl
Cwl_39_52 word39_52 gnd C_wl
Rw40_52 word40_52 word39_52 R_wl
Cwl_40_52 word40_52 gnd C_wl
Rw41_52 word41_52 word40_52 R_wl
Cwl_41_52 word41_52 gnd C_wl
Rw42_52 word42_52 word41_52 R_wl
Cwl_42_52 word42_52 gnd C_wl
Rw43_52 word43_52 word42_52 R_wl
Cwl_43_52 word43_52 gnd C_wl
Rw44_52 word44_52 word43_52 R_wl
Cwl_44_52 word44_52 gnd C_wl
Rw45_52 word45_52 word44_52 R_wl
Cwl_45_52 word45_52 gnd C_wl
Rw46_52 word46_52 word45_52 R_wl
Cwl_46_52 word46_52 gnd C_wl
Rw47_52 word47_52 word46_52 R_wl
Cwl_47_52 word47_52 gnd C_wl
Rw48_52 word48_52 word47_52 R_wl
Cwl_48_52 word48_52 gnd C_wl
Rw49_52 word49_52 word48_52 R_wl
Cwl_49_52 word49_52 gnd C_wl
Rw50_52 word50_52 word49_52 R_wl
Cwl_50_52 word50_52 gnd C_wl
Rw51_52 word51_52 word50_52 R_wl
Cwl_51_52 word51_52 gnd C_wl
Rw52_52 word52_52 word51_52 R_wl
Cwl_52_52 word52_52 gnd C_wl
Rw53_52 word53_52 word52_52 R_wl
Cwl_53_52 word53_52 gnd C_wl
Rw54_52 word54_52 word53_52 R_wl
Cwl_54_52 word54_52 gnd C_wl
Rw55_52 word55_52 word54_52 R_wl
Cwl_55_52 word55_52 gnd C_wl
Rw56_52 word56_52 word55_52 R_wl
Cwl_56_52 word56_52 gnd C_wl
Rw57_52 word57_52 word56_52 R_wl
Cwl_57_52 word57_52 gnd C_wl
Rw58_52 word58_52 word57_52 R_wl
Cwl_58_52 word58_52 gnd C_wl
Rw59_52 word59_52 word58_52 R_wl
Cwl_59_52 word59_52 gnd C_wl
Rw60_52 word60_52 word59_52 R_wl
Cwl_60_52 word60_52 gnd C_wl
Rw61_52 word61_52 word60_52 R_wl
Cwl_61_52 word61_52 gnd C_wl
Rw62_52 word62_52 word61_52 R_wl
Cwl_62_52 word62_52 gnd C_wl
Rw63_52 word63_52 word62_52 R_wl
Cwl_63_52 word63_52 gnd C_wl
Rw64_52 word64_52 word63_52 R_wl
Cwl_64_52 word64_52 gnd C_wl
Rw65_52 word65_52 word64_52 R_wl
Cwl_65_52 word65_52 gnd C_wl
Rw66_52 word66_52 word65_52 R_wl
Cwl_66_52 word66_52 gnd C_wl
Rw67_52 word67_52 word66_52 R_wl
Cwl_67_52 word67_52 gnd C_wl
Rw68_52 word68_52 word67_52 R_wl
Cwl_68_52 word68_52 gnd C_wl
Rw69_52 word69_52 word68_52 R_wl
Cwl_69_52 word69_52 gnd C_wl
Rw70_52 word70_52 word69_52 R_wl
Cwl_70_52 word70_52 gnd C_wl
Rw71_52 word71_52 word70_52 R_wl
Cwl_71_52 word71_52 gnd C_wl
Rw72_52 word72_52 word71_52 R_wl
Cwl_72_52 word72_52 gnd C_wl
Rw73_52 word73_52 word72_52 R_wl
Cwl_73_52 word73_52 gnd C_wl
Rw74_52 word74_52 word73_52 R_wl
Cwl_74_52 word74_52 gnd C_wl
Rw75_52 word75_52 word74_52 R_wl
Cwl_75_52 word75_52 gnd C_wl
Rw76_52 word76_52 word75_52 R_wl
Cwl_76_52 word76_52 gnd C_wl
Rw77_52 word77_52 word76_52 R_wl
Cwl_77_52 word77_52 gnd C_wl
Rw78_52 word78_52 word77_52 R_wl
Cwl_78_52 word78_52 gnd C_wl
Rw79_52 word79_52 word78_52 R_wl
Cwl_79_52 word79_52 gnd C_wl
Rw80_52 word80_52 word79_52 R_wl
Cwl_80_52 word80_52 gnd C_wl
Rw81_52 word81_52 word80_52 R_wl
Cwl_81_52 word81_52 gnd C_wl
Rw82_52 word82_52 word81_52 R_wl
Cwl_82_52 word82_52 gnd C_wl
Rw83_52 word83_52 word82_52 R_wl
Cwl_83_52 word83_52 gnd C_wl
Rw84_52 word84_52 word83_52 R_wl
Cwl_84_52 word84_52 gnd C_wl
Rw85_52 word85_52 word84_52 R_wl
Cwl_85_52 word85_52 gnd C_wl
Rw86_52 word86_52 word85_52 R_wl
Cwl_86_52 word86_52 gnd C_wl
Rw87_52 word87_52 word86_52 R_wl
Cwl_87_52 word87_52 gnd C_wl
Rw88_52 word88_52 word87_52 R_wl
Cwl_88_52 word88_52 gnd C_wl
Rw89_52 word89_52 word88_52 R_wl
Cwl_89_52 word89_52 gnd C_wl
Rw90_52 word90_52 word89_52 R_wl
Cwl_90_52 word90_52 gnd C_wl
Rw91_52 word91_52 word90_52 R_wl
Cwl_91_52 word91_52 gnd C_wl
Rw92_52 word92_52 word91_52 R_wl
Cwl_92_52 word92_52 gnd C_wl
Rw93_52 word93_52 word92_52 R_wl
Cwl_93_52 word93_52 gnd C_wl
Rw94_52 word94_52 word93_52 R_wl
Cwl_94_52 word94_52 gnd C_wl
Rw95_52 word95_52 word94_52 R_wl
Cwl_95_52 word95_52 gnd C_wl
Rw96_52 word96_52 word95_52 R_wl
Cwl_96_52 word96_52 gnd C_wl
Rw97_52 word97_52 word96_52 R_wl
Cwl_97_52 word97_52 gnd C_wl
Rw98_52 word98_52 word97_52 R_wl
Cwl_98_52 word98_52 gnd C_wl
Rw99_52 word99_52 word98_52 R_wl
Cwl_99_52 word99_52 gnd C_wl
Vwl_53 word_53 0 0
Rw0_53 word_53 word0_53 R_wl
Cwl_0_53 word0_53 gnd C_wl
Rw1_53 word1_53 word0_53 R_wl
Cwl_1_53 word1_53 gnd C_wl
Rw2_53 word2_53 word1_53 R_wl
Cwl_2_53 word2_53 gnd C_wl
Rw3_53 word3_53 word2_53 R_wl
Cwl_3_53 word3_53 gnd C_wl
Rw4_53 word4_53 word3_53 R_wl
Cwl_4_53 word4_53 gnd C_wl
Rw5_53 word5_53 word4_53 R_wl
Cwl_5_53 word5_53 gnd C_wl
Rw6_53 word6_53 word5_53 R_wl
Cwl_6_53 word6_53 gnd C_wl
Rw7_53 word7_53 word6_53 R_wl
Cwl_7_53 word7_53 gnd C_wl
Rw8_53 word8_53 word7_53 R_wl
Cwl_8_53 word8_53 gnd C_wl
Rw9_53 word9_53 word8_53 R_wl
Cwl_9_53 word9_53 gnd C_wl
Rw10_53 word10_53 word9_53 R_wl
Cwl_10_53 word10_53 gnd C_wl
Rw11_53 word11_53 word10_53 R_wl
Cwl_11_53 word11_53 gnd C_wl
Rw12_53 word12_53 word11_53 R_wl
Cwl_12_53 word12_53 gnd C_wl
Rw13_53 word13_53 word12_53 R_wl
Cwl_13_53 word13_53 gnd C_wl
Rw14_53 word14_53 word13_53 R_wl
Cwl_14_53 word14_53 gnd C_wl
Rw15_53 word15_53 word14_53 R_wl
Cwl_15_53 word15_53 gnd C_wl
Rw16_53 word16_53 word15_53 R_wl
Cwl_16_53 word16_53 gnd C_wl
Rw17_53 word17_53 word16_53 R_wl
Cwl_17_53 word17_53 gnd C_wl
Rw18_53 word18_53 word17_53 R_wl
Cwl_18_53 word18_53 gnd C_wl
Rw19_53 word19_53 word18_53 R_wl
Cwl_19_53 word19_53 gnd C_wl
Rw20_53 word20_53 word19_53 R_wl
Cwl_20_53 word20_53 gnd C_wl
Rw21_53 word21_53 word20_53 R_wl
Cwl_21_53 word21_53 gnd C_wl
Rw22_53 word22_53 word21_53 R_wl
Cwl_22_53 word22_53 gnd C_wl
Rw23_53 word23_53 word22_53 R_wl
Cwl_23_53 word23_53 gnd C_wl
Rw24_53 word24_53 word23_53 R_wl
Cwl_24_53 word24_53 gnd C_wl
Rw25_53 word25_53 word24_53 R_wl
Cwl_25_53 word25_53 gnd C_wl
Rw26_53 word26_53 word25_53 R_wl
Cwl_26_53 word26_53 gnd C_wl
Rw27_53 word27_53 word26_53 R_wl
Cwl_27_53 word27_53 gnd C_wl
Rw28_53 word28_53 word27_53 R_wl
Cwl_28_53 word28_53 gnd C_wl
Rw29_53 word29_53 word28_53 R_wl
Cwl_29_53 word29_53 gnd C_wl
Rw30_53 word30_53 word29_53 R_wl
Cwl_30_53 word30_53 gnd C_wl
Rw31_53 word31_53 word30_53 R_wl
Cwl_31_53 word31_53 gnd C_wl
Rw32_53 word32_53 word31_53 R_wl
Cwl_32_53 word32_53 gnd C_wl
Rw33_53 word33_53 word32_53 R_wl
Cwl_33_53 word33_53 gnd C_wl
Rw34_53 word34_53 word33_53 R_wl
Cwl_34_53 word34_53 gnd C_wl
Rw35_53 word35_53 word34_53 R_wl
Cwl_35_53 word35_53 gnd C_wl
Rw36_53 word36_53 word35_53 R_wl
Cwl_36_53 word36_53 gnd C_wl
Rw37_53 word37_53 word36_53 R_wl
Cwl_37_53 word37_53 gnd C_wl
Rw38_53 word38_53 word37_53 R_wl
Cwl_38_53 word38_53 gnd C_wl
Rw39_53 word39_53 word38_53 R_wl
Cwl_39_53 word39_53 gnd C_wl
Rw40_53 word40_53 word39_53 R_wl
Cwl_40_53 word40_53 gnd C_wl
Rw41_53 word41_53 word40_53 R_wl
Cwl_41_53 word41_53 gnd C_wl
Rw42_53 word42_53 word41_53 R_wl
Cwl_42_53 word42_53 gnd C_wl
Rw43_53 word43_53 word42_53 R_wl
Cwl_43_53 word43_53 gnd C_wl
Rw44_53 word44_53 word43_53 R_wl
Cwl_44_53 word44_53 gnd C_wl
Rw45_53 word45_53 word44_53 R_wl
Cwl_45_53 word45_53 gnd C_wl
Rw46_53 word46_53 word45_53 R_wl
Cwl_46_53 word46_53 gnd C_wl
Rw47_53 word47_53 word46_53 R_wl
Cwl_47_53 word47_53 gnd C_wl
Rw48_53 word48_53 word47_53 R_wl
Cwl_48_53 word48_53 gnd C_wl
Rw49_53 word49_53 word48_53 R_wl
Cwl_49_53 word49_53 gnd C_wl
Rw50_53 word50_53 word49_53 R_wl
Cwl_50_53 word50_53 gnd C_wl
Rw51_53 word51_53 word50_53 R_wl
Cwl_51_53 word51_53 gnd C_wl
Rw52_53 word52_53 word51_53 R_wl
Cwl_52_53 word52_53 gnd C_wl
Rw53_53 word53_53 word52_53 R_wl
Cwl_53_53 word53_53 gnd C_wl
Rw54_53 word54_53 word53_53 R_wl
Cwl_54_53 word54_53 gnd C_wl
Rw55_53 word55_53 word54_53 R_wl
Cwl_55_53 word55_53 gnd C_wl
Rw56_53 word56_53 word55_53 R_wl
Cwl_56_53 word56_53 gnd C_wl
Rw57_53 word57_53 word56_53 R_wl
Cwl_57_53 word57_53 gnd C_wl
Rw58_53 word58_53 word57_53 R_wl
Cwl_58_53 word58_53 gnd C_wl
Rw59_53 word59_53 word58_53 R_wl
Cwl_59_53 word59_53 gnd C_wl
Rw60_53 word60_53 word59_53 R_wl
Cwl_60_53 word60_53 gnd C_wl
Rw61_53 word61_53 word60_53 R_wl
Cwl_61_53 word61_53 gnd C_wl
Rw62_53 word62_53 word61_53 R_wl
Cwl_62_53 word62_53 gnd C_wl
Rw63_53 word63_53 word62_53 R_wl
Cwl_63_53 word63_53 gnd C_wl
Rw64_53 word64_53 word63_53 R_wl
Cwl_64_53 word64_53 gnd C_wl
Rw65_53 word65_53 word64_53 R_wl
Cwl_65_53 word65_53 gnd C_wl
Rw66_53 word66_53 word65_53 R_wl
Cwl_66_53 word66_53 gnd C_wl
Rw67_53 word67_53 word66_53 R_wl
Cwl_67_53 word67_53 gnd C_wl
Rw68_53 word68_53 word67_53 R_wl
Cwl_68_53 word68_53 gnd C_wl
Rw69_53 word69_53 word68_53 R_wl
Cwl_69_53 word69_53 gnd C_wl
Rw70_53 word70_53 word69_53 R_wl
Cwl_70_53 word70_53 gnd C_wl
Rw71_53 word71_53 word70_53 R_wl
Cwl_71_53 word71_53 gnd C_wl
Rw72_53 word72_53 word71_53 R_wl
Cwl_72_53 word72_53 gnd C_wl
Rw73_53 word73_53 word72_53 R_wl
Cwl_73_53 word73_53 gnd C_wl
Rw74_53 word74_53 word73_53 R_wl
Cwl_74_53 word74_53 gnd C_wl
Rw75_53 word75_53 word74_53 R_wl
Cwl_75_53 word75_53 gnd C_wl
Rw76_53 word76_53 word75_53 R_wl
Cwl_76_53 word76_53 gnd C_wl
Rw77_53 word77_53 word76_53 R_wl
Cwl_77_53 word77_53 gnd C_wl
Rw78_53 word78_53 word77_53 R_wl
Cwl_78_53 word78_53 gnd C_wl
Rw79_53 word79_53 word78_53 R_wl
Cwl_79_53 word79_53 gnd C_wl
Rw80_53 word80_53 word79_53 R_wl
Cwl_80_53 word80_53 gnd C_wl
Rw81_53 word81_53 word80_53 R_wl
Cwl_81_53 word81_53 gnd C_wl
Rw82_53 word82_53 word81_53 R_wl
Cwl_82_53 word82_53 gnd C_wl
Rw83_53 word83_53 word82_53 R_wl
Cwl_83_53 word83_53 gnd C_wl
Rw84_53 word84_53 word83_53 R_wl
Cwl_84_53 word84_53 gnd C_wl
Rw85_53 word85_53 word84_53 R_wl
Cwl_85_53 word85_53 gnd C_wl
Rw86_53 word86_53 word85_53 R_wl
Cwl_86_53 word86_53 gnd C_wl
Rw87_53 word87_53 word86_53 R_wl
Cwl_87_53 word87_53 gnd C_wl
Rw88_53 word88_53 word87_53 R_wl
Cwl_88_53 word88_53 gnd C_wl
Rw89_53 word89_53 word88_53 R_wl
Cwl_89_53 word89_53 gnd C_wl
Rw90_53 word90_53 word89_53 R_wl
Cwl_90_53 word90_53 gnd C_wl
Rw91_53 word91_53 word90_53 R_wl
Cwl_91_53 word91_53 gnd C_wl
Rw92_53 word92_53 word91_53 R_wl
Cwl_92_53 word92_53 gnd C_wl
Rw93_53 word93_53 word92_53 R_wl
Cwl_93_53 word93_53 gnd C_wl
Rw94_53 word94_53 word93_53 R_wl
Cwl_94_53 word94_53 gnd C_wl
Rw95_53 word95_53 word94_53 R_wl
Cwl_95_53 word95_53 gnd C_wl
Rw96_53 word96_53 word95_53 R_wl
Cwl_96_53 word96_53 gnd C_wl
Rw97_53 word97_53 word96_53 R_wl
Cwl_97_53 word97_53 gnd C_wl
Rw98_53 word98_53 word97_53 R_wl
Cwl_98_53 word98_53 gnd C_wl
Rw99_53 word99_53 word98_53 R_wl
Cwl_99_53 word99_53 gnd C_wl
Vwl_54 word_54 0 0
Rw0_54 word_54 word0_54 R_wl
Cwl_0_54 word0_54 gnd C_wl
Rw1_54 word1_54 word0_54 R_wl
Cwl_1_54 word1_54 gnd C_wl
Rw2_54 word2_54 word1_54 R_wl
Cwl_2_54 word2_54 gnd C_wl
Rw3_54 word3_54 word2_54 R_wl
Cwl_3_54 word3_54 gnd C_wl
Rw4_54 word4_54 word3_54 R_wl
Cwl_4_54 word4_54 gnd C_wl
Rw5_54 word5_54 word4_54 R_wl
Cwl_5_54 word5_54 gnd C_wl
Rw6_54 word6_54 word5_54 R_wl
Cwl_6_54 word6_54 gnd C_wl
Rw7_54 word7_54 word6_54 R_wl
Cwl_7_54 word7_54 gnd C_wl
Rw8_54 word8_54 word7_54 R_wl
Cwl_8_54 word8_54 gnd C_wl
Rw9_54 word9_54 word8_54 R_wl
Cwl_9_54 word9_54 gnd C_wl
Rw10_54 word10_54 word9_54 R_wl
Cwl_10_54 word10_54 gnd C_wl
Rw11_54 word11_54 word10_54 R_wl
Cwl_11_54 word11_54 gnd C_wl
Rw12_54 word12_54 word11_54 R_wl
Cwl_12_54 word12_54 gnd C_wl
Rw13_54 word13_54 word12_54 R_wl
Cwl_13_54 word13_54 gnd C_wl
Rw14_54 word14_54 word13_54 R_wl
Cwl_14_54 word14_54 gnd C_wl
Rw15_54 word15_54 word14_54 R_wl
Cwl_15_54 word15_54 gnd C_wl
Rw16_54 word16_54 word15_54 R_wl
Cwl_16_54 word16_54 gnd C_wl
Rw17_54 word17_54 word16_54 R_wl
Cwl_17_54 word17_54 gnd C_wl
Rw18_54 word18_54 word17_54 R_wl
Cwl_18_54 word18_54 gnd C_wl
Rw19_54 word19_54 word18_54 R_wl
Cwl_19_54 word19_54 gnd C_wl
Rw20_54 word20_54 word19_54 R_wl
Cwl_20_54 word20_54 gnd C_wl
Rw21_54 word21_54 word20_54 R_wl
Cwl_21_54 word21_54 gnd C_wl
Rw22_54 word22_54 word21_54 R_wl
Cwl_22_54 word22_54 gnd C_wl
Rw23_54 word23_54 word22_54 R_wl
Cwl_23_54 word23_54 gnd C_wl
Rw24_54 word24_54 word23_54 R_wl
Cwl_24_54 word24_54 gnd C_wl
Rw25_54 word25_54 word24_54 R_wl
Cwl_25_54 word25_54 gnd C_wl
Rw26_54 word26_54 word25_54 R_wl
Cwl_26_54 word26_54 gnd C_wl
Rw27_54 word27_54 word26_54 R_wl
Cwl_27_54 word27_54 gnd C_wl
Rw28_54 word28_54 word27_54 R_wl
Cwl_28_54 word28_54 gnd C_wl
Rw29_54 word29_54 word28_54 R_wl
Cwl_29_54 word29_54 gnd C_wl
Rw30_54 word30_54 word29_54 R_wl
Cwl_30_54 word30_54 gnd C_wl
Rw31_54 word31_54 word30_54 R_wl
Cwl_31_54 word31_54 gnd C_wl
Rw32_54 word32_54 word31_54 R_wl
Cwl_32_54 word32_54 gnd C_wl
Rw33_54 word33_54 word32_54 R_wl
Cwl_33_54 word33_54 gnd C_wl
Rw34_54 word34_54 word33_54 R_wl
Cwl_34_54 word34_54 gnd C_wl
Rw35_54 word35_54 word34_54 R_wl
Cwl_35_54 word35_54 gnd C_wl
Rw36_54 word36_54 word35_54 R_wl
Cwl_36_54 word36_54 gnd C_wl
Rw37_54 word37_54 word36_54 R_wl
Cwl_37_54 word37_54 gnd C_wl
Rw38_54 word38_54 word37_54 R_wl
Cwl_38_54 word38_54 gnd C_wl
Rw39_54 word39_54 word38_54 R_wl
Cwl_39_54 word39_54 gnd C_wl
Rw40_54 word40_54 word39_54 R_wl
Cwl_40_54 word40_54 gnd C_wl
Rw41_54 word41_54 word40_54 R_wl
Cwl_41_54 word41_54 gnd C_wl
Rw42_54 word42_54 word41_54 R_wl
Cwl_42_54 word42_54 gnd C_wl
Rw43_54 word43_54 word42_54 R_wl
Cwl_43_54 word43_54 gnd C_wl
Rw44_54 word44_54 word43_54 R_wl
Cwl_44_54 word44_54 gnd C_wl
Rw45_54 word45_54 word44_54 R_wl
Cwl_45_54 word45_54 gnd C_wl
Rw46_54 word46_54 word45_54 R_wl
Cwl_46_54 word46_54 gnd C_wl
Rw47_54 word47_54 word46_54 R_wl
Cwl_47_54 word47_54 gnd C_wl
Rw48_54 word48_54 word47_54 R_wl
Cwl_48_54 word48_54 gnd C_wl
Rw49_54 word49_54 word48_54 R_wl
Cwl_49_54 word49_54 gnd C_wl
Rw50_54 word50_54 word49_54 R_wl
Cwl_50_54 word50_54 gnd C_wl
Rw51_54 word51_54 word50_54 R_wl
Cwl_51_54 word51_54 gnd C_wl
Rw52_54 word52_54 word51_54 R_wl
Cwl_52_54 word52_54 gnd C_wl
Rw53_54 word53_54 word52_54 R_wl
Cwl_53_54 word53_54 gnd C_wl
Rw54_54 word54_54 word53_54 R_wl
Cwl_54_54 word54_54 gnd C_wl
Rw55_54 word55_54 word54_54 R_wl
Cwl_55_54 word55_54 gnd C_wl
Rw56_54 word56_54 word55_54 R_wl
Cwl_56_54 word56_54 gnd C_wl
Rw57_54 word57_54 word56_54 R_wl
Cwl_57_54 word57_54 gnd C_wl
Rw58_54 word58_54 word57_54 R_wl
Cwl_58_54 word58_54 gnd C_wl
Rw59_54 word59_54 word58_54 R_wl
Cwl_59_54 word59_54 gnd C_wl
Rw60_54 word60_54 word59_54 R_wl
Cwl_60_54 word60_54 gnd C_wl
Rw61_54 word61_54 word60_54 R_wl
Cwl_61_54 word61_54 gnd C_wl
Rw62_54 word62_54 word61_54 R_wl
Cwl_62_54 word62_54 gnd C_wl
Rw63_54 word63_54 word62_54 R_wl
Cwl_63_54 word63_54 gnd C_wl
Rw64_54 word64_54 word63_54 R_wl
Cwl_64_54 word64_54 gnd C_wl
Rw65_54 word65_54 word64_54 R_wl
Cwl_65_54 word65_54 gnd C_wl
Rw66_54 word66_54 word65_54 R_wl
Cwl_66_54 word66_54 gnd C_wl
Rw67_54 word67_54 word66_54 R_wl
Cwl_67_54 word67_54 gnd C_wl
Rw68_54 word68_54 word67_54 R_wl
Cwl_68_54 word68_54 gnd C_wl
Rw69_54 word69_54 word68_54 R_wl
Cwl_69_54 word69_54 gnd C_wl
Rw70_54 word70_54 word69_54 R_wl
Cwl_70_54 word70_54 gnd C_wl
Rw71_54 word71_54 word70_54 R_wl
Cwl_71_54 word71_54 gnd C_wl
Rw72_54 word72_54 word71_54 R_wl
Cwl_72_54 word72_54 gnd C_wl
Rw73_54 word73_54 word72_54 R_wl
Cwl_73_54 word73_54 gnd C_wl
Rw74_54 word74_54 word73_54 R_wl
Cwl_74_54 word74_54 gnd C_wl
Rw75_54 word75_54 word74_54 R_wl
Cwl_75_54 word75_54 gnd C_wl
Rw76_54 word76_54 word75_54 R_wl
Cwl_76_54 word76_54 gnd C_wl
Rw77_54 word77_54 word76_54 R_wl
Cwl_77_54 word77_54 gnd C_wl
Rw78_54 word78_54 word77_54 R_wl
Cwl_78_54 word78_54 gnd C_wl
Rw79_54 word79_54 word78_54 R_wl
Cwl_79_54 word79_54 gnd C_wl
Rw80_54 word80_54 word79_54 R_wl
Cwl_80_54 word80_54 gnd C_wl
Rw81_54 word81_54 word80_54 R_wl
Cwl_81_54 word81_54 gnd C_wl
Rw82_54 word82_54 word81_54 R_wl
Cwl_82_54 word82_54 gnd C_wl
Rw83_54 word83_54 word82_54 R_wl
Cwl_83_54 word83_54 gnd C_wl
Rw84_54 word84_54 word83_54 R_wl
Cwl_84_54 word84_54 gnd C_wl
Rw85_54 word85_54 word84_54 R_wl
Cwl_85_54 word85_54 gnd C_wl
Rw86_54 word86_54 word85_54 R_wl
Cwl_86_54 word86_54 gnd C_wl
Rw87_54 word87_54 word86_54 R_wl
Cwl_87_54 word87_54 gnd C_wl
Rw88_54 word88_54 word87_54 R_wl
Cwl_88_54 word88_54 gnd C_wl
Rw89_54 word89_54 word88_54 R_wl
Cwl_89_54 word89_54 gnd C_wl
Rw90_54 word90_54 word89_54 R_wl
Cwl_90_54 word90_54 gnd C_wl
Rw91_54 word91_54 word90_54 R_wl
Cwl_91_54 word91_54 gnd C_wl
Rw92_54 word92_54 word91_54 R_wl
Cwl_92_54 word92_54 gnd C_wl
Rw93_54 word93_54 word92_54 R_wl
Cwl_93_54 word93_54 gnd C_wl
Rw94_54 word94_54 word93_54 R_wl
Cwl_94_54 word94_54 gnd C_wl
Rw95_54 word95_54 word94_54 R_wl
Cwl_95_54 word95_54 gnd C_wl
Rw96_54 word96_54 word95_54 R_wl
Cwl_96_54 word96_54 gnd C_wl
Rw97_54 word97_54 word96_54 R_wl
Cwl_97_54 word97_54 gnd C_wl
Rw98_54 word98_54 word97_54 R_wl
Cwl_98_54 word98_54 gnd C_wl
Rw99_54 word99_54 word98_54 R_wl
Cwl_99_54 word99_54 gnd C_wl
Vwl_55 word_55 0 0
Rw0_55 word_55 word0_55 R_wl
Cwl_0_55 word0_55 gnd C_wl
Rw1_55 word1_55 word0_55 R_wl
Cwl_1_55 word1_55 gnd C_wl
Rw2_55 word2_55 word1_55 R_wl
Cwl_2_55 word2_55 gnd C_wl
Rw3_55 word3_55 word2_55 R_wl
Cwl_3_55 word3_55 gnd C_wl
Rw4_55 word4_55 word3_55 R_wl
Cwl_4_55 word4_55 gnd C_wl
Rw5_55 word5_55 word4_55 R_wl
Cwl_5_55 word5_55 gnd C_wl
Rw6_55 word6_55 word5_55 R_wl
Cwl_6_55 word6_55 gnd C_wl
Rw7_55 word7_55 word6_55 R_wl
Cwl_7_55 word7_55 gnd C_wl
Rw8_55 word8_55 word7_55 R_wl
Cwl_8_55 word8_55 gnd C_wl
Rw9_55 word9_55 word8_55 R_wl
Cwl_9_55 word9_55 gnd C_wl
Rw10_55 word10_55 word9_55 R_wl
Cwl_10_55 word10_55 gnd C_wl
Rw11_55 word11_55 word10_55 R_wl
Cwl_11_55 word11_55 gnd C_wl
Rw12_55 word12_55 word11_55 R_wl
Cwl_12_55 word12_55 gnd C_wl
Rw13_55 word13_55 word12_55 R_wl
Cwl_13_55 word13_55 gnd C_wl
Rw14_55 word14_55 word13_55 R_wl
Cwl_14_55 word14_55 gnd C_wl
Rw15_55 word15_55 word14_55 R_wl
Cwl_15_55 word15_55 gnd C_wl
Rw16_55 word16_55 word15_55 R_wl
Cwl_16_55 word16_55 gnd C_wl
Rw17_55 word17_55 word16_55 R_wl
Cwl_17_55 word17_55 gnd C_wl
Rw18_55 word18_55 word17_55 R_wl
Cwl_18_55 word18_55 gnd C_wl
Rw19_55 word19_55 word18_55 R_wl
Cwl_19_55 word19_55 gnd C_wl
Rw20_55 word20_55 word19_55 R_wl
Cwl_20_55 word20_55 gnd C_wl
Rw21_55 word21_55 word20_55 R_wl
Cwl_21_55 word21_55 gnd C_wl
Rw22_55 word22_55 word21_55 R_wl
Cwl_22_55 word22_55 gnd C_wl
Rw23_55 word23_55 word22_55 R_wl
Cwl_23_55 word23_55 gnd C_wl
Rw24_55 word24_55 word23_55 R_wl
Cwl_24_55 word24_55 gnd C_wl
Rw25_55 word25_55 word24_55 R_wl
Cwl_25_55 word25_55 gnd C_wl
Rw26_55 word26_55 word25_55 R_wl
Cwl_26_55 word26_55 gnd C_wl
Rw27_55 word27_55 word26_55 R_wl
Cwl_27_55 word27_55 gnd C_wl
Rw28_55 word28_55 word27_55 R_wl
Cwl_28_55 word28_55 gnd C_wl
Rw29_55 word29_55 word28_55 R_wl
Cwl_29_55 word29_55 gnd C_wl
Rw30_55 word30_55 word29_55 R_wl
Cwl_30_55 word30_55 gnd C_wl
Rw31_55 word31_55 word30_55 R_wl
Cwl_31_55 word31_55 gnd C_wl
Rw32_55 word32_55 word31_55 R_wl
Cwl_32_55 word32_55 gnd C_wl
Rw33_55 word33_55 word32_55 R_wl
Cwl_33_55 word33_55 gnd C_wl
Rw34_55 word34_55 word33_55 R_wl
Cwl_34_55 word34_55 gnd C_wl
Rw35_55 word35_55 word34_55 R_wl
Cwl_35_55 word35_55 gnd C_wl
Rw36_55 word36_55 word35_55 R_wl
Cwl_36_55 word36_55 gnd C_wl
Rw37_55 word37_55 word36_55 R_wl
Cwl_37_55 word37_55 gnd C_wl
Rw38_55 word38_55 word37_55 R_wl
Cwl_38_55 word38_55 gnd C_wl
Rw39_55 word39_55 word38_55 R_wl
Cwl_39_55 word39_55 gnd C_wl
Rw40_55 word40_55 word39_55 R_wl
Cwl_40_55 word40_55 gnd C_wl
Rw41_55 word41_55 word40_55 R_wl
Cwl_41_55 word41_55 gnd C_wl
Rw42_55 word42_55 word41_55 R_wl
Cwl_42_55 word42_55 gnd C_wl
Rw43_55 word43_55 word42_55 R_wl
Cwl_43_55 word43_55 gnd C_wl
Rw44_55 word44_55 word43_55 R_wl
Cwl_44_55 word44_55 gnd C_wl
Rw45_55 word45_55 word44_55 R_wl
Cwl_45_55 word45_55 gnd C_wl
Rw46_55 word46_55 word45_55 R_wl
Cwl_46_55 word46_55 gnd C_wl
Rw47_55 word47_55 word46_55 R_wl
Cwl_47_55 word47_55 gnd C_wl
Rw48_55 word48_55 word47_55 R_wl
Cwl_48_55 word48_55 gnd C_wl
Rw49_55 word49_55 word48_55 R_wl
Cwl_49_55 word49_55 gnd C_wl
Rw50_55 word50_55 word49_55 R_wl
Cwl_50_55 word50_55 gnd C_wl
Rw51_55 word51_55 word50_55 R_wl
Cwl_51_55 word51_55 gnd C_wl
Rw52_55 word52_55 word51_55 R_wl
Cwl_52_55 word52_55 gnd C_wl
Rw53_55 word53_55 word52_55 R_wl
Cwl_53_55 word53_55 gnd C_wl
Rw54_55 word54_55 word53_55 R_wl
Cwl_54_55 word54_55 gnd C_wl
Rw55_55 word55_55 word54_55 R_wl
Cwl_55_55 word55_55 gnd C_wl
Rw56_55 word56_55 word55_55 R_wl
Cwl_56_55 word56_55 gnd C_wl
Rw57_55 word57_55 word56_55 R_wl
Cwl_57_55 word57_55 gnd C_wl
Rw58_55 word58_55 word57_55 R_wl
Cwl_58_55 word58_55 gnd C_wl
Rw59_55 word59_55 word58_55 R_wl
Cwl_59_55 word59_55 gnd C_wl
Rw60_55 word60_55 word59_55 R_wl
Cwl_60_55 word60_55 gnd C_wl
Rw61_55 word61_55 word60_55 R_wl
Cwl_61_55 word61_55 gnd C_wl
Rw62_55 word62_55 word61_55 R_wl
Cwl_62_55 word62_55 gnd C_wl
Rw63_55 word63_55 word62_55 R_wl
Cwl_63_55 word63_55 gnd C_wl
Rw64_55 word64_55 word63_55 R_wl
Cwl_64_55 word64_55 gnd C_wl
Rw65_55 word65_55 word64_55 R_wl
Cwl_65_55 word65_55 gnd C_wl
Rw66_55 word66_55 word65_55 R_wl
Cwl_66_55 word66_55 gnd C_wl
Rw67_55 word67_55 word66_55 R_wl
Cwl_67_55 word67_55 gnd C_wl
Rw68_55 word68_55 word67_55 R_wl
Cwl_68_55 word68_55 gnd C_wl
Rw69_55 word69_55 word68_55 R_wl
Cwl_69_55 word69_55 gnd C_wl
Rw70_55 word70_55 word69_55 R_wl
Cwl_70_55 word70_55 gnd C_wl
Rw71_55 word71_55 word70_55 R_wl
Cwl_71_55 word71_55 gnd C_wl
Rw72_55 word72_55 word71_55 R_wl
Cwl_72_55 word72_55 gnd C_wl
Rw73_55 word73_55 word72_55 R_wl
Cwl_73_55 word73_55 gnd C_wl
Rw74_55 word74_55 word73_55 R_wl
Cwl_74_55 word74_55 gnd C_wl
Rw75_55 word75_55 word74_55 R_wl
Cwl_75_55 word75_55 gnd C_wl
Rw76_55 word76_55 word75_55 R_wl
Cwl_76_55 word76_55 gnd C_wl
Rw77_55 word77_55 word76_55 R_wl
Cwl_77_55 word77_55 gnd C_wl
Rw78_55 word78_55 word77_55 R_wl
Cwl_78_55 word78_55 gnd C_wl
Rw79_55 word79_55 word78_55 R_wl
Cwl_79_55 word79_55 gnd C_wl
Rw80_55 word80_55 word79_55 R_wl
Cwl_80_55 word80_55 gnd C_wl
Rw81_55 word81_55 word80_55 R_wl
Cwl_81_55 word81_55 gnd C_wl
Rw82_55 word82_55 word81_55 R_wl
Cwl_82_55 word82_55 gnd C_wl
Rw83_55 word83_55 word82_55 R_wl
Cwl_83_55 word83_55 gnd C_wl
Rw84_55 word84_55 word83_55 R_wl
Cwl_84_55 word84_55 gnd C_wl
Rw85_55 word85_55 word84_55 R_wl
Cwl_85_55 word85_55 gnd C_wl
Rw86_55 word86_55 word85_55 R_wl
Cwl_86_55 word86_55 gnd C_wl
Rw87_55 word87_55 word86_55 R_wl
Cwl_87_55 word87_55 gnd C_wl
Rw88_55 word88_55 word87_55 R_wl
Cwl_88_55 word88_55 gnd C_wl
Rw89_55 word89_55 word88_55 R_wl
Cwl_89_55 word89_55 gnd C_wl
Rw90_55 word90_55 word89_55 R_wl
Cwl_90_55 word90_55 gnd C_wl
Rw91_55 word91_55 word90_55 R_wl
Cwl_91_55 word91_55 gnd C_wl
Rw92_55 word92_55 word91_55 R_wl
Cwl_92_55 word92_55 gnd C_wl
Rw93_55 word93_55 word92_55 R_wl
Cwl_93_55 word93_55 gnd C_wl
Rw94_55 word94_55 word93_55 R_wl
Cwl_94_55 word94_55 gnd C_wl
Rw95_55 word95_55 word94_55 R_wl
Cwl_95_55 word95_55 gnd C_wl
Rw96_55 word96_55 word95_55 R_wl
Cwl_96_55 word96_55 gnd C_wl
Rw97_55 word97_55 word96_55 R_wl
Cwl_97_55 word97_55 gnd C_wl
Rw98_55 word98_55 word97_55 R_wl
Cwl_98_55 word98_55 gnd C_wl
Rw99_55 word99_55 word98_55 R_wl
Cwl_99_55 word99_55 gnd C_wl
Vwl_56 word_56 0 0
Rw0_56 word_56 word0_56 R_wl
Cwl_0_56 word0_56 gnd C_wl
Rw1_56 word1_56 word0_56 R_wl
Cwl_1_56 word1_56 gnd C_wl
Rw2_56 word2_56 word1_56 R_wl
Cwl_2_56 word2_56 gnd C_wl
Rw3_56 word3_56 word2_56 R_wl
Cwl_3_56 word3_56 gnd C_wl
Rw4_56 word4_56 word3_56 R_wl
Cwl_4_56 word4_56 gnd C_wl
Rw5_56 word5_56 word4_56 R_wl
Cwl_5_56 word5_56 gnd C_wl
Rw6_56 word6_56 word5_56 R_wl
Cwl_6_56 word6_56 gnd C_wl
Rw7_56 word7_56 word6_56 R_wl
Cwl_7_56 word7_56 gnd C_wl
Rw8_56 word8_56 word7_56 R_wl
Cwl_8_56 word8_56 gnd C_wl
Rw9_56 word9_56 word8_56 R_wl
Cwl_9_56 word9_56 gnd C_wl
Rw10_56 word10_56 word9_56 R_wl
Cwl_10_56 word10_56 gnd C_wl
Rw11_56 word11_56 word10_56 R_wl
Cwl_11_56 word11_56 gnd C_wl
Rw12_56 word12_56 word11_56 R_wl
Cwl_12_56 word12_56 gnd C_wl
Rw13_56 word13_56 word12_56 R_wl
Cwl_13_56 word13_56 gnd C_wl
Rw14_56 word14_56 word13_56 R_wl
Cwl_14_56 word14_56 gnd C_wl
Rw15_56 word15_56 word14_56 R_wl
Cwl_15_56 word15_56 gnd C_wl
Rw16_56 word16_56 word15_56 R_wl
Cwl_16_56 word16_56 gnd C_wl
Rw17_56 word17_56 word16_56 R_wl
Cwl_17_56 word17_56 gnd C_wl
Rw18_56 word18_56 word17_56 R_wl
Cwl_18_56 word18_56 gnd C_wl
Rw19_56 word19_56 word18_56 R_wl
Cwl_19_56 word19_56 gnd C_wl
Rw20_56 word20_56 word19_56 R_wl
Cwl_20_56 word20_56 gnd C_wl
Rw21_56 word21_56 word20_56 R_wl
Cwl_21_56 word21_56 gnd C_wl
Rw22_56 word22_56 word21_56 R_wl
Cwl_22_56 word22_56 gnd C_wl
Rw23_56 word23_56 word22_56 R_wl
Cwl_23_56 word23_56 gnd C_wl
Rw24_56 word24_56 word23_56 R_wl
Cwl_24_56 word24_56 gnd C_wl
Rw25_56 word25_56 word24_56 R_wl
Cwl_25_56 word25_56 gnd C_wl
Rw26_56 word26_56 word25_56 R_wl
Cwl_26_56 word26_56 gnd C_wl
Rw27_56 word27_56 word26_56 R_wl
Cwl_27_56 word27_56 gnd C_wl
Rw28_56 word28_56 word27_56 R_wl
Cwl_28_56 word28_56 gnd C_wl
Rw29_56 word29_56 word28_56 R_wl
Cwl_29_56 word29_56 gnd C_wl
Rw30_56 word30_56 word29_56 R_wl
Cwl_30_56 word30_56 gnd C_wl
Rw31_56 word31_56 word30_56 R_wl
Cwl_31_56 word31_56 gnd C_wl
Rw32_56 word32_56 word31_56 R_wl
Cwl_32_56 word32_56 gnd C_wl
Rw33_56 word33_56 word32_56 R_wl
Cwl_33_56 word33_56 gnd C_wl
Rw34_56 word34_56 word33_56 R_wl
Cwl_34_56 word34_56 gnd C_wl
Rw35_56 word35_56 word34_56 R_wl
Cwl_35_56 word35_56 gnd C_wl
Rw36_56 word36_56 word35_56 R_wl
Cwl_36_56 word36_56 gnd C_wl
Rw37_56 word37_56 word36_56 R_wl
Cwl_37_56 word37_56 gnd C_wl
Rw38_56 word38_56 word37_56 R_wl
Cwl_38_56 word38_56 gnd C_wl
Rw39_56 word39_56 word38_56 R_wl
Cwl_39_56 word39_56 gnd C_wl
Rw40_56 word40_56 word39_56 R_wl
Cwl_40_56 word40_56 gnd C_wl
Rw41_56 word41_56 word40_56 R_wl
Cwl_41_56 word41_56 gnd C_wl
Rw42_56 word42_56 word41_56 R_wl
Cwl_42_56 word42_56 gnd C_wl
Rw43_56 word43_56 word42_56 R_wl
Cwl_43_56 word43_56 gnd C_wl
Rw44_56 word44_56 word43_56 R_wl
Cwl_44_56 word44_56 gnd C_wl
Rw45_56 word45_56 word44_56 R_wl
Cwl_45_56 word45_56 gnd C_wl
Rw46_56 word46_56 word45_56 R_wl
Cwl_46_56 word46_56 gnd C_wl
Rw47_56 word47_56 word46_56 R_wl
Cwl_47_56 word47_56 gnd C_wl
Rw48_56 word48_56 word47_56 R_wl
Cwl_48_56 word48_56 gnd C_wl
Rw49_56 word49_56 word48_56 R_wl
Cwl_49_56 word49_56 gnd C_wl
Rw50_56 word50_56 word49_56 R_wl
Cwl_50_56 word50_56 gnd C_wl
Rw51_56 word51_56 word50_56 R_wl
Cwl_51_56 word51_56 gnd C_wl
Rw52_56 word52_56 word51_56 R_wl
Cwl_52_56 word52_56 gnd C_wl
Rw53_56 word53_56 word52_56 R_wl
Cwl_53_56 word53_56 gnd C_wl
Rw54_56 word54_56 word53_56 R_wl
Cwl_54_56 word54_56 gnd C_wl
Rw55_56 word55_56 word54_56 R_wl
Cwl_55_56 word55_56 gnd C_wl
Rw56_56 word56_56 word55_56 R_wl
Cwl_56_56 word56_56 gnd C_wl
Rw57_56 word57_56 word56_56 R_wl
Cwl_57_56 word57_56 gnd C_wl
Rw58_56 word58_56 word57_56 R_wl
Cwl_58_56 word58_56 gnd C_wl
Rw59_56 word59_56 word58_56 R_wl
Cwl_59_56 word59_56 gnd C_wl
Rw60_56 word60_56 word59_56 R_wl
Cwl_60_56 word60_56 gnd C_wl
Rw61_56 word61_56 word60_56 R_wl
Cwl_61_56 word61_56 gnd C_wl
Rw62_56 word62_56 word61_56 R_wl
Cwl_62_56 word62_56 gnd C_wl
Rw63_56 word63_56 word62_56 R_wl
Cwl_63_56 word63_56 gnd C_wl
Rw64_56 word64_56 word63_56 R_wl
Cwl_64_56 word64_56 gnd C_wl
Rw65_56 word65_56 word64_56 R_wl
Cwl_65_56 word65_56 gnd C_wl
Rw66_56 word66_56 word65_56 R_wl
Cwl_66_56 word66_56 gnd C_wl
Rw67_56 word67_56 word66_56 R_wl
Cwl_67_56 word67_56 gnd C_wl
Rw68_56 word68_56 word67_56 R_wl
Cwl_68_56 word68_56 gnd C_wl
Rw69_56 word69_56 word68_56 R_wl
Cwl_69_56 word69_56 gnd C_wl
Rw70_56 word70_56 word69_56 R_wl
Cwl_70_56 word70_56 gnd C_wl
Rw71_56 word71_56 word70_56 R_wl
Cwl_71_56 word71_56 gnd C_wl
Rw72_56 word72_56 word71_56 R_wl
Cwl_72_56 word72_56 gnd C_wl
Rw73_56 word73_56 word72_56 R_wl
Cwl_73_56 word73_56 gnd C_wl
Rw74_56 word74_56 word73_56 R_wl
Cwl_74_56 word74_56 gnd C_wl
Rw75_56 word75_56 word74_56 R_wl
Cwl_75_56 word75_56 gnd C_wl
Rw76_56 word76_56 word75_56 R_wl
Cwl_76_56 word76_56 gnd C_wl
Rw77_56 word77_56 word76_56 R_wl
Cwl_77_56 word77_56 gnd C_wl
Rw78_56 word78_56 word77_56 R_wl
Cwl_78_56 word78_56 gnd C_wl
Rw79_56 word79_56 word78_56 R_wl
Cwl_79_56 word79_56 gnd C_wl
Rw80_56 word80_56 word79_56 R_wl
Cwl_80_56 word80_56 gnd C_wl
Rw81_56 word81_56 word80_56 R_wl
Cwl_81_56 word81_56 gnd C_wl
Rw82_56 word82_56 word81_56 R_wl
Cwl_82_56 word82_56 gnd C_wl
Rw83_56 word83_56 word82_56 R_wl
Cwl_83_56 word83_56 gnd C_wl
Rw84_56 word84_56 word83_56 R_wl
Cwl_84_56 word84_56 gnd C_wl
Rw85_56 word85_56 word84_56 R_wl
Cwl_85_56 word85_56 gnd C_wl
Rw86_56 word86_56 word85_56 R_wl
Cwl_86_56 word86_56 gnd C_wl
Rw87_56 word87_56 word86_56 R_wl
Cwl_87_56 word87_56 gnd C_wl
Rw88_56 word88_56 word87_56 R_wl
Cwl_88_56 word88_56 gnd C_wl
Rw89_56 word89_56 word88_56 R_wl
Cwl_89_56 word89_56 gnd C_wl
Rw90_56 word90_56 word89_56 R_wl
Cwl_90_56 word90_56 gnd C_wl
Rw91_56 word91_56 word90_56 R_wl
Cwl_91_56 word91_56 gnd C_wl
Rw92_56 word92_56 word91_56 R_wl
Cwl_92_56 word92_56 gnd C_wl
Rw93_56 word93_56 word92_56 R_wl
Cwl_93_56 word93_56 gnd C_wl
Rw94_56 word94_56 word93_56 R_wl
Cwl_94_56 word94_56 gnd C_wl
Rw95_56 word95_56 word94_56 R_wl
Cwl_95_56 word95_56 gnd C_wl
Rw96_56 word96_56 word95_56 R_wl
Cwl_96_56 word96_56 gnd C_wl
Rw97_56 word97_56 word96_56 R_wl
Cwl_97_56 word97_56 gnd C_wl
Rw98_56 word98_56 word97_56 R_wl
Cwl_98_56 word98_56 gnd C_wl
Rw99_56 word99_56 word98_56 R_wl
Cwl_99_56 word99_56 gnd C_wl
Vwl_57 word_57 0 0
Rw0_57 word_57 word0_57 R_wl
Cwl_0_57 word0_57 gnd C_wl
Rw1_57 word1_57 word0_57 R_wl
Cwl_1_57 word1_57 gnd C_wl
Rw2_57 word2_57 word1_57 R_wl
Cwl_2_57 word2_57 gnd C_wl
Rw3_57 word3_57 word2_57 R_wl
Cwl_3_57 word3_57 gnd C_wl
Rw4_57 word4_57 word3_57 R_wl
Cwl_4_57 word4_57 gnd C_wl
Rw5_57 word5_57 word4_57 R_wl
Cwl_5_57 word5_57 gnd C_wl
Rw6_57 word6_57 word5_57 R_wl
Cwl_6_57 word6_57 gnd C_wl
Rw7_57 word7_57 word6_57 R_wl
Cwl_7_57 word7_57 gnd C_wl
Rw8_57 word8_57 word7_57 R_wl
Cwl_8_57 word8_57 gnd C_wl
Rw9_57 word9_57 word8_57 R_wl
Cwl_9_57 word9_57 gnd C_wl
Rw10_57 word10_57 word9_57 R_wl
Cwl_10_57 word10_57 gnd C_wl
Rw11_57 word11_57 word10_57 R_wl
Cwl_11_57 word11_57 gnd C_wl
Rw12_57 word12_57 word11_57 R_wl
Cwl_12_57 word12_57 gnd C_wl
Rw13_57 word13_57 word12_57 R_wl
Cwl_13_57 word13_57 gnd C_wl
Rw14_57 word14_57 word13_57 R_wl
Cwl_14_57 word14_57 gnd C_wl
Rw15_57 word15_57 word14_57 R_wl
Cwl_15_57 word15_57 gnd C_wl
Rw16_57 word16_57 word15_57 R_wl
Cwl_16_57 word16_57 gnd C_wl
Rw17_57 word17_57 word16_57 R_wl
Cwl_17_57 word17_57 gnd C_wl
Rw18_57 word18_57 word17_57 R_wl
Cwl_18_57 word18_57 gnd C_wl
Rw19_57 word19_57 word18_57 R_wl
Cwl_19_57 word19_57 gnd C_wl
Rw20_57 word20_57 word19_57 R_wl
Cwl_20_57 word20_57 gnd C_wl
Rw21_57 word21_57 word20_57 R_wl
Cwl_21_57 word21_57 gnd C_wl
Rw22_57 word22_57 word21_57 R_wl
Cwl_22_57 word22_57 gnd C_wl
Rw23_57 word23_57 word22_57 R_wl
Cwl_23_57 word23_57 gnd C_wl
Rw24_57 word24_57 word23_57 R_wl
Cwl_24_57 word24_57 gnd C_wl
Rw25_57 word25_57 word24_57 R_wl
Cwl_25_57 word25_57 gnd C_wl
Rw26_57 word26_57 word25_57 R_wl
Cwl_26_57 word26_57 gnd C_wl
Rw27_57 word27_57 word26_57 R_wl
Cwl_27_57 word27_57 gnd C_wl
Rw28_57 word28_57 word27_57 R_wl
Cwl_28_57 word28_57 gnd C_wl
Rw29_57 word29_57 word28_57 R_wl
Cwl_29_57 word29_57 gnd C_wl
Rw30_57 word30_57 word29_57 R_wl
Cwl_30_57 word30_57 gnd C_wl
Rw31_57 word31_57 word30_57 R_wl
Cwl_31_57 word31_57 gnd C_wl
Rw32_57 word32_57 word31_57 R_wl
Cwl_32_57 word32_57 gnd C_wl
Rw33_57 word33_57 word32_57 R_wl
Cwl_33_57 word33_57 gnd C_wl
Rw34_57 word34_57 word33_57 R_wl
Cwl_34_57 word34_57 gnd C_wl
Rw35_57 word35_57 word34_57 R_wl
Cwl_35_57 word35_57 gnd C_wl
Rw36_57 word36_57 word35_57 R_wl
Cwl_36_57 word36_57 gnd C_wl
Rw37_57 word37_57 word36_57 R_wl
Cwl_37_57 word37_57 gnd C_wl
Rw38_57 word38_57 word37_57 R_wl
Cwl_38_57 word38_57 gnd C_wl
Rw39_57 word39_57 word38_57 R_wl
Cwl_39_57 word39_57 gnd C_wl
Rw40_57 word40_57 word39_57 R_wl
Cwl_40_57 word40_57 gnd C_wl
Rw41_57 word41_57 word40_57 R_wl
Cwl_41_57 word41_57 gnd C_wl
Rw42_57 word42_57 word41_57 R_wl
Cwl_42_57 word42_57 gnd C_wl
Rw43_57 word43_57 word42_57 R_wl
Cwl_43_57 word43_57 gnd C_wl
Rw44_57 word44_57 word43_57 R_wl
Cwl_44_57 word44_57 gnd C_wl
Rw45_57 word45_57 word44_57 R_wl
Cwl_45_57 word45_57 gnd C_wl
Rw46_57 word46_57 word45_57 R_wl
Cwl_46_57 word46_57 gnd C_wl
Rw47_57 word47_57 word46_57 R_wl
Cwl_47_57 word47_57 gnd C_wl
Rw48_57 word48_57 word47_57 R_wl
Cwl_48_57 word48_57 gnd C_wl
Rw49_57 word49_57 word48_57 R_wl
Cwl_49_57 word49_57 gnd C_wl
Rw50_57 word50_57 word49_57 R_wl
Cwl_50_57 word50_57 gnd C_wl
Rw51_57 word51_57 word50_57 R_wl
Cwl_51_57 word51_57 gnd C_wl
Rw52_57 word52_57 word51_57 R_wl
Cwl_52_57 word52_57 gnd C_wl
Rw53_57 word53_57 word52_57 R_wl
Cwl_53_57 word53_57 gnd C_wl
Rw54_57 word54_57 word53_57 R_wl
Cwl_54_57 word54_57 gnd C_wl
Rw55_57 word55_57 word54_57 R_wl
Cwl_55_57 word55_57 gnd C_wl
Rw56_57 word56_57 word55_57 R_wl
Cwl_56_57 word56_57 gnd C_wl
Rw57_57 word57_57 word56_57 R_wl
Cwl_57_57 word57_57 gnd C_wl
Rw58_57 word58_57 word57_57 R_wl
Cwl_58_57 word58_57 gnd C_wl
Rw59_57 word59_57 word58_57 R_wl
Cwl_59_57 word59_57 gnd C_wl
Rw60_57 word60_57 word59_57 R_wl
Cwl_60_57 word60_57 gnd C_wl
Rw61_57 word61_57 word60_57 R_wl
Cwl_61_57 word61_57 gnd C_wl
Rw62_57 word62_57 word61_57 R_wl
Cwl_62_57 word62_57 gnd C_wl
Rw63_57 word63_57 word62_57 R_wl
Cwl_63_57 word63_57 gnd C_wl
Rw64_57 word64_57 word63_57 R_wl
Cwl_64_57 word64_57 gnd C_wl
Rw65_57 word65_57 word64_57 R_wl
Cwl_65_57 word65_57 gnd C_wl
Rw66_57 word66_57 word65_57 R_wl
Cwl_66_57 word66_57 gnd C_wl
Rw67_57 word67_57 word66_57 R_wl
Cwl_67_57 word67_57 gnd C_wl
Rw68_57 word68_57 word67_57 R_wl
Cwl_68_57 word68_57 gnd C_wl
Rw69_57 word69_57 word68_57 R_wl
Cwl_69_57 word69_57 gnd C_wl
Rw70_57 word70_57 word69_57 R_wl
Cwl_70_57 word70_57 gnd C_wl
Rw71_57 word71_57 word70_57 R_wl
Cwl_71_57 word71_57 gnd C_wl
Rw72_57 word72_57 word71_57 R_wl
Cwl_72_57 word72_57 gnd C_wl
Rw73_57 word73_57 word72_57 R_wl
Cwl_73_57 word73_57 gnd C_wl
Rw74_57 word74_57 word73_57 R_wl
Cwl_74_57 word74_57 gnd C_wl
Rw75_57 word75_57 word74_57 R_wl
Cwl_75_57 word75_57 gnd C_wl
Rw76_57 word76_57 word75_57 R_wl
Cwl_76_57 word76_57 gnd C_wl
Rw77_57 word77_57 word76_57 R_wl
Cwl_77_57 word77_57 gnd C_wl
Rw78_57 word78_57 word77_57 R_wl
Cwl_78_57 word78_57 gnd C_wl
Rw79_57 word79_57 word78_57 R_wl
Cwl_79_57 word79_57 gnd C_wl
Rw80_57 word80_57 word79_57 R_wl
Cwl_80_57 word80_57 gnd C_wl
Rw81_57 word81_57 word80_57 R_wl
Cwl_81_57 word81_57 gnd C_wl
Rw82_57 word82_57 word81_57 R_wl
Cwl_82_57 word82_57 gnd C_wl
Rw83_57 word83_57 word82_57 R_wl
Cwl_83_57 word83_57 gnd C_wl
Rw84_57 word84_57 word83_57 R_wl
Cwl_84_57 word84_57 gnd C_wl
Rw85_57 word85_57 word84_57 R_wl
Cwl_85_57 word85_57 gnd C_wl
Rw86_57 word86_57 word85_57 R_wl
Cwl_86_57 word86_57 gnd C_wl
Rw87_57 word87_57 word86_57 R_wl
Cwl_87_57 word87_57 gnd C_wl
Rw88_57 word88_57 word87_57 R_wl
Cwl_88_57 word88_57 gnd C_wl
Rw89_57 word89_57 word88_57 R_wl
Cwl_89_57 word89_57 gnd C_wl
Rw90_57 word90_57 word89_57 R_wl
Cwl_90_57 word90_57 gnd C_wl
Rw91_57 word91_57 word90_57 R_wl
Cwl_91_57 word91_57 gnd C_wl
Rw92_57 word92_57 word91_57 R_wl
Cwl_92_57 word92_57 gnd C_wl
Rw93_57 word93_57 word92_57 R_wl
Cwl_93_57 word93_57 gnd C_wl
Rw94_57 word94_57 word93_57 R_wl
Cwl_94_57 word94_57 gnd C_wl
Rw95_57 word95_57 word94_57 R_wl
Cwl_95_57 word95_57 gnd C_wl
Rw96_57 word96_57 word95_57 R_wl
Cwl_96_57 word96_57 gnd C_wl
Rw97_57 word97_57 word96_57 R_wl
Cwl_97_57 word97_57 gnd C_wl
Rw98_57 word98_57 word97_57 R_wl
Cwl_98_57 word98_57 gnd C_wl
Rw99_57 word99_57 word98_57 R_wl
Cwl_99_57 word99_57 gnd C_wl
Vwl_58 word_58 0 0
Rw0_58 word_58 word0_58 R_wl
Cwl_0_58 word0_58 gnd C_wl
Rw1_58 word1_58 word0_58 R_wl
Cwl_1_58 word1_58 gnd C_wl
Rw2_58 word2_58 word1_58 R_wl
Cwl_2_58 word2_58 gnd C_wl
Rw3_58 word3_58 word2_58 R_wl
Cwl_3_58 word3_58 gnd C_wl
Rw4_58 word4_58 word3_58 R_wl
Cwl_4_58 word4_58 gnd C_wl
Rw5_58 word5_58 word4_58 R_wl
Cwl_5_58 word5_58 gnd C_wl
Rw6_58 word6_58 word5_58 R_wl
Cwl_6_58 word6_58 gnd C_wl
Rw7_58 word7_58 word6_58 R_wl
Cwl_7_58 word7_58 gnd C_wl
Rw8_58 word8_58 word7_58 R_wl
Cwl_8_58 word8_58 gnd C_wl
Rw9_58 word9_58 word8_58 R_wl
Cwl_9_58 word9_58 gnd C_wl
Rw10_58 word10_58 word9_58 R_wl
Cwl_10_58 word10_58 gnd C_wl
Rw11_58 word11_58 word10_58 R_wl
Cwl_11_58 word11_58 gnd C_wl
Rw12_58 word12_58 word11_58 R_wl
Cwl_12_58 word12_58 gnd C_wl
Rw13_58 word13_58 word12_58 R_wl
Cwl_13_58 word13_58 gnd C_wl
Rw14_58 word14_58 word13_58 R_wl
Cwl_14_58 word14_58 gnd C_wl
Rw15_58 word15_58 word14_58 R_wl
Cwl_15_58 word15_58 gnd C_wl
Rw16_58 word16_58 word15_58 R_wl
Cwl_16_58 word16_58 gnd C_wl
Rw17_58 word17_58 word16_58 R_wl
Cwl_17_58 word17_58 gnd C_wl
Rw18_58 word18_58 word17_58 R_wl
Cwl_18_58 word18_58 gnd C_wl
Rw19_58 word19_58 word18_58 R_wl
Cwl_19_58 word19_58 gnd C_wl
Rw20_58 word20_58 word19_58 R_wl
Cwl_20_58 word20_58 gnd C_wl
Rw21_58 word21_58 word20_58 R_wl
Cwl_21_58 word21_58 gnd C_wl
Rw22_58 word22_58 word21_58 R_wl
Cwl_22_58 word22_58 gnd C_wl
Rw23_58 word23_58 word22_58 R_wl
Cwl_23_58 word23_58 gnd C_wl
Rw24_58 word24_58 word23_58 R_wl
Cwl_24_58 word24_58 gnd C_wl
Rw25_58 word25_58 word24_58 R_wl
Cwl_25_58 word25_58 gnd C_wl
Rw26_58 word26_58 word25_58 R_wl
Cwl_26_58 word26_58 gnd C_wl
Rw27_58 word27_58 word26_58 R_wl
Cwl_27_58 word27_58 gnd C_wl
Rw28_58 word28_58 word27_58 R_wl
Cwl_28_58 word28_58 gnd C_wl
Rw29_58 word29_58 word28_58 R_wl
Cwl_29_58 word29_58 gnd C_wl
Rw30_58 word30_58 word29_58 R_wl
Cwl_30_58 word30_58 gnd C_wl
Rw31_58 word31_58 word30_58 R_wl
Cwl_31_58 word31_58 gnd C_wl
Rw32_58 word32_58 word31_58 R_wl
Cwl_32_58 word32_58 gnd C_wl
Rw33_58 word33_58 word32_58 R_wl
Cwl_33_58 word33_58 gnd C_wl
Rw34_58 word34_58 word33_58 R_wl
Cwl_34_58 word34_58 gnd C_wl
Rw35_58 word35_58 word34_58 R_wl
Cwl_35_58 word35_58 gnd C_wl
Rw36_58 word36_58 word35_58 R_wl
Cwl_36_58 word36_58 gnd C_wl
Rw37_58 word37_58 word36_58 R_wl
Cwl_37_58 word37_58 gnd C_wl
Rw38_58 word38_58 word37_58 R_wl
Cwl_38_58 word38_58 gnd C_wl
Rw39_58 word39_58 word38_58 R_wl
Cwl_39_58 word39_58 gnd C_wl
Rw40_58 word40_58 word39_58 R_wl
Cwl_40_58 word40_58 gnd C_wl
Rw41_58 word41_58 word40_58 R_wl
Cwl_41_58 word41_58 gnd C_wl
Rw42_58 word42_58 word41_58 R_wl
Cwl_42_58 word42_58 gnd C_wl
Rw43_58 word43_58 word42_58 R_wl
Cwl_43_58 word43_58 gnd C_wl
Rw44_58 word44_58 word43_58 R_wl
Cwl_44_58 word44_58 gnd C_wl
Rw45_58 word45_58 word44_58 R_wl
Cwl_45_58 word45_58 gnd C_wl
Rw46_58 word46_58 word45_58 R_wl
Cwl_46_58 word46_58 gnd C_wl
Rw47_58 word47_58 word46_58 R_wl
Cwl_47_58 word47_58 gnd C_wl
Rw48_58 word48_58 word47_58 R_wl
Cwl_48_58 word48_58 gnd C_wl
Rw49_58 word49_58 word48_58 R_wl
Cwl_49_58 word49_58 gnd C_wl
Rw50_58 word50_58 word49_58 R_wl
Cwl_50_58 word50_58 gnd C_wl
Rw51_58 word51_58 word50_58 R_wl
Cwl_51_58 word51_58 gnd C_wl
Rw52_58 word52_58 word51_58 R_wl
Cwl_52_58 word52_58 gnd C_wl
Rw53_58 word53_58 word52_58 R_wl
Cwl_53_58 word53_58 gnd C_wl
Rw54_58 word54_58 word53_58 R_wl
Cwl_54_58 word54_58 gnd C_wl
Rw55_58 word55_58 word54_58 R_wl
Cwl_55_58 word55_58 gnd C_wl
Rw56_58 word56_58 word55_58 R_wl
Cwl_56_58 word56_58 gnd C_wl
Rw57_58 word57_58 word56_58 R_wl
Cwl_57_58 word57_58 gnd C_wl
Rw58_58 word58_58 word57_58 R_wl
Cwl_58_58 word58_58 gnd C_wl
Rw59_58 word59_58 word58_58 R_wl
Cwl_59_58 word59_58 gnd C_wl
Rw60_58 word60_58 word59_58 R_wl
Cwl_60_58 word60_58 gnd C_wl
Rw61_58 word61_58 word60_58 R_wl
Cwl_61_58 word61_58 gnd C_wl
Rw62_58 word62_58 word61_58 R_wl
Cwl_62_58 word62_58 gnd C_wl
Rw63_58 word63_58 word62_58 R_wl
Cwl_63_58 word63_58 gnd C_wl
Rw64_58 word64_58 word63_58 R_wl
Cwl_64_58 word64_58 gnd C_wl
Rw65_58 word65_58 word64_58 R_wl
Cwl_65_58 word65_58 gnd C_wl
Rw66_58 word66_58 word65_58 R_wl
Cwl_66_58 word66_58 gnd C_wl
Rw67_58 word67_58 word66_58 R_wl
Cwl_67_58 word67_58 gnd C_wl
Rw68_58 word68_58 word67_58 R_wl
Cwl_68_58 word68_58 gnd C_wl
Rw69_58 word69_58 word68_58 R_wl
Cwl_69_58 word69_58 gnd C_wl
Rw70_58 word70_58 word69_58 R_wl
Cwl_70_58 word70_58 gnd C_wl
Rw71_58 word71_58 word70_58 R_wl
Cwl_71_58 word71_58 gnd C_wl
Rw72_58 word72_58 word71_58 R_wl
Cwl_72_58 word72_58 gnd C_wl
Rw73_58 word73_58 word72_58 R_wl
Cwl_73_58 word73_58 gnd C_wl
Rw74_58 word74_58 word73_58 R_wl
Cwl_74_58 word74_58 gnd C_wl
Rw75_58 word75_58 word74_58 R_wl
Cwl_75_58 word75_58 gnd C_wl
Rw76_58 word76_58 word75_58 R_wl
Cwl_76_58 word76_58 gnd C_wl
Rw77_58 word77_58 word76_58 R_wl
Cwl_77_58 word77_58 gnd C_wl
Rw78_58 word78_58 word77_58 R_wl
Cwl_78_58 word78_58 gnd C_wl
Rw79_58 word79_58 word78_58 R_wl
Cwl_79_58 word79_58 gnd C_wl
Rw80_58 word80_58 word79_58 R_wl
Cwl_80_58 word80_58 gnd C_wl
Rw81_58 word81_58 word80_58 R_wl
Cwl_81_58 word81_58 gnd C_wl
Rw82_58 word82_58 word81_58 R_wl
Cwl_82_58 word82_58 gnd C_wl
Rw83_58 word83_58 word82_58 R_wl
Cwl_83_58 word83_58 gnd C_wl
Rw84_58 word84_58 word83_58 R_wl
Cwl_84_58 word84_58 gnd C_wl
Rw85_58 word85_58 word84_58 R_wl
Cwl_85_58 word85_58 gnd C_wl
Rw86_58 word86_58 word85_58 R_wl
Cwl_86_58 word86_58 gnd C_wl
Rw87_58 word87_58 word86_58 R_wl
Cwl_87_58 word87_58 gnd C_wl
Rw88_58 word88_58 word87_58 R_wl
Cwl_88_58 word88_58 gnd C_wl
Rw89_58 word89_58 word88_58 R_wl
Cwl_89_58 word89_58 gnd C_wl
Rw90_58 word90_58 word89_58 R_wl
Cwl_90_58 word90_58 gnd C_wl
Rw91_58 word91_58 word90_58 R_wl
Cwl_91_58 word91_58 gnd C_wl
Rw92_58 word92_58 word91_58 R_wl
Cwl_92_58 word92_58 gnd C_wl
Rw93_58 word93_58 word92_58 R_wl
Cwl_93_58 word93_58 gnd C_wl
Rw94_58 word94_58 word93_58 R_wl
Cwl_94_58 word94_58 gnd C_wl
Rw95_58 word95_58 word94_58 R_wl
Cwl_95_58 word95_58 gnd C_wl
Rw96_58 word96_58 word95_58 R_wl
Cwl_96_58 word96_58 gnd C_wl
Rw97_58 word97_58 word96_58 R_wl
Cwl_97_58 word97_58 gnd C_wl
Rw98_58 word98_58 word97_58 R_wl
Cwl_98_58 word98_58 gnd C_wl
Rw99_58 word99_58 word98_58 R_wl
Cwl_99_58 word99_58 gnd C_wl
Vwl_59 word_59 0 0
Rw0_59 word_59 word0_59 R_wl
Cwl_0_59 word0_59 gnd C_wl
Rw1_59 word1_59 word0_59 R_wl
Cwl_1_59 word1_59 gnd C_wl
Rw2_59 word2_59 word1_59 R_wl
Cwl_2_59 word2_59 gnd C_wl
Rw3_59 word3_59 word2_59 R_wl
Cwl_3_59 word3_59 gnd C_wl
Rw4_59 word4_59 word3_59 R_wl
Cwl_4_59 word4_59 gnd C_wl
Rw5_59 word5_59 word4_59 R_wl
Cwl_5_59 word5_59 gnd C_wl
Rw6_59 word6_59 word5_59 R_wl
Cwl_6_59 word6_59 gnd C_wl
Rw7_59 word7_59 word6_59 R_wl
Cwl_7_59 word7_59 gnd C_wl
Rw8_59 word8_59 word7_59 R_wl
Cwl_8_59 word8_59 gnd C_wl
Rw9_59 word9_59 word8_59 R_wl
Cwl_9_59 word9_59 gnd C_wl
Rw10_59 word10_59 word9_59 R_wl
Cwl_10_59 word10_59 gnd C_wl
Rw11_59 word11_59 word10_59 R_wl
Cwl_11_59 word11_59 gnd C_wl
Rw12_59 word12_59 word11_59 R_wl
Cwl_12_59 word12_59 gnd C_wl
Rw13_59 word13_59 word12_59 R_wl
Cwl_13_59 word13_59 gnd C_wl
Rw14_59 word14_59 word13_59 R_wl
Cwl_14_59 word14_59 gnd C_wl
Rw15_59 word15_59 word14_59 R_wl
Cwl_15_59 word15_59 gnd C_wl
Rw16_59 word16_59 word15_59 R_wl
Cwl_16_59 word16_59 gnd C_wl
Rw17_59 word17_59 word16_59 R_wl
Cwl_17_59 word17_59 gnd C_wl
Rw18_59 word18_59 word17_59 R_wl
Cwl_18_59 word18_59 gnd C_wl
Rw19_59 word19_59 word18_59 R_wl
Cwl_19_59 word19_59 gnd C_wl
Rw20_59 word20_59 word19_59 R_wl
Cwl_20_59 word20_59 gnd C_wl
Rw21_59 word21_59 word20_59 R_wl
Cwl_21_59 word21_59 gnd C_wl
Rw22_59 word22_59 word21_59 R_wl
Cwl_22_59 word22_59 gnd C_wl
Rw23_59 word23_59 word22_59 R_wl
Cwl_23_59 word23_59 gnd C_wl
Rw24_59 word24_59 word23_59 R_wl
Cwl_24_59 word24_59 gnd C_wl
Rw25_59 word25_59 word24_59 R_wl
Cwl_25_59 word25_59 gnd C_wl
Rw26_59 word26_59 word25_59 R_wl
Cwl_26_59 word26_59 gnd C_wl
Rw27_59 word27_59 word26_59 R_wl
Cwl_27_59 word27_59 gnd C_wl
Rw28_59 word28_59 word27_59 R_wl
Cwl_28_59 word28_59 gnd C_wl
Rw29_59 word29_59 word28_59 R_wl
Cwl_29_59 word29_59 gnd C_wl
Rw30_59 word30_59 word29_59 R_wl
Cwl_30_59 word30_59 gnd C_wl
Rw31_59 word31_59 word30_59 R_wl
Cwl_31_59 word31_59 gnd C_wl
Rw32_59 word32_59 word31_59 R_wl
Cwl_32_59 word32_59 gnd C_wl
Rw33_59 word33_59 word32_59 R_wl
Cwl_33_59 word33_59 gnd C_wl
Rw34_59 word34_59 word33_59 R_wl
Cwl_34_59 word34_59 gnd C_wl
Rw35_59 word35_59 word34_59 R_wl
Cwl_35_59 word35_59 gnd C_wl
Rw36_59 word36_59 word35_59 R_wl
Cwl_36_59 word36_59 gnd C_wl
Rw37_59 word37_59 word36_59 R_wl
Cwl_37_59 word37_59 gnd C_wl
Rw38_59 word38_59 word37_59 R_wl
Cwl_38_59 word38_59 gnd C_wl
Rw39_59 word39_59 word38_59 R_wl
Cwl_39_59 word39_59 gnd C_wl
Rw40_59 word40_59 word39_59 R_wl
Cwl_40_59 word40_59 gnd C_wl
Rw41_59 word41_59 word40_59 R_wl
Cwl_41_59 word41_59 gnd C_wl
Rw42_59 word42_59 word41_59 R_wl
Cwl_42_59 word42_59 gnd C_wl
Rw43_59 word43_59 word42_59 R_wl
Cwl_43_59 word43_59 gnd C_wl
Rw44_59 word44_59 word43_59 R_wl
Cwl_44_59 word44_59 gnd C_wl
Rw45_59 word45_59 word44_59 R_wl
Cwl_45_59 word45_59 gnd C_wl
Rw46_59 word46_59 word45_59 R_wl
Cwl_46_59 word46_59 gnd C_wl
Rw47_59 word47_59 word46_59 R_wl
Cwl_47_59 word47_59 gnd C_wl
Rw48_59 word48_59 word47_59 R_wl
Cwl_48_59 word48_59 gnd C_wl
Rw49_59 word49_59 word48_59 R_wl
Cwl_49_59 word49_59 gnd C_wl
Rw50_59 word50_59 word49_59 R_wl
Cwl_50_59 word50_59 gnd C_wl
Rw51_59 word51_59 word50_59 R_wl
Cwl_51_59 word51_59 gnd C_wl
Rw52_59 word52_59 word51_59 R_wl
Cwl_52_59 word52_59 gnd C_wl
Rw53_59 word53_59 word52_59 R_wl
Cwl_53_59 word53_59 gnd C_wl
Rw54_59 word54_59 word53_59 R_wl
Cwl_54_59 word54_59 gnd C_wl
Rw55_59 word55_59 word54_59 R_wl
Cwl_55_59 word55_59 gnd C_wl
Rw56_59 word56_59 word55_59 R_wl
Cwl_56_59 word56_59 gnd C_wl
Rw57_59 word57_59 word56_59 R_wl
Cwl_57_59 word57_59 gnd C_wl
Rw58_59 word58_59 word57_59 R_wl
Cwl_58_59 word58_59 gnd C_wl
Rw59_59 word59_59 word58_59 R_wl
Cwl_59_59 word59_59 gnd C_wl
Rw60_59 word60_59 word59_59 R_wl
Cwl_60_59 word60_59 gnd C_wl
Rw61_59 word61_59 word60_59 R_wl
Cwl_61_59 word61_59 gnd C_wl
Rw62_59 word62_59 word61_59 R_wl
Cwl_62_59 word62_59 gnd C_wl
Rw63_59 word63_59 word62_59 R_wl
Cwl_63_59 word63_59 gnd C_wl
Rw64_59 word64_59 word63_59 R_wl
Cwl_64_59 word64_59 gnd C_wl
Rw65_59 word65_59 word64_59 R_wl
Cwl_65_59 word65_59 gnd C_wl
Rw66_59 word66_59 word65_59 R_wl
Cwl_66_59 word66_59 gnd C_wl
Rw67_59 word67_59 word66_59 R_wl
Cwl_67_59 word67_59 gnd C_wl
Rw68_59 word68_59 word67_59 R_wl
Cwl_68_59 word68_59 gnd C_wl
Rw69_59 word69_59 word68_59 R_wl
Cwl_69_59 word69_59 gnd C_wl
Rw70_59 word70_59 word69_59 R_wl
Cwl_70_59 word70_59 gnd C_wl
Rw71_59 word71_59 word70_59 R_wl
Cwl_71_59 word71_59 gnd C_wl
Rw72_59 word72_59 word71_59 R_wl
Cwl_72_59 word72_59 gnd C_wl
Rw73_59 word73_59 word72_59 R_wl
Cwl_73_59 word73_59 gnd C_wl
Rw74_59 word74_59 word73_59 R_wl
Cwl_74_59 word74_59 gnd C_wl
Rw75_59 word75_59 word74_59 R_wl
Cwl_75_59 word75_59 gnd C_wl
Rw76_59 word76_59 word75_59 R_wl
Cwl_76_59 word76_59 gnd C_wl
Rw77_59 word77_59 word76_59 R_wl
Cwl_77_59 word77_59 gnd C_wl
Rw78_59 word78_59 word77_59 R_wl
Cwl_78_59 word78_59 gnd C_wl
Rw79_59 word79_59 word78_59 R_wl
Cwl_79_59 word79_59 gnd C_wl
Rw80_59 word80_59 word79_59 R_wl
Cwl_80_59 word80_59 gnd C_wl
Rw81_59 word81_59 word80_59 R_wl
Cwl_81_59 word81_59 gnd C_wl
Rw82_59 word82_59 word81_59 R_wl
Cwl_82_59 word82_59 gnd C_wl
Rw83_59 word83_59 word82_59 R_wl
Cwl_83_59 word83_59 gnd C_wl
Rw84_59 word84_59 word83_59 R_wl
Cwl_84_59 word84_59 gnd C_wl
Rw85_59 word85_59 word84_59 R_wl
Cwl_85_59 word85_59 gnd C_wl
Rw86_59 word86_59 word85_59 R_wl
Cwl_86_59 word86_59 gnd C_wl
Rw87_59 word87_59 word86_59 R_wl
Cwl_87_59 word87_59 gnd C_wl
Rw88_59 word88_59 word87_59 R_wl
Cwl_88_59 word88_59 gnd C_wl
Rw89_59 word89_59 word88_59 R_wl
Cwl_89_59 word89_59 gnd C_wl
Rw90_59 word90_59 word89_59 R_wl
Cwl_90_59 word90_59 gnd C_wl
Rw91_59 word91_59 word90_59 R_wl
Cwl_91_59 word91_59 gnd C_wl
Rw92_59 word92_59 word91_59 R_wl
Cwl_92_59 word92_59 gnd C_wl
Rw93_59 word93_59 word92_59 R_wl
Cwl_93_59 word93_59 gnd C_wl
Rw94_59 word94_59 word93_59 R_wl
Cwl_94_59 word94_59 gnd C_wl
Rw95_59 word95_59 word94_59 R_wl
Cwl_95_59 word95_59 gnd C_wl
Rw96_59 word96_59 word95_59 R_wl
Cwl_96_59 word96_59 gnd C_wl
Rw97_59 word97_59 word96_59 R_wl
Cwl_97_59 word97_59 gnd C_wl
Rw98_59 word98_59 word97_59 R_wl
Cwl_98_59 word98_59 gnd C_wl
Rw99_59 word99_59 word98_59 R_wl
Cwl_99_59 word99_59 gnd C_wl
Vwl_60 word_60 0 0
Rw0_60 word_60 word0_60 R_wl
Cwl_0_60 word0_60 gnd C_wl
Rw1_60 word1_60 word0_60 R_wl
Cwl_1_60 word1_60 gnd C_wl
Rw2_60 word2_60 word1_60 R_wl
Cwl_2_60 word2_60 gnd C_wl
Rw3_60 word3_60 word2_60 R_wl
Cwl_3_60 word3_60 gnd C_wl
Rw4_60 word4_60 word3_60 R_wl
Cwl_4_60 word4_60 gnd C_wl
Rw5_60 word5_60 word4_60 R_wl
Cwl_5_60 word5_60 gnd C_wl
Rw6_60 word6_60 word5_60 R_wl
Cwl_6_60 word6_60 gnd C_wl
Rw7_60 word7_60 word6_60 R_wl
Cwl_7_60 word7_60 gnd C_wl
Rw8_60 word8_60 word7_60 R_wl
Cwl_8_60 word8_60 gnd C_wl
Rw9_60 word9_60 word8_60 R_wl
Cwl_9_60 word9_60 gnd C_wl
Rw10_60 word10_60 word9_60 R_wl
Cwl_10_60 word10_60 gnd C_wl
Rw11_60 word11_60 word10_60 R_wl
Cwl_11_60 word11_60 gnd C_wl
Rw12_60 word12_60 word11_60 R_wl
Cwl_12_60 word12_60 gnd C_wl
Rw13_60 word13_60 word12_60 R_wl
Cwl_13_60 word13_60 gnd C_wl
Rw14_60 word14_60 word13_60 R_wl
Cwl_14_60 word14_60 gnd C_wl
Rw15_60 word15_60 word14_60 R_wl
Cwl_15_60 word15_60 gnd C_wl
Rw16_60 word16_60 word15_60 R_wl
Cwl_16_60 word16_60 gnd C_wl
Rw17_60 word17_60 word16_60 R_wl
Cwl_17_60 word17_60 gnd C_wl
Rw18_60 word18_60 word17_60 R_wl
Cwl_18_60 word18_60 gnd C_wl
Rw19_60 word19_60 word18_60 R_wl
Cwl_19_60 word19_60 gnd C_wl
Rw20_60 word20_60 word19_60 R_wl
Cwl_20_60 word20_60 gnd C_wl
Rw21_60 word21_60 word20_60 R_wl
Cwl_21_60 word21_60 gnd C_wl
Rw22_60 word22_60 word21_60 R_wl
Cwl_22_60 word22_60 gnd C_wl
Rw23_60 word23_60 word22_60 R_wl
Cwl_23_60 word23_60 gnd C_wl
Rw24_60 word24_60 word23_60 R_wl
Cwl_24_60 word24_60 gnd C_wl
Rw25_60 word25_60 word24_60 R_wl
Cwl_25_60 word25_60 gnd C_wl
Rw26_60 word26_60 word25_60 R_wl
Cwl_26_60 word26_60 gnd C_wl
Rw27_60 word27_60 word26_60 R_wl
Cwl_27_60 word27_60 gnd C_wl
Rw28_60 word28_60 word27_60 R_wl
Cwl_28_60 word28_60 gnd C_wl
Rw29_60 word29_60 word28_60 R_wl
Cwl_29_60 word29_60 gnd C_wl
Rw30_60 word30_60 word29_60 R_wl
Cwl_30_60 word30_60 gnd C_wl
Rw31_60 word31_60 word30_60 R_wl
Cwl_31_60 word31_60 gnd C_wl
Rw32_60 word32_60 word31_60 R_wl
Cwl_32_60 word32_60 gnd C_wl
Rw33_60 word33_60 word32_60 R_wl
Cwl_33_60 word33_60 gnd C_wl
Rw34_60 word34_60 word33_60 R_wl
Cwl_34_60 word34_60 gnd C_wl
Rw35_60 word35_60 word34_60 R_wl
Cwl_35_60 word35_60 gnd C_wl
Rw36_60 word36_60 word35_60 R_wl
Cwl_36_60 word36_60 gnd C_wl
Rw37_60 word37_60 word36_60 R_wl
Cwl_37_60 word37_60 gnd C_wl
Rw38_60 word38_60 word37_60 R_wl
Cwl_38_60 word38_60 gnd C_wl
Rw39_60 word39_60 word38_60 R_wl
Cwl_39_60 word39_60 gnd C_wl
Rw40_60 word40_60 word39_60 R_wl
Cwl_40_60 word40_60 gnd C_wl
Rw41_60 word41_60 word40_60 R_wl
Cwl_41_60 word41_60 gnd C_wl
Rw42_60 word42_60 word41_60 R_wl
Cwl_42_60 word42_60 gnd C_wl
Rw43_60 word43_60 word42_60 R_wl
Cwl_43_60 word43_60 gnd C_wl
Rw44_60 word44_60 word43_60 R_wl
Cwl_44_60 word44_60 gnd C_wl
Rw45_60 word45_60 word44_60 R_wl
Cwl_45_60 word45_60 gnd C_wl
Rw46_60 word46_60 word45_60 R_wl
Cwl_46_60 word46_60 gnd C_wl
Rw47_60 word47_60 word46_60 R_wl
Cwl_47_60 word47_60 gnd C_wl
Rw48_60 word48_60 word47_60 R_wl
Cwl_48_60 word48_60 gnd C_wl
Rw49_60 word49_60 word48_60 R_wl
Cwl_49_60 word49_60 gnd C_wl
Rw50_60 word50_60 word49_60 R_wl
Cwl_50_60 word50_60 gnd C_wl
Rw51_60 word51_60 word50_60 R_wl
Cwl_51_60 word51_60 gnd C_wl
Rw52_60 word52_60 word51_60 R_wl
Cwl_52_60 word52_60 gnd C_wl
Rw53_60 word53_60 word52_60 R_wl
Cwl_53_60 word53_60 gnd C_wl
Rw54_60 word54_60 word53_60 R_wl
Cwl_54_60 word54_60 gnd C_wl
Rw55_60 word55_60 word54_60 R_wl
Cwl_55_60 word55_60 gnd C_wl
Rw56_60 word56_60 word55_60 R_wl
Cwl_56_60 word56_60 gnd C_wl
Rw57_60 word57_60 word56_60 R_wl
Cwl_57_60 word57_60 gnd C_wl
Rw58_60 word58_60 word57_60 R_wl
Cwl_58_60 word58_60 gnd C_wl
Rw59_60 word59_60 word58_60 R_wl
Cwl_59_60 word59_60 gnd C_wl
Rw60_60 word60_60 word59_60 R_wl
Cwl_60_60 word60_60 gnd C_wl
Rw61_60 word61_60 word60_60 R_wl
Cwl_61_60 word61_60 gnd C_wl
Rw62_60 word62_60 word61_60 R_wl
Cwl_62_60 word62_60 gnd C_wl
Rw63_60 word63_60 word62_60 R_wl
Cwl_63_60 word63_60 gnd C_wl
Rw64_60 word64_60 word63_60 R_wl
Cwl_64_60 word64_60 gnd C_wl
Rw65_60 word65_60 word64_60 R_wl
Cwl_65_60 word65_60 gnd C_wl
Rw66_60 word66_60 word65_60 R_wl
Cwl_66_60 word66_60 gnd C_wl
Rw67_60 word67_60 word66_60 R_wl
Cwl_67_60 word67_60 gnd C_wl
Rw68_60 word68_60 word67_60 R_wl
Cwl_68_60 word68_60 gnd C_wl
Rw69_60 word69_60 word68_60 R_wl
Cwl_69_60 word69_60 gnd C_wl
Rw70_60 word70_60 word69_60 R_wl
Cwl_70_60 word70_60 gnd C_wl
Rw71_60 word71_60 word70_60 R_wl
Cwl_71_60 word71_60 gnd C_wl
Rw72_60 word72_60 word71_60 R_wl
Cwl_72_60 word72_60 gnd C_wl
Rw73_60 word73_60 word72_60 R_wl
Cwl_73_60 word73_60 gnd C_wl
Rw74_60 word74_60 word73_60 R_wl
Cwl_74_60 word74_60 gnd C_wl
Rw75_60 word75_60 word74_60 R_wl
Cwl_75_60 word75_60 gnd C_wl
Rw76_60 word76_60 word75_60 R_wl
Cwl_76_60 word76_60 gnd C_wl
Rw77_60 word77_60 word76_60 R_wl
Cwl_77_60 word77_60 gnd C_wl
Rw78_60 word78_60 word77_60 R_wl
Cwl_78_60 word78_60 gnd C_wl
Rw79_60 word79_60 word78_60 R_wl
Cwl_79_60 word79_60 gnd C_wl
Rw80_60 word80_60 word79_60 R_wl
Cwl_80_60 word80_60 gnd C_wl
Rw81_60 word81_60 word80_60 R_wl
Cwl_81_60 word81_60 gnd C_wl
Rw82_60 word82_60 word81_60 R_wl
Cwl_82_60 word82_60 gnd C_wl
Rw83_60 word83_60 word82_60 R_wl
Cwl_83_60 word83_60 gnd C_wl
Rw84_60 word84_60 word83_60 R_wl
Cwl_84_60 word84_60 gnd C_wl
Rw85_60 word85_60 word84_60 R_wl
Cwl_85_60 word85_60 gnd C_wl
Rw86_60 word86_60 word85_60 R_wl
Cwl_86_60 word86_60 gnd C_wl
Rw87_60 word87_60 word86_60 R_wl
Cwl_87_60 word87_60 gnd C_wl
Rw88_60 word88_60 word87_60 R_wl
Cwl_88_60 word88_60 gnd C_wl
Rw89_60 word89_60 word88_60 R_wl
Cwl_89_60 word89_60 gnd C_wl
Rw90_60 word90_60 word89_60 R_wl
Cwl_90_60 word90_60 gnd C_wl
Rw91_60 word91_60 word90_60 R_wl
Cwl_91_60 word91_60 gnd C_wl
Rw92_60 word92_60 word91_60 R_wl
Cwl_92_60 word92_60 gnd C_wl
Rw93_60 word93_60 word92_60 R_wl
Cwl_93_60 word93_60 gnd C_wl
Rw94_60 word94_60 word93_60 R_wl
Cwl_94_60 word94_60 gnd C_wl
Rw95_60 word95_60 word94_60 R_wl
Cwl_95_60 word95_60 gnd C_wl
Rw96_60 word96_60 word95_60 R_wl
Cwl_96_60 word96_60 gnd C_wl
Rw97_60 word97_60 word96_60 R_wl
Cwl_97_60 word97_60 gnd C_wl
Rw98_60 word98_60 word97_60 R_wl
Cwl_98_60 word98_60 gnd C_wl
Rw99_60 word99_60 word98_60 R_wl
Cwl_99_60 word99_60 gnd C_wl
Vwl_61 word_61 0 0
Rw0_61 word_61 word0_61 R_wl
Cwl_0_61 word0_61 gnd C_wl
Rw1_61 word1_61 word0_61 R_wl
Cwl_1_61 word1_61 gnd C_wl
Rw2_61 word2_61 word1_61 R_wl
Cwl_2_61 word2_61 gnd C_wl
Rw3_61 word3_61 word2_61 R_wl
Cwl_3_61 word3_61 gnd C_wl
Rw4_61 word4_61 word3_61 R_wl
Cwl_4_61 word4_61 gnd C_wl
Rw5_61 word5_61 word4_61 R_wl
Cwl_5_61 word5_61 gnd C_wl
Rw6_61 word6_61 word5_61 R_wl
Cwl_6_61 word6_61 gnd C_wl
Rw7_61 word7_61 word6_61 R_wl
Cwl_7_61 word7_61 gnd C_wl
Rw8_61 word8_61 word7_61 R_wl
Cwl_8_61 word8_61 gnd C_wl
Rw9_61 word9_61 word8_61 R_wl
Cwl_9_61 word9_61 gnd C_wl
Rw10_61 word10_61 word9_61 R_wl
Cwl_10_61 word10_61 gnd C_wl
Rw11_61 word11_61 word10_61 R_wl
Cwl_11_61 word11_61 gnd C_wl
Rw12_61 word12_61 word11_61 R_wl
Cwl_12_61 word12_61 gnd C_wl
Rw13_61 word13_61 word12_61 R_wl
Cwl_13_61 word13_61 gnd C_wl
Rw14_61 word14_61 word13_61 R_wl
Cwl_14_61 word14_61 gnd C_wl
Rw15_61 word15_61 word14_61 R_wl
Cwl_15_61 word15_61 gnd C_wl
Rw16_61 word16_61 word15_61 R_wl
Cwl_16_61 word16_61 gnd C_wl
Rw17_61 word17_61 word16_61 R_wl
Cwl_17_61 word17_61 gnd C_wl
Rw18_61 word18_61 word17_61 R_wl
Cwl_18_61 word18_61 gnd C_wl
Rw19_61 word19_61 word18_61 R_wl
Cwl_19_61 word19_61 gnd C_wl
Rw20_61 word20_61 word19_61 R_wl
Cwl_20_61 word20_61 gnd C_wl
Rw21_61 word21_61 word20_61 R_wl
Cwl_21_61 word21_61 gnd C_wl
Rw22_61 word22_61 word21_61 R_wl
Cwl_22_61 word22_61 gnd C_wl
Rw23_61 word23_61 word22_61 R_wl
Cwl_23_61 word23_61 gnd C_wl
Rw24_61 word24_61 word23_61 R_wl
Cwl_24_61 word24_61 gnd C_wl
Rw25_61 word25_61 word24_61 R_wl
Cwl_25_61 word25_61 gnd C_wl
Rw26_61 word26_61 word25_61 R_wl
Cwl_26_61 word26_61 gnd C_wl
Rw27_61 word27_61 word26_61 R_wl
Cwl_27_61 word27_61 gnd C_wl
Rw28_61 word28_61 word27_61 R_wl
Cwl_28_61 word28_61 gnd C_wl
Rw29_61 word29_61 word28_61 R_wl
Cwl_29_61 word29_61 gnd C_wl
Rw30_61 word30_61 word29_61 R_wl
Cwl_30_61 word30_61 gnd C_wl
Rw31_61 word31_61 word30_61 R_wl
Cwl_31_61 word31_61 gnd C_wl
Rw32_61 word32_61 word31_61 R_wl
Cwl_32_61 word32_61 gnd C_wl
Rw33_61 word33_61 word32_61 R_wl
Cwl_33_61 word33_61 gnd C_wl
Rw34_61 word34_61 word33_61 R_wl
Cwl_34_61 word34_61 gnd C_wl
Rw35_61 word35_61 word34_61 R_wl
Cwl_35_61 word35_61 gnd C_wl
Rw36_61 word36_61 word35_61 R_wl
Cwl_36_61 word36_61 gnd C_wl
Rw37_61 word37_61 word36_61 R_wl
Cwl_37_61 word37_61 gnd C_wl
Rw38_61 word38_61 word37_61 R_wl
Cwl_38_61 word38_61 gnd C_wl
Rw39_61 word39_61 word38_61 R_wl
Cwl_39_61 word39_61 gnd C_wl
Rw40_61 word40_61 word39_61 R_wl
Cwl_40_61 word40_61 gnd C_wl
Rw41_61 word41_61 word40_61 R_wl
Cwl_41_61 word41_61 gnd C_wl
Rw42_61 word42_61 word41_61 R_wl
Cwl_42_61 word42_61 gnd C_wl
Rw43_61 word43_61 word42_61 R_wl
Cwl_43_61 word43_61 gnd C_wl
Rw44_61 word44_61 word43_61 R_wl
Cwl_44_61 word44_61 gnd C_wl
Rw45_61 word45_61 word44_61 R_wl
Cwl_45_61 word45_61 gnd C_wl
Rw46_61 word46_61 word45_61 R_wl
Cwl_46_61 word46_61 gnd C_wl
Rw47_61 word47_61 word46_61 R_wl
Cwl_47_61 word47_61 gnd C_wl
Rw48_61 word48_61 word47_61 R_wl
Cwl_48_61 word48_61 gnd C_wl
Rw49_61 word49_61 word48_61 R_wl
Cwl_49_61 word49_61 gnd C_wl
Rw50_61 word50_61 word49_61 R_wl
Cwl_50_61 word50_61 gnd C_wl
Rw51_61 word51_61 word50_61 R_wl
Cwl_51_61 word51_61 gnd C_wl
Rw52_61 word52_61 word51_61 R_wl
Cwl_52_61 word52_61 gnd C_wl
Rw53_61 word53_61 word52_61 R_wl
Cwl_53_61 word53_61 gnd C_wl
Rw54_61 word54_61 word53_61 R_wl
Cwl_54_61 word54_61 gnd C_wl
Rw55_61 word55_61 word54_61 R_wl
Cwl_55_61 word55_61 gnd C_wl
Rw56_61 word56_61 word55_61 R_wl
Cwl_56_61 word56_61 gnd C_wl
Rw57_61 word57_61 word56_61 R_wl
Cwl_57_61 word57_61 gnd C_wl
Rw58_61 word58_61 word57_61 R_wl
Cwl_58_61 word58_61 gnd C_wl
Rw59_61 word59_61 word58_61 R_wl
Cwl_59_61 word59_61 gnd C_wl
Rw60_61 word60_61 word59_61 R_wl
Cwl_60_61 word60_61 gnd C_wl
Rw61_61 word61_61 word60_61 R_wl
Cwl_61_61 word61_61 gnd C_wl
Rw62_61 word62_61 word61_61 R_wl
Cwl_62_61 word62_61 gnd C_wl
Rw63_61 word63_61 word62_61 R_wl
Cwl_63_61 word63_61 gnd C_wl
Rw64_61 word64_61 word63_61 R_wl
Cwl_64_61 word64_61 gnd C_wl
Rw65_61 word65_61 word64_61 R_wl
Cwl_65_61 word65_61 gnd C_wl
Rw66_61 word66_61 word65_61 R_wl
Cwl_66_61 word66_61 gnd C_wl
Rw67_61 word67_61 word66_61 R_wl
Cwl_67_61 word67_61 gnd C_wl
Rw68_61 word68_61 word67_61 R_wl
Cwl_68_61 word68_61 gnd C_wl
Rw69_61 word69_61 word68_61 R_wl
Cwl_69_61 word69_61 gnd C_wl
Rw70_61 word70_61 word69_61 R_wl
Cwl_70_61 word70_61 gnd C_wl
Rw71_61 word71_61 word70_61 R_wl
Cwl_71_61 word71_61 gnd C_wl
Rw72_61 word72_61 word71_61 R_wl
Cwl_72_61 word72_61 gnd C_wl
Rw73_61 word73_61 word72_61 R_wl
Cwl_73_61 word73_61 gnd C_wl
Rw74_61 word74_61 word73_61 R_wl
Cwl_74_61 word74_61 gnd C_wl
Rw75_61 word75_61 word74_61 R_wl
Cwl_75_61 word75_61 gnd C_wl
Rw76_61 word76_61 word75_61 R_wl
Cwl_76_61 word76_61 gnd C_wl
Rw77_61 word77_61 word76_61 R_wl
Cwl_77_61 word77_61 gnd C_wl
Rw78_61 word78_61 word77_61 R_wl
Cwl_78_61 word78_61 gnd C_wl
Rw79_61 word79_61 word78_61 R_wl
Cwl_79_61 word79_61 gnd C_wl
Rw80_61 word80_61 word79_61 R_wl
Cwl_80_61 word80_61 gnd C_wl
Rw81_61 word81_61 word80_61 R_wl
Cwl_81_61 word81_61 gnd C_wl
Rw82_61 word82_61 word81_61 R_wl
Cwl_82_61 word82_61 gnd C_wl
Rw83_61 word83_61 word82_61 R_wl
Cwl_83_61 word83_61 gnd C_wl
Rw84_61 word84_61 word83_61 R_wl
Cwl_84_61 word84_61 gnd C_wl
Rw85_61 word85_61 word84_61 R_wl
Cwl_85_61 word85_61 gnd C_wl
Rw86_61 word86_61 word85_61 R_wl
Cwl_86_61 word86_61 gnd C_wl
Rw87_61 word87_61 word86_61 R_wl
Cwl_87_61 word87_61 gnd C_wl
Rw88_61 word88_61 word87_61 R_wl
Cwl_88_61 word88_61 gnd C_wl
Rw89_61 word89_61 word88_61 R_wl
Cwl_89_61 word89_61 gnd C_wl
Rw90_61 word90_61 word89_61 R_wl
Cwl_90_61 word90_61 gnd C_wl
Rw91_61 word91_61 word90_61 R_wl
Cwl_91_61 word91_61 gnd C_wl
Rw92_61 word92_61 word91_61 R_wl
Cwl_92_61 word92_61 gnd C_wl
Rw93_61 word93_61 word92_61 R_wl
Cwl_93_61 word93_61 gnd C_wl
Rw94_61 word94_61 word93_61 R_wl
Cwl_94_61 word94_61 gnd C_wl
Rw95_61 word95_61 word94_61 R_wl
Cwl_95_61 word95_61 gnd C_wl
Rw96_61 word96_61 word95_61 R_wl
Cwl_96_61 word96_61 gnd C_wl
Rw97_61 word97_61 word96_61 R_wl
Cwl_97_61 word97_61 gnd C_wl
Rw98_61 word98_61 word97_61 R_wl
Cwl_98_61 word98_61 gnd C_wl
Rw99_61 word99_61 word98_61 R_wl
Cwl_99_61 word99_61 gnd C_wl
Vwl_62 word_62 0 0
Rw0_62 word_62 word0_62 R_wl
Cwl_0_62 word0_62 gnd C_wl
Rw1_62 word1_62 word0_62 R_wl
Cwl_1_62 word1_62 gnd C_wl
Rw2_62 word2_62 word1_62 R_wl
Cwl_2_62 word2_62 gnd C_wl
Rw3_62 word3_62 word2_62 R_wl
Cwl_3_62 word3_62 gnd C_wl
Rw4_62 word4_62 word3_62 R_wl
Cwl_4_62 word4_62 gnd C_wl
Rw5_62 word5_62 word4_62 R_wl
Cwl_5_62 word5_62 gnd C_wl
Rw6_62 word6_62 word5_62 R_wl
Cwl_6_62 word6_62 gnd C_wl
Rw7_62 word7_62 word6_62 R_wl
Cwl_7_62 word7_62 gnd C_wl
Rw8_62 word8_62 word7_62 R_wl
Cwl_8_62 word8_62 gnd C_wl
Rw9_62 word9_62 word8_62 R_wl
Cwl_9_62 word9_62 gnd C_wl
Rw10_62 word10_62 word9_62 R_wl
Cwl_10_62 word10_62 gnd C_wl
Rw11_62 word11_62 word10_62 R_wl
Cwl_11_62 word11_62 gnd C_wl
Rw12_62 word12_62 word11_62 R_wl
Cwl_12_62 word12_62 gnd C_wl
Rw13_62 word13_62 word12_62 R_wl
Cwl_13_62 word13_62 gnd C_wl
Rw14_62 word14_62 word13_62 R_wl
Cwl_14_62 word14_62 gnd C_wl
Rw15_62 word15_62 word14_62 R_wl
Cwl_15_62 word15_62 gnd C_wl
Rw16_62 word16_62 word15_62 R_wl
Cwl_16_62 word16_62 gnd C_wl
Rw17_62 word17_62 word16_62 R_wl
Cwl_17_62 word17_62 gnd C_wl
Rw18_62 word18_62 word17_62 R_wl
Cwl_18_62 word18_62 gnd C_wl
Rw19_62 word19_62 word18_62 R_wl
Cwl_19_62 word19_62 gnd C_wl
Rw20_62 word20_62 word19_62 R_wl
Cwl_20_62 word20_62 gnd C_wl
Rw21_62 word21_62 word20_62 R_wl
Cwl_21_62 word21_62 gnd C_wl
Rw22_62 word22_62 word21_62 R_wl
Cwl_22_62 word22_62 gnd C_wl
Rw23_62 word23_62 word22_62 R_wl
Cwl_23_62 word23_62 gnd C_wl
Rw24_62 word24_62 word23_62 R_wl
Cwl_24_62 word24_62 gnd C_wl
Rw25_62 word25_62 word24_62 R_wl
Cwl_25_62 word25_62 gnd C_wl
Rw26_62 word26_62 word25_62 R_wl
Cwl_26_62 word26_62 gnd C_wl
Rw27_62 word27_62 word26_62 R_wl
Cwl_27_62 word27_62 gnd C_wl
Rw28_62 word28_62 word27_62 R_wl
Cwl_28_62 word28_62 gnd C_wl
Rw29_62 word29_62 word28_62 R_wl
Cwl_29_62 word29_62 gnd C_wl
Rw30_62 word30_62 word29_62 R_wl
Cwl_30_62 word30_62 gnd C_wl
Rw31_62 word31_62 word30_62 R_wl
Cwl_31_62 word31_62 gnd C_wl
Rw32_62 word32_62 word31_62 R_wl
Cwl_32_62 word32_62 gnd C_wl
Rw33_62 word33_62 word32_62 R_wl
Cwl_33_62 word33_62 gnd C_wl
Rw34_62 word34_62 word33_62 R_wl
Cwl_34_62 word34_62 gnd C_wl
Rw35_62 word35_62 word34_62 R_wl
Cwl_35_62 word35_62 gnd C_wl
Rw36_62 word36_62 word35_62 R_wl
Cwl_36_62 word36_62 gnd C_wl
Rw37_62 word37_62 word36_62 R_wl
Cwl_37_62 word37_62 gnd C_wl
Rw38_62 word38_62 word37_62 R_wl
Cwl_38_62 word38_62 gnd C_wl
Rw39_62 word39_62 word38_62 R_wl
Cwl_39_62 word39_62 gnd C_wl
Rw40_62 word40_62 word39_62 R_wl
Cwl_40_62 word40_62 gnd C_wl
Rw41_62 word41_62 word40_62 R_wl
Cwl_41_62 word41_62 gnd C_wl
Rw42_62 word42_62 word41_62 R_wl
Cwl_42_62 word42_62 gnd C_wl
Rw43_62 word43_62 word42_62 R_wl
Cwl_43_62 word43_62 gnd C_wl
Rw44_62 word44_62 word43_62 R_wl
Cwl_44_62 word44_62 gnd C_wl
Rw45_62 word45_62 word44_62 R_wl
Cwl_45_62 word45_62 gnd C_wl
Rw46_62 word46_62 word45_62 R_wl
Cwl_46_62 word46_62 gnd C_wl
Rw47_62 word47_62 word46_62 R_wl
Cwl_47_62 word47_62 gnd C_wl
Rw48_62 word48_62 word47_62 R_wl
Cwl_48_62 word48_62 gnd C_wl
Rw49_62 word49_62 word48_62 R_wl
Cwl_49_62 word49_62 gnd C_wl
Rw50_62 word50_62 word49_62 R_wl
Cwl_50_62 word50_62 gnd C_wl
Rw51_62 word51_62 word50_62 R_wl
Cwl_51_62 word51_62 gnd C_wl
Rw52_62 word52_62 word51_62 R_wl
Cwl_52_62 word52_62 gnd C_wl
Rw53_62 word53_62 word52_62 R_wl
Cwl_53_62 word53_62 gnd C_wl
Rw54_62 word54_62 word53_62 R_wl
Cwl_54_62 word54_62 gnd C_wl
Rw55_62 word55_62 word54_62 R_wl
Cwl_55_62 word55_62 gnd C_wl
Rw56_62 word56_62 word55_62 R_wl
Cwl_56_62 word56_62 gnd C_wl
Rw57_62 word57_62 word56_62 R_wl
Cwl_57_62 word57_62 gnd C_wl
Rw58_62 word58_62 word57_62 R_wl
Cwl_58_62 word58_62 gnd C_wl
Rw59_62 word59_62 word58_62 R_wl
Cwl_59_62 word59_62 gnd C_wl
Rw60_62 word60_62 word59_62 R_wl
Cwl_60_62 word60_62 gnd C_wl
Rw61_62 word61_62 word60_62 R_wl
Cwl_61_62 word61_62 gnd C_wl
Rw62_62 word62_62 word61_62 R_wl
Cwl_62_62 word62_62 gnd C_wl
Rw63_62 word63_62 word62_62 R_wl
Cwl_63_62 word63_62 gnd C_wl
Rw64_62 word64_62 word63_62 R_wl
Cwl_64_62 word64_62 gnd C_wl
Rw65_62 word65_62 word64_62 R_wl
Cwl_65_62 word65_62 gnd C_wl
Rw66_62 word66_62 word65_62 R_wl
Cwl_66_62 word66_62 gnd C_wl
Rw67_62 word67_62 word66_62 R_wl
Cwl_67_62 word67_62 gnd C_wl
Rw68_62 word68_62 word67_62 R_wl
Cwl_68_62 word68_62 gnd C_wl
Rw69_62 word69_62 word68_62 R_wl
Cwl_69_62 word69_62 gnd C_wl
Rw70_62 word70_62 word69_62 R_wl
Cwl_70_62 word70_62 gnd C_wl
Rw71_62 word71_62 word70_62 R_wl
Cwl_71_62 word71_62 gnd C_wl
Rw72_62 word72_62 word71_62 R_wl
Cwl_72_62 word72_62 gnd C_wl
Rw73_62 word73_62 word72_62 R_wl
Cwl_73_62 word73_62 gnd C_wl
Rw74_62 word74_62 word73_62 R_wl
Cwl_74_62 word74_62 gnd C_wl
Rw75_62 word75_62 word74_62 R_wl
Cwl_75_62 word75_62 gnd C_wl
Rw76_62 word76_62 word75_62 R_wl
Cwl_76_62 word76_62 gnd C_wl
Rw77_62 word77_62 word76_62 R_wl
Cwl_77_62 word77_62 gnd C_wl
Rw78_62 word78_62 word77_62 R_wl
Cwl_78_62 word78_62 gnd C_wl
Rw79_62 word79_62 word78_62 R_wl
Cwl_79_62 word79_62 gnd C_wl
Rw80_62 word80_62 word79_62 R_wl
Cwl_80_62 word80_62 gnd C_wl
Rw81_62 word81_62 word80_62 R_wl
Cwl_81_62 word81_62 gnd C_wl
Rw82_62 word82_62 word81_62 R_wl
Cwl_82_62 word82_62 gnd C_wl
Rw83_62 word83_62 word82_62 R_wl
Cwl_83_62 word83_62 gnd C_wl
Rw84_62 word84_62 word83_62 R_wl
Cwl_84_62 word84_62 gnd C_wl
Rw85_62 word85_62 word84_62 R_wl
Cwl_85_62 word85_62 gnd C_wl
Rw86_62 word86_62 word85_62 R_wl
Cwl_86_62 word86_62 gnd C_wl
Rw87_62 word87_62 word86_62 R_wl
Cwl_87_62 word87_62 gnd C_wl
Rw88_62 word88_62 word87_62 R_wl
Cwl_88_62 word88_62 gnd C_wl
Rw89_62 word89_62 word88_62 R_wl
Cwl_89_62 word89_62 gnd C_wl
Rw90_62 word90_62 word89_62 R_wl
Cwl_90_62 word90_62 gnd C_wl
Rw91_62 word91_62 word90_62 R_wl
Cwl_91_62 word91_62 gnd C_wl
Rw92_62 word92_62 word91_62 R_wl
Cwl_92_62 word92_62 gnd C_wl
Rw93_62 word93_62 word92_62 R_wl
Cwl_93_62 word93_62 gnd C_wl
Rw94_62 word94_62 word93_62 R_wl
Cwl_94_62 word94_62 gnd C_wl
Rw95_62 word95_62 word94_62 R_wl
Cwl_95_62 word95_62 gnd C_wl
Rw96_62 word96_62 word95_62 R_wl
Cwl_96_62 word96_62 gnd C_wl
Rw97_62 word97_62 word96_62 R_wl
Cwl_97_62 word97_62 gnd C_wl
Rw98_62 word98_62 word97_62 R_wl
Cwl_98_62 word98_62 gnd C_wl
Rw99_62 word99_62 word98_62 R_wl
Cwl_99_62 word99_62 gnd C_wl
Vwl_63 word_63 0 0
Rw0_63 word_63 word0_63 R_wl
Cwl_0_63 word0_63 gnd C_wl
Rw1_63 word1_63 word0_63 R_wl
Cwl_1_63 word1_63 gnd C_wl
Rw2_63 word2_63 word1_63 R_wl
Cwl_2_63 word2_63 gnd C_wl
Rw3_63 word3_63 word2_63 R_wl
Cwl_3_63 word3_63 gnd C_wl
Rw4_63 word4_63 word3_63 R_wl
Cwl_4_63 word4_63 gnd C_wl
Rw5_63 word5_63 word4_63 R_wl
Cwl_5_63 word5_63 gnd C_wl
Rw6_63 word6_63 word5_63 R_wl
Cwl_6_63 word6_63 gnd C_wl
Rw7_63 word7_63 word6_63 R_wl
Cwl_7_63 word7_63 gnd C_wl
Rw8_63 word8_63 word7_63 R_wl
Cwl_8_63 word8_63 gnd C_wl
Rw9_63 word9_63 word8_63 R_wl
Cwl_9_63 word9_63 gnd C_wl
Rw10_63 word10_63 word9_63 R_wl
Cwl_10_63 word10_63 gnd C_wl
Rw11_63 word11_63 word10_63 R_wl
Cwl_11_63 word11_63 gnd C_wl
Rw12_63 word12_63 word11_63 R_wl
Cwl_12_63 word12_63 gnd C_wl
Rw13_63 word13_63 word12_63 R_wl
Cwl_13_63 word13_63 gnd C_wl
Rw14_63 word14_63 word13_63 R_wl
Cwl_14_63 word14_63 gnd C_wl
Rw15_63 word15_63 word14_63 R_wl
Cwl_15_63 word15_63 gnd C_wl
Rw16_63 word16_63 word15_63 R_wl
Cwl_16_63 word16_63 gnd C_wl
Rw17_63 word17_63 word16_63 R_wl
Cwl_17_63 word17_63 gnd C_wl
Rw18_63 word18_63 word17_63 R_wl
Cwl_18_63 word18_63 gnd C_wl
Rw19_63 word19_63 word18_63 R_wl
Cwl_19_63 word19_63 gnd C_wl
Rw20_63 word20_63 word19_63 R_wl
Cwl_20_63 word20_63 gnd C_wl
Rw21_63 word21_63 word20_63 R_wl
Cwl_21_63 word21_63 gnd C_wl
Rw22_63 word22_63 word21_63 R_wl
Cwl_22_63 word22_63 gnd C_wl
Rw23_63 word23_63 word22_63 R_wl
Cwl_23_63 word23_63 gnd C_wl
Rw24_63 word24_63 word23_63 R_wl
Cwl_24_63 word24_63 gnd C_wl
Rw25_63 word25_63 word24_63 R_wl
Cwl_25_63 word25_63 gnd C_wl
Rw26_63 word26_63 word25_63 R_wl
Cwl_26_63 word26_63 gnd C_wl
Rw27_63 word27_63 word26_63 R_wl
Cwl_27_63 word27_63 gnd C_wl
Rw28_63 word28_63 word27_63 R_wl
Cwl_28_63 word28_63 gnd C_wl
Rw29_63 word29_63 word28_63 R_wl
Cwl_29_63 word29_63 gnd C_wl
Rw30_63 word30_63 word29_63 R_wl
Cwl_30_63 word30_63 gnd C_wl
Rw31_63 word31_63 word30_63 R_wl
Cwl_31_63 word31_63 gnd C_wl
Rw32_63 word32_63 word31_63 R_wl
Cwl_32_63 word32_63 gnd C_wl
Rw33_63 word33_63 word32_63 R_wl
Cwl_33_63 word33_63 gnd C_wl
Rw34_63 word34_63 word33_63 R_wl
Cwl_34_63 word34_63 gnd C_wl
Rw35_63 word35_63 word34_63 R_wl
Cwl_35_63 word35_63 gnd C_wl
Rw36_63 word36_63 word35_63 R_wl
Cwl_36_63 word36_63 gnd C_wl
Rw37_63 word37_63 word36_63 R_wl
Cwl_37_63 word37_63 gnd C_wl
Rw38_63 word38_63 word37_63 R_wl
Cwl_38_63 word38_63 gnd C_wl
Rw39_63 word39_63 word38_63 R_wl
Cwl_39_63 word39_63 gnd C_wl
Rw40_63 word40_63 word39_63 R_wl
Cwl_40_63 word40_63 gnd C_wl
Rw41_63 word41_63 word40_63 R_wl
Cwl_41_63 word41_63 gnd C_wl
Rw42_63 word42_63 word41_63 R_wl
Cwl_42_63 word42_63 gnd C_wl
Rw43_63 word43_63 word42_63 R_wl
Cwl_43_63 word43_63 gnd C_wl
Rw44_63 word44_63 word43_63 R_wl
Cwl_44_63 word44_63 gnd C_wl
Rw45_63 word45_63 word44_63 R_wl
Cwl_45_63 word45_63 gnd C_wl
Rw46_63 word46_63 word45_63 R_wl
Cwl_46_63 word46_63 gnd C_wl
Rw47_63 word47_63 word46_63 R_wl
Cwl_47_63 word47_63 gnd C_wl
Rw48_63 word48_63 word47_63 R_wl
Cwl_48_63 word48_63 gnd C_wl
Rw49_63 word49_63 word48_63 R_wl
Cwl_49_63 word49_63 gnd C_wl
Rw50_63 word50_63 word49_63 R_wl
Cwl_50_63 word50_63 gnd C_wl
Rw51_63 word51_63 word50_63 R_wl
Cwl_51_63 word51_63 gnd C_wl
Rw52_63 word52_63 word51_63 R_wl
Cwl_52_63 word52_63 gnd C_wl
Rw53_63 word53_63 word52_63 R_wl
Cwl_53_63 word53_63 gnd C_wl
Rw54_63 word54_63 word53_63 R_wl
Cwl_54_63 word54_63 gnd C_wl
Rw55_63 word55_63 word54_63 R_wl
Cwl_55_63 word55_63 gnd C_wl
Rw56_63 word56_63 word55_63 R_wl
Cwl_56_63 word56_63 gnd C_wl
Rw57_63 word57_63 word56_63 R_wl
Cwl_57_63 word57_63 gnd C_wl
Rw58_63 word58_63 word57_63 R_wl
Cwl_58_63 word58_63 gnd C_wl
Rw59_63 word59_63 word58_63 R_wl
Cwl_59_63 word59_63 gnd C_wl
Rw60_63 word60_63 word59_63 R_wl
Cwl_60_63 word60_63 gnd C_wl
Rw61_63 word61_63 word60_63 R_wl
Cwl_61_63 word61_63 gnd C_wl
Rw62_63 word62_63 word61_63 R_wl
Cwl_62_63 word62_63 gnd C_wl
Rw63_63 word63_63 word62_63 R_wl
Cwl_63_63 word63_63 gnd C_wl
Rw64_63 word64_63 word63_63 R_wl
Cwl_64_63 word64_63 gnd C_wl
Rw65_63 word65_63 word64_63 R_wl
Cwl_65_63 word65_63 gnd C_wl
Rw66_63 word66_63 word65_63 R_wl
Cwl_66_63 word66_63 gnd C_wl
Rw67_63 word67_63 word66_63 R_wl
Cwl_67_63 word67_63 gnd C_wl
Rw68_63 word68_63 word67_63 R_wl
Cwl_68_63 word68_63 gnd C_wl
Rw69_63 word69_63 word68_63 R_wl
Cwl_69_63 word69_63 gnd C_wl
Rw70_63 word70_63 word69_63 R_wl
Cwl_70_63 word70_63 gnd C_wl
Rw71_63 word71_63 word70_63 R_wl
Cwl_71_63 word71_63 gnd C_wl
Rw72_63 word72_63 word71_63 R_wl
Cwl_72_63 word72_63 gnd C_wl
Rw73_63 word73_63 word72_63 R_wl
Cwl_73_63 word73_63 gnd C_wl
Rw74_63 word74_63 word73_63 R_wl
Cwl_74_63 word74_63 gnd C_wl
Rw75_63 word75_63 word74_63 R_wl
Cwl_75_63 word75_63 gnd C_wl
Rw76_63 word76_63 word75_63 R_wl
Cwl_76_63 word76_63 gnd C_wl
Rw77_63 word77_63 word76_63 R_wl
Cwl_77_63 word77_63 gnd C_wl
Rw78_63 word78_63 word77_63 R_wl
Cwl_78_63 word78_63 gnd C_wl
Rw79_63 word79_63 word78_63 R_wl
Cwl_79_63 word79_63 gnd C_wl
Rw80_63 word80_63 word79_63 R_wl
Cwl_80_63 word80_63 gnd C_wl
Rw81_63 word81_63 word80_63 R_wl
Cwl_81_63 word81_63 gnd C_wl
Rw82_63 word82_63 word81_63 R_wl
Cwl_82_63 word82_63 gnd C_wl
Rw83_63 word83_63 word82_63 R_wl
Cwl_83_63 word83_63 gnd C_wl
Rw84_63 word84_63 word83_63 R_wl
Cwl_84_63 word84_63 gnd C_wl
Rw85_63 word85_63 word84_63 R_wl
Cwl_85_63 word85_63 gnd C_wl
Rw86_63 word86_63 word85_63 R_wl
Cwl_86_63 word86_63 gnd C_wl
Rw87_63 word87_63 word86_63 R_wl
Cwl_87_63 word87_63 gnd C_wl
Rw88_63 word88_63 word87_63 R_wl
Cwl_88_63 word88_63 gnd C_wl
Rw89_63 word89_63 word88_63 R_wl
Cwl_89_63 word89_63 gnd C_wl
Rw90_63 word90_63 word89_63 R_wl
Cwl_90_63 word90_63 gnd C_wl
Rw91_63 word91_63 word90_63 R_wl
Cwl_91_63 word91_63 gnd C_wl
Rw92_63 word92_63 word91_63 R_wl
Cwl_92_63 word92_63 gnd C_wl
Rw93_63 word93_63 word92_63 R_wl
Cwl_93_63 word93_63 gnd C_wl
Rw94_63 word94_63 word93_63 R_wl
Cwl_94_63 word94_63 gnd C_wl
Rw95_63 word95_63 word94_63 R_wl
Cwl_95_63 word95_63 gnd C_wl
Rw96_63 word96_63 word95_63 R_wl
Cwl_96_63 word96_63 gnd C_wl
Rw97_63 word97_63 word96_63 R_wl
Cwl_97_63 word97_63 gnd C_wl
Rw98_63 word98_63 word97_63 R_wl
Cwl_98_63 word98_63 gnd C_wl
Rw99_63 word99_63 word98_63 R_wl
Cwl_99_63 word99_63 gnd C_wl
Vwl_64 word_64 0 0
Rw0_64 word_64 word0_64 R_wl
Cwl_0_64 word0_64 gnd C_wl
Rw1_64 word1_64 word0_64 R_wl
Cwl_1_64 word1_64 gnd C_wl
Rw2_64 word2_64 word1_64 R_wl
Cwl_2_64 word2_64 gnd C_wl
Rw3_64 word3_64 word2_64 R_wl
Cwl_3_64 word3_64 gnd C_wl
Rw4_64 word4_64 word3_64 R_wl
Cwl_4_64 word4_64 gnd C_wl
Rw5_64 word5_64 word4_64 R_wl
Cwl_5_64 word5_64 gnd C_wl
Rw6_64 word6_64 word5_64 R_wl
Cwl_6_64 word6_64 gnd C_wl
Rw7_64 word7_64 word6_64 R_wl
Cwl_7_64 word7_64 gnd C_wl
Rw8_64 word8_64 word7_64 R_wl
Cwl_8_64 word8_64 gnd C_wl
Rw9_64 word9_64 word8_64 R_wl
Cwl_9_64 word9_64 gnd C_wl
Rw10_64 word10_64 word9_64 R_wl
Cwl_10_64 word10_64 gnd C_wl
Rw11_64 word11_64 word10_64 R_wl
Cwl_11_64 word11_64 gnd C_wl
Rw12_64 word12_64 word11_64 R_wl
Cwl_12_64 word12_64 gnd C_wl
Rw13_64 word13_64 word12_64 R_wl
Cwl_13_64 word13_64 gnd C_wl
Rw14_64 word14_64 word13_64 R_wl
Cwl_14_64 word14_64 gnd C_wl
Rw15_64 word15_64 word14_64 R_wl
Cwl_15_64 word15_64 gnd C_wl
Rw16_64 word16_64 word15_64 R_wl
Cwl_16_64 word16_64 gnd C_wl
Rw17_64 word17_64 word16_64 R_wl
Cwl_17_64 word17_64 gnd C_wl
Rw18_64 word18_64 word17_64 R_wl
Cwl_18_64 word18_64 gnd C_wl
Rw19_64 word19_64 word18_64 R_wl
Cwl_19_64 word19_64 gnd C_wl
Rw20_64 word20_64 word19_64 R_wl
Cwl_20_64 word20_64 gnd C_wl
Rw21_64 word21_64 word20_64 R_wl
Cwl_21_64 word21_64 gnd C_wl
Rw22_64 word22_64 word21_64 R_wl
Cwl_22_64 word22_64 gnd C_wl
Rw23_64 word23_64 word22_64 R_wl
Cwl_23_64 word23_64 gnd C_wl
Rw24_64 word24_64 word23_64 R_wl
Cwl_24_64 word24_64 gnd C_wl
Rw25_64 word25_64 word24_64 R_wl
Cwl_25_64 word25_64 gnd C_wl
Rw26_64 word26_64 word25_64 R_wl
Cwl_26_64 word26_64 gnd C_wl
Rw27_64 word27_64 word26_64 R_wl
Cwl_27_64 word27_64 gnd C_wl
Rw28_64 word28_64 word27_64 R_wl
Cwl_28_64 word28_64 gnd C_wl
Rw29_64 word29_64 word28_64 R_wl
Cwl_29_64 word29_64 gnd C_wl
Rw30_64 word30_64 word29_64 R_wl
Cwl_30_64 word30_64 gnd C_wl
Rw31_64 word31_64 word30_64 R_wl
Cwl_31_64 word31_64 gnd C_wl
Rw32_64 word32_64 word31_64 R_wl
Cwl_32_64 word32_64 gnd C_wl
Rw33_64 word33_64 word32_64 R_wl
Cwl_33_64 word33_64 gnd C_wl
Rw34_64 word34_64 word33_64 R_wl
Cwl_34_64 word34_64 gnd C_wl
Rw35_64 word35_64 word34_64 R_wl
Cwl_35_64 word35_64 gnd C_wl
Rw36_64 word36_64 word35_64 R_wl
Cwl_36_64 word36_64 gnd C_wl
Rw37_64 word37_64 word36_64 R_wl
Cwl_37_64 word37_64 gnd C_wl
Rw38_64 word38_64 word37_64 R_wl
Cwl_38_64 word38_64 gnd C_wl
Rw39_64 word39_64 word38_64 R_wl
Cwl_39_64 word39_64 gnd C_wl
Rw40_64 word40_64 word39_64 R_wl
Cwl_40_64 word40_64 gnd C_wl
Rw41_64 word41_64 word40_64 R_wl
Cwl_41_64 word41_64 gnd C_wl
Rw42_64 word42_64 word41_64 R_wl
Cwl_42_64 word42_64 gnd C_wl
Rw43_64 word43_64 word42_64 R_wl
Cwl_43_64 word43_64 gnd C_wl
Rw44_64 word44_64 word43_64 R_wl
Cwl_44_64 word44_64 gnd C_wl
Rw45_64 word45_64 word44_64 R_wl
Cwl_45_64 word45_64 gnd C_wl
Rw46_64 word46_64 word45_64 R_wl
Cwl_46_64 word46_64 gnd C_wl
Rw47_64 word47_64 word46_64 R_wl
Cwl_47_64 word47_64 gnd C_wl
Rw48_64 word48_64 word47_64 R_wl
Cwl_48_64 word48_64 gnd C_wl
Rw49_64 word49_64 word48_64 R_wl
Cwl_49_64 word49_64 gnd C_wl
Rw50_64 word50_64 word49_64 R_wl
Cwl_50_64 word50_64 gnd C_wl
Rw51_64 word51_64 word50_64 R_wl
Cwl_51_64 word51_64 gnd C_wl
Rw52_64 word52_64 word51_64 R_wl
Cwl_52_64 word52_64 gnd C_wl
Rw53_64 word53_64 word52_64 R_wl
Cwl_53_64 word53_64 gnd C_wl
Rw54_64 word54_64 word53_64 R_wl
Cwl_54_64 word54_64 gnd C_wl
Rw55_64 word55_64 word54_64 R_wl
Cwl_55_64 word55_64 gnd C_wl
Rw56_64 word56_64 word55_64 R_wl
Cwl_56_64 word56_64 gnd C_wl
Rw57_64 word57_64 word56_64 R_wl
Cwl_57_64 word57_64 gnd C_wl
Rw58_64 word58_64 word57_64 R_wl
Cwl_58_64 word58_64 gnd C_wl
Rw59_64 word59_64 word58_64 R_wl
Cwl_59_64 word59_64 gnd C_wl
Rw60_64 word60_64 word59_64 R_wl
Cwl_60_64 word60_64 gnd C_wl
Rw61_64 word61_64 word60_64 R_wl
Cwl_61_64 word61_64 gnd C_wl
Rw62_64 word62_64 word61_64 R_wl
Cwl_62_64 word62_64 gnd C_wl
Rw63_64 word63_64 word62_64 R_wl
Cwl_63_64 word63_64 gnd C_wl
Rw64_64 word64_64 word63_64 R_wl
Cwl_64_64 word64_64 gnd C_wl
Rw65_64 word65_64 word64_64 R_wl
Cwl_65_64 word65_64 gnd C_wl
Rw66_64 word66_64 word65_64 R_wl
Cwl_66_64 word66_64 gnd C_wl
Rw67_64 word67_64 word66_64 R_wl
Cwl_67_64 word67_64 gnd C_wl
Rw68_64 word68_64 word67_64 R_wl
Cwl_68_64 word68_64 gnd C_wl
Rw69_64 word69_64 word68_64 R_wl
Cwl_69_64 word69_64 gnd C_wl
Rw70_64 word70_64 word69_64 R_wl
Cwl_70_64 word70_64 gnd C_wl
Rw71_64 word71_64 word70_64 R_wl
Cwl_71_64 word71_64 gnd C_wl
Rw72_64 word72_64 word71_64 R_wl
Cwl_72_64 word72_64 gnd C_wl
Rw73_64 word73_64 word72_64 R_wl
Cwl_73_64 word73_64 gnd C_wl
Rw74_64 word74_64 word73_64 R_wl
Cwl_74_64 word74_64 gnd C_wl
Rw75_64 word75_64 word74_64 R_wl
Cwl_75_64 word75_64 gnd C_wl
Rw76_64 word76_64 word75_64 R_wl
Cwl_76_64 word76_64 gnd C_wl
Rw77_64 word77_64 word76_64 R_wl
Cwl_77_64 word77_64 gnd C_wl
Rw78_64 word78_64 word77_64 R_wl
Cwl_78_64 word78_64 gnd C_wl
Rw79_64 word79_64 word78_64 R_wl
Cwl_79_64 word79_64 gnd C_wl
Rw80_64 word80_64 word79_64 R_wl
Cwl_80_64 word80_64 gnd C_wl
Rw81_64 word81_64 word80_64 R_wl
Cwl_81_64 word81_64 gnd C_wl
Rw82_64 word82_64 word81_64 R_wl
Cwl_82_64 word82_64 gnd C_wl
Rw83_64 word83_64 word82_64 R_wl
Cwl_83_64 word83_64 gnd C_wl
Rw84_64 word84_64 word83_64 R_wl
Cwl_84_64 word84_64 gnd C_wl
Rw85_64 word85_64 word84_64 R_wl
Cwl_85_64 word85_64 gnd C_wl
Rw86_64 word86_64 word85_64 R_wl
Cwl_86_64 word86_64 gnd C_wl
Rw87_64 word87_64 word86_64 R_wl
Cwl_87_64 word87_64 gnd C_wl
Rw88_64 word88_64 word87_64 R_wl
Cwl_88_64 word88_64 gnd C_wl
Rw89_64 word89_64 word88_64 R_wl
Cwl_89_64 word89_64 gnd C_wl
Rw90_64 word90_64 word89_64 R_wl
Cwl_90_64 word90_64 gnd C_wl
Rw91_64 word91_64 word90_64 R_wl
Cwl_91_64 word91_64 gnd C_wl
Rw92_64 word92_64 word91_64 R_wl
Cwl_92_64 word92_64 gnd C_wl
Rw93_64 word93_64 word92_64 R_wl
Cwl_93_64 word93_64 gnd C_wl
Rw94_64 word94_64 word93_64 R_wl
Cwl_94_64 word94_64 gnd C_wl
Rw95_64 word95_64 word94_64 R_wl
Cwl_95_64 word95_64 gnd C_wl
Rw96_64 word96_64 word95_64 R_wl
Cwl_96_64 word96_64 gnd C_wl
Rw97_64 word97_64 word96_64 R_wl
Cwl_97_64 word97_64 gnd C_wl
Rw98_64 word98_64 word97_64 R_wl
Cwl_98_64 word98_64 gnd C_wl
Rw99_64 word99_64 word98_64 R_wl
Cwl_99_64 word99_64 gnd C_wl
Vwl_65 word_65 0 0
Rw0_65 word_65 word0_65 R_wl
Cwl_0_65 word0_65 gnd C_wl
Rw1_65 word1_65 word0_65 R_wl
Cwl_1_65 word1_65 gnd C_wl
Rw2_65 word2_65 word1_65 R_wl
Cwl_2_65 word2_65 gnd C_wl
Rw3_65 word3_65 word2_65 R_wl
Cwl_3_65 word3_65 gnd C_wl
Rw4_65 word4_65 word3_65 R_wl
Cwl_4_65 word4_65 gnd C_wl
Rw5_65 word5_65 word4_65 R_wl
Cwl_5_65 word5_65 gnd C_wl
Rw6_65 word6_65 word5_65 R_wl
Cwl_6_65 word6_65 gnd C_wl
Rw7_65 word7_65 word6_65 R_wl
Cwl_7_65 word7_65 gnd C_wl
Rw8_65 word8_65 word7_65 R_wl
Cwl_8_65 word8_65 gnd C_wl
Rw9_65 word9_65 word8_65 R_wl
Cwl_9_65 word9_65 gnd C_wl
Rw10_65 word10_65 word9_65 R_wl
Cwl_10_65 word10_65 gnd C_wl
Rw11_65 word11_65 word10_65 R_wl
Cwl_11_65 word11_65 gnd C_wl
Rw12_65 word12_65 word11_65 R_wl
Cwl_12_65 word12_65 gnd C_wl
Rw13_65 word13_65 word12_65 R_wl
Cwl_13_65 word13_65 gnd C_wl
Rw14_65 word14_65 word13_65 R_wl
Cwl_14_65 word14_65 gnd C_wl
Rw15_65 word15_65 word14_65 R_wl
Cwl_15_65 word15_65 gnd C_wl
Rw16_65 word16_65 word15_65 R_wl
Cwl_16_65 word16_65 gnd C_wl
Rw17_65 word17_65 word16_65 R_wl
Cwl_17_65 word17_65 gnd C_wl
Rw18_65 word18_65 word17_65 R_wl
Cwl_18_65 word18_65 gnd C_wl
Rw19_65 word19_65 word18_65 R_wl
Cwl_19_65 word19_65 gnd C_wl
Rw20_65 word20_65 word19_65 R_wl
Cwl_20_65 word20_65 gnd C_wl
Rw21_65 word21_65 word20_65 R_wl
Cwl_21_65 word21_65 gnd C_wl
Rw22_65 word22_65 word21_65 R_wl
Cwl_22_65 word22_65 gnd C_wl
Rw23_65 word23_65 word22_65 R_wl
Cwl_23_65 word23_65 gnd C_wl
Rw24_65 word24_65 word23_65 R_wl
Cwl_24_65 word24_65 gnd C_wl
Rw25_65 word25_65 word24_65 R_wl
Cwl_25_65 word25_65 gnd C_wl
Rw26_65 word26_65 word25_65 R_wl
Cwl_26_65 word26_65 gnd C_wl
Rw27_65 word27_65 word26_65 R_wl
Cwl_27_65 word27_65 gnd C_wl
Rw28_65 word28_65 word27_65 R_wl
Cwl_28_65 word28_65 gnd C_wl
Rw29_65 word29_65 word28_65 R_wl
Cwl_29_65 word29_65 gnd C_wl
Rw30_65 word30_65 word29_65 R_wl
Cwl_30_65 word30_65 gnd C_wl
Rw31_65 word31_65 word30_65 R_wl
Cwl_31_65 word31_65 gnd C_wl
Rw32_65 word32_65 word31_65 R_wl
Cwl_32_65 word32_65 gnd C_wl
Rw33_65 word33_65 word32_65 R_wl
Cwl_33_65 word33_65 gnd C_wl
Rw34_65 word34_65 word33_65 R_wl
Cwl_34_65 word34_65 gnd C_wl
Rw35_65 word35_65 word34_65 R_wl
Cwl_35_65 word35_65 gnd C_wl
Rw36_65 word36_65 word35_65 R_wl
Cwl_36_65 word36_65 gnd C_wl
Rw37_65 word37_65 word36_65 R_wl
Cwl_37_65 word37_65 gnd C_wl
Rw38_65 word38_65 word37_65 R_wl
Cwl_38_65 word38_65 gnd C_wl
Rw39_65 word39_65 word38_65 R_wl
Cwl_39_65 word39_65 gnd C_wl
Rw40_65 word40_65 word39_65 R_wl
Cwl_40_65 word40_65 gnd C_wl
Rw41_65 word41_65 word40_65 R_wl
Cwl_41_65 word41_65 gnd C_wl
Rw42_65 word42_65 word41_65 R_wl
Cwl_42_65 word42_65 gnd C_wl
Rw43_65 word43_65 word42_65 R_wl
Cwl_43_65 word43_65 gnd C_wl
Rw44_65 word44_65 word43_65 R_wl
Cwl_44_65 word44_65 gnd C_wl
Rw45_65 word45_65 word44_65 R_wl
Cwl_45_65 word45_65 gnd C_wl
Rw46_65 word46_65 word45_65 R_wl
Cwl_46_65 word46_65 gnd C_wl
Rw47_65 word47_65 word46_65 R_wl
Cwl_47_65 word47_65 gnd C_wl
Rw48_65 word48_65 word47_65 R_wl
Cwl_48_65 word48_65 gnd C_wl
Rw49_65 word49_65 word48_65 R_wl
Cwl_49_65 word49_65 gnd C_wl
Rw50_65 word50_65 word49_65 R_wl
Cwl_50_65 word50_65 gnd C_wl
Rw51_65 word51_65 word50_65 R_wl
Cwl_51_65 word51_65 gnd C_wl
Rw52_65 word52_65 word51_65 R_wl
Cwl_52_65 word52_65 gnd C_wl
Rw53_65 word53_65 word52_65 R_wl
Cwl_53_65 word53_65 gnd C_wl
Rw54_65 word54_65 word53_65 R_wl
Cwl_54_65 word54_65 gnd C_wl
Rw55_65 word55_65 word54_65 R_wl
Cwl_55_65 word55_65 gnd C_wl
Rw56_65 word56_65 word55_65 R_wl
Cwl_56_65 word56_65 gnd C_wl
Rw57_65 word57_65 word56_65 R_wl
Cwl_57_65 word57_65 gnd C_wl
Rw58_65 word58_65 word57_65 R_wl
Cwl_58_65 word58_65 gnd C_wl
Rw59_65 word59_65 word58_65 R_wl
Cwl_59_65 word59_65 gnd C_wl
Rw60_65 word60_65 word59_65 R_wl
Cwl_60_65 word60_65 gnd C_wl
Rw61_65 word61_65 word60_65 R_wl
Cwl_61_65 word61_65 gnd C_wl
Rw62_65 word62_65 word61_65 R_wl
Cwl_62_65 word62_65 gnd C_wl
Rw63_65 word63_65 word62_65 R_wl
Cwl_63_65 word63_65 gnd C_wl
Rw64_65 word64_65 word63_65 R_wl
Cwl_64_65 word64_65 gnd C_wl
Rw65_65 word65_65 word64_65 R_wl
Cwl_65_65 word65_65 gnd C_wl
Rw66_65 word66_65 word65_65 R_wl
Cwl_66_65 word66_65 gnd C_wl
Rw67_65 word67_65 word66_65 R_wl
Cwl_67_65 word67_65 gnd C_wl
Rw68_65 word68_65 word67_65 R_wl
Cwl_68_65 word68_65 gnd C_wl
Rw69_65 word69_65 word68_65 R_wl
Cwl_69_65 word69_65 gnd C_wl
Rw70_65 word70_65 word69_65 R_wl
Cwl_70_65 word70_65 gnd C_wl
Rw71_65 word71_65 word70_65 R_wl
Cwl_71_65 word71_65 gnd C_wl
Rw72_65 word72_65 word71_65 R_wl
Cwl_72_65 word72_65 gnd C_wl
Rw73_65 word73_65 word72_65 R_wl
Cwl_73_65 word73_65 gnd C_wl
Rw74_65 word74_65 word73_65 R_wl
Cwl_74_65 word74_65 gnd C_wl
Rw75_65 word75_65 word74_65 R_wl
Cwl_75_65 word75_65 gnd C_wl
Rw76_65 word76_65 word75_65 R_wl
Cwl_76_65 word76_65 gnd C_wl
Rw77_65 word77_65 word76_65 R_wl
Cwl_77_65 word77_65 gnd C_wl
Rw78_65 word78_65 word77_65 R_wl
Cwl_78_65 word78_65 gnd C_wl
Rw79_65 word79_65 word78_65 R_wl
Cwl_79_65 word79_65 gnd C_wl
Rw80_65 word80_65 word79_65 R_wl
Cwl_80_65 word80_65 gnd C_wl
Rw81_65 word81_65 word80_65 R_wl
Cwl_81_65 word81_65 gnd C_wl
Rw82_65 word82_65 word81_65 R_wl
Cwl_82_65 word82_65 gnd C_wl
Rw83_65 word83_65 word82_65 R_wl
Cwl_83_65 word83_65 gnd C_wl
Rw84_65 word84_65 word83_65 R_wl
Cwl_84_65 word84_65 gnd C_wl
Rw85_65 word85_65 word84_65 R_wl
Cwl_85_65 word85_65 gnd C_wl
Rw86_65 word86_65 word85_65 R_wl
Cwl_86_65 word86_65 gnd C_wl
Rw87_65 word87_65 word86_65 R_wl
Cwl_87_65 word87_65 gnd C_wl
Rw88_65 word88_65 word87_65 R_wl
Cwl_88_65 word88_65 gnd C_wl
Rw89_65 word89_65 word88_65 R_wl
Cwl_89_65 word89_65 gnd C_wl
Rw90_65 word90_65 word89_65 R_wl
Cwl_90_65 word90_65 gnd C_wl
Rw91_65 word91_65 word90_65 R_wl
Cwl_91_65 word91_65 gnd C_wl
Rw92_65 word92_65 word91_65 R_wl
Cwl_92_65 word92_65 gnd C_wl
Rw93_65 word93_65 word92_65 R_wl
Cwl_93_65 word93_65 gnd C_wl
Rw94_65 word94_65 word93_65 R_wl
Cwl_94_65 word94_65 gnd C_wl
Rw95_65 word95_65 word94_65 R_wl
Cwl_95_65 word95_65 gnd C_wl
Rw96_65 word96_65 word95_65 R_wl
Cwl_96_65 word96_65 gnd C_wl
Rw97_65 word97_65 word96_65 R_wl
Cwl_97_65 word97_65 gnd C_wl
Rw98_65 word98_65 word97_65 R_wl
Cwl_98_65 word98_65 gnd C_wl
Rw99_65 word99_65 word98_65 R_wl
Cwl_99_65 word99_65 gnd C_wl
Vwl_66 word_66 0 0
Rw0_66 word_66 word0_66 R_wl
Cwl_0_66 word0_66 gnd C_wl
Rw1_66 word1_66 word0_66 R_wl
Cwl_1_66 word1_66 gnd C_wl
Rw2_66 word2_66 word1_66 R_wl
Cwl_2_66 word2_66 gnd C_wl
Rw3_66 word3_66 word2_66 R_wl
Cwl_3_66 word3_66 gnd C_wl
Rw4_66 word4_66 word3_66 R_wl
Cwl_4_66 word4_66 gnd C_wl
Rw5_66 word5_66 word4_66 R_wl
Cwl_5_66 word5_66 gnd C_wl
Rw6_66 word6_66 word5_66 R_wl
Cwl_6_66 word6_66 gnd C_wl
Rw7_66 word7_66 word6_66 R_wl
Cwl_7_66 word7_66 gnd C_wl
Rw8_66 word8_66 word7_66 R_wl
Cwl_8_66 word8_66 gnd C_wl
Rw9_66 word9_66 word8_66 R_wl
Cwl_9_66 word9_66 gnd C_wl
Rw10_66 word10_66 word9_66 R_wl
Cwl_10_66 word10_66 gnd C_wl
Rw11_66 word11_66 word10_66 R_wl
Cwl_11_66 word11_66 gnd C_wl
Rw12_66 word12_66 word11_66 R_wl
Cwl_12_66 word12_66 gnd C_wl
Rw13_66 word13_66 word12_66 R_wl
Cwl_13_66 word13_66 gnd C_wl
Rw14_66 word14_66 word13_66 R_wl
Cwl_14_66 word14_66 gnd C_wl
Rw15_66 word15_66 word14_66 R_wl
Cwl_15_66 word15_66 gnd C_wl
Rw16_66 word16_66 word15_66 R_wl
Cwl_16_66 word16_66 gnd C_wl
Rw17_66 word17_66 word16_66 R_wl
Cwl_17_66 word17_66 gnd C_wl
Rw18_66 word18_66 word17_66 R_wl
Cwl_18_66 word18_66 gnd C_wl
Rw19_66 word19_66 word18_66 R_wl
Cwl_19_66 word19_66 gnd C_wl
Rw20_66 word20_66 word19_66 R_wl
Cwl_20_66 word20_66 gnd C_wl
Rw21_66 word21_66 word20_66 R_wl
Cwl_21_66 word21_66 gnd C_wl
Rw22_66 word22_66 word21_66 R_wl
Cwl_22_66 word22_66 gnd C_wl
Rw23_66 word23_66 word22_66 R_wl
Cwl_23_66 word23_66 gnd C_wl
Rw24_66 word24_66 word23_66 R_wl
Cwl_24_66 word24_66 gnd C_wl
Rw25_66 word25_66 word24_66 R_wl
Cwl_25_66 word25_66 gnd C_wl
Rw26_66 word26_66 word25_66 R_wl
Cwl_26_66 word26_66 gnd C_wl
Rw27_66 word27_66 word26_66 R_wl
Cwl_27_66 word27_66 gnd C_wl
Rw28_66 word28_66 word27_66 R_wl
Cwl_28_66 word28_66 gnd C_wl
Rw29_66 word29_66 word28_66 R_wl
Cwl_29_66 word29_66 gnd C_wl
Rw30_66 word30_66 word29_66 R_wl
Cwl_30_66 word30_66 gnd C_wl
Rw31_66 word31_66 word30_66 R_wl
Cwl_31_66 word31_66 gnd C_wl
Rw32_66 word32_66 word31_66 R_wl
Cwl_32_66 word32_66 gnd C_wl
Rw33_66 word33_66 word32_66 R_wl
Cwl_33_66 word33_66 gnd C_wl
Rw34_66 word34_66 word33_66 R_wl
Cwl_34_66 word34_66 gnd C_wl
Rw35_66 word35_66 word34_66 R_wl
Cwl_35_66 word35_66 gnd C_wl
Rw36_66 word36_66 word35_66 R_wl
Cwl_36_66 word36_66 gnd C_wl
Rw37_66 word37_66 word36_66 R_wl
Cwl_37_66 word37_66 gnd C_wl
Rw38_66 word38_66 word37_66 R_wl
Cwl_38_66 word38_66 gnd C_wl
Rw39_66 word39_66 word38_66 R_wl
Cwl_39_66 word39_66 gnd C_wl
Rw40_66 word40_66 word39_66 R_wl
Cwl_40_66 word40_66 gnd C_wl
Rw41_66 word41_66 word40_66 R_wl
Cwl_41_66 word41_66 gnd C_wl
Rw42_66 word42_66 word41_66 R_wl
Cwl_42_66 word42_66 gnd C_wl
Rw43_66 word43_66 word42_66 R_wl
Cwl_43_66 word43_66 gnd C_wl
Rw44_66 word44_66 word43_66 R_wl
Cwl_44_66 word44_66 gnd C_wl
Rw45_66 word45_66 word44_66 R_wl
Cwl_45_66 word45_66 gnd C_wl
Rw46_66 word46_66 word45_66 R_wl
Cwl_46_66 word46_66 gnd C_wl
Rw47_66 word47_66 word46_66 R_wl
Cwl_47_66 word47_66 gnd C_wl
Rw48_66 word48_66 word47_66 R_wl
Cwl_48_66 word48_66 gnd C_wl
Rw49_66 word49_66 word48_66 R_wl
Cwl_49_66 word49_66 gnd C_wl
Rw50_66 word50_66 word49_66 R_wl
Cwl_50_66 word50_66 gnd C_wl
Rw51_66 word51_66 word50_66 R_wl
Cwl_51_66 word51_66 gnd C_wl
Rw52_66 word52_66 word51_66 R_wl
Cwl_52_66 word52_66 gnd C_wl
Rw53_66 word53_66 word52_66 R_wl
Cwl_53_66 word53_66 gnd C_wl
Rw54_66 word54_66 word53_66 R_wl
Cwl_54_66 word54_66 gnd C_wl
Rw55_66 word55_66 word54_66 R_wl
Cwl_55_66 word55_66 gnd C_wl
Rw56_66 word56_66 word55_66 R_wl
Cwl_56_66 word56_66 gnd C_wl
Rw57_66 word57_66 word56_66 R_wl
Cwl_57_66 word57_66 gnd C_wl
Rw58_66 word58_66 word57_66 R_wl
Cwl_58_66 word58_66 gnd C_wl
Rw59_66 word59_66 word58_66 R_wl
Cwl_59_66 word59_66 gnd C_wl
Rw60_66 word60_66 word59_66 R_wl
Cwl_60_66 word60_66 gnd C_wl
Rw61_66 word61_66 word60_66 R_wl
Cwl_61_66 word61_66 gnd C_wl
Rw62_66 word62_66 word61_66 R_wl
Cwl_62_66 word62_66 gnd C_wl
Rw63_66 word63_66 word62_66 R_wl
Cwl_63_66 word63_66 gnd C_wl
Rw64_66 word64_66 word63_66 R_wl
Cwl_64_66 word64_66 gnd C_wl
Rw65_66 word65_66 word64_66 R_wl
Cwl_65_66 word65_66 gnd C_wl
Rw66_66 word66_66 word65_66 R_wl
Cwl_66_66 word66_66 gnd C_wl
Rw67_66 word67_66 word66_66 R_wl
Cwl_67_66 word67_66 gnd C_wl
Rw68_66 word68_66 word67_66 R_wl
Cwl_68_66 word68_66 gnd C_wl
Rw69_66 word69_66 word68_66 R_wl
Cwl_69_66 word69_66 gnd C_wl
Rw70_66 word70_66 word69_66 R_wl
Cwl_70_66 word70_66 gnd C_wl
Rw71_66 word71_66 word70_66 R_wl
Cwl_71_66 word71_66 gnd C_wl
Rw72_66 word72_66 word71_66 R_wl
Cwl_72_66 word72_66 gnd C_wl
Rw73_66 word73_66 word72_66 R_wl
Cwl_73_66 word73_66 gnd C_wl
Rw74_66 word74_66 word73_66 R_wl
Cwl_74_66 word74_66 gnd C_wl
Rw75_66 word75_66 word74_66 R_wl
Cwl_75_66 word75_66 gnd C_wl
Rw76_66 word76_66 word75_66 R_wl
Cwl_76_66 word76_66 gnd C_wl
Rw77_66 word77_66 word76_66 R_wl
Cwl_77_66 word77_66 gnd C_wl
Rw78_66 word78_66 word77_66 R_wl
Cwl_78_66 word78_66 gnd C_wl
Rw79_66 word79_66 word78_66 R_wl
Cwl_79_66 word79_66 gnd C_wl
Rw80_66 word80_66 word79_66 R_wl
Cwl_80_66 word80_66 gnd C_wl
Rw81_66 word81_66 word80_66 R_wl
Cwl_81_66 word81_66 gnd C_wl
Rw82_66 word82_66 word81_66 R_wl
Cwl_82_66 word82_66 gnd C_wl
Rw83_66 word83_66 word82_66 R_wl
Cwl_83_66 word83_66 gnd C_wl
Rw84_66 word84_66 word83_66 R_wl
Cwl_84_66 word84_66 gnd C_wl
Rw85_66 word85_66 word84_66 R_wl
Cwl_85_66 word85_66 gnd C_wl
Rw86_66 word86_66 word85_66 R_wl
Cwl_86_66 word86_66 gnd C_wl
Rw87_66 word87_66 word86_66 R_wl
Cwl_87_66 word87_66 gnd C_wl
Rw88_66 word88_66 word87_66 R_wl
Cwl_88_66 word88_66 gnd C_wl
Rw89_66 word89_66 word88_66 R_wl
Cwl_89_66 word89_66 gnd C_wl
Rw90_66 word90_66 word89_66 R_wl
Cwl_90_66 word90_66 gnd C_wl
Rw91_66 word91_66 word90_66 R_wl
Cwl_91_66 word91_66 gnd C_wl
Rw92_66 word92_66 word91_66 R_wl
Cwl_92_66 word92_66 gnd C_wl
Rw93_66 word93_66 word92_66 R_wl
Cwl_93_66 word93_66 gnd C_wl
Rw94_66 word94_66 word93_66 R_wl
Cwl_94_66 word94_66 gnd C_wl
Rw95_66 word95_66 word94_66 R_wl
Cwl_95_66 word95_66 gnd C_wl
Rw96_66 word96_66 word95_66 R_wl
Cwl_96_66 word96_66 gnd C_wl
Rw97_66 word97_66 word96_66 R_wl
Cwl_97_66 word97_66 gnd C_wl
Rw98_66 word98_66 word97_66 R_wl
Cwl_98_66 word98_66 gnd C_wl
Rw99_66 word99_66 word98_66 R_wl
Cwl_99_66 word99_66 gnd C_wl
Vwl_67 word_67 0 0
Rw0_67 word_67 word0_67 R_wl
Cwl_0_67 word0_67 gnd C_wl
Rw1_67 word1_67 word0_67 R_wl
Cwl_1_67 word1_67 gnd C_wl
Rw2_67 word2_67 word1_67 R_wl
Cwl_2_67 word2_67 gnd C_wl
Rw3_67 word3_67 word2_67 R_wl
Cwl_3_67 word3_67 gnd C_wl
Rw4_67 word4_67 word3_67 R_wl
Cwl_4_67 word4_67 gnd C_wl
Rw5_67 word5_67 word4_67 R_wl
Cwl_5_67 word5_67 gnd C_wl
Rw6_67 word6_67 word5_67 R_wl
Cwl_6_67 word6_67 gnd C_wl
Rw7_67 word7_67 word6_67 R_wl
Cwl_7_67 word7_67 gnd C_wl
Rw8_67 word8_67 word7_67 R_wl
Cwl_8_67 word8_67 gnd C_wl
Rw9_67 word9_67 word8_67 R_wl
Cwl_9_67 word9_67 gnd C_wl
Rw10_67 word10_67 word9_67 R_wl
Cwl_10_67 word10_67 gnd C_wl
Rw11_67 word11_67 word10_67 R_wl
Cwl_11_67 word11_67 gnd C_wl
Rw12_67 word12_67 word11_67 R_wl
Cwl_12_67 word12_67 gnd C_wl
Rw13_67 word13_67 word12_67 R_wl
Cwl_13_67 word13_67 gnd C_wl
Rw14_67 word14_67 word13_67 R_wl
Cwl_14_67 word14_67 gnd C_wl
Rw15_67 word15_67 word14_67 R_wl
Cwl_15_67 word15_67 gnd C_wl
Rw16_67 word16_67 word15_67 R_wl
Cwl_16_67 word16_67 gnd C_wl
Rw17_67 word17_67 word16_67 R_wl
Cwl_17_67 word17_67 gnd C_wl
Rw18_67 word18_67 word17_67 R_wl
Cwl_18_67 word18_67 gnd C_wl
Rw19_67 word19_67 word18_67 R_wl
Cwl_19_67 word19_67 gnd C_wl
Rw20_67 word20_67 word19_67 R_wl
Cwl_20_67 word20_67 gnd C_wl
Rw21_67 word21_67 word20_67 R_wl
Cwl_21_67 word21_67 gnd C_wl
Rw22_67 word22_67 word21_67 R_wl
Cwl_22_67 word22_67 gnd C_wl
Rw23_67 word23_67 word22_67 R_wl
Cwl_23_67 word23_67 gnd C_wl
Rw24_67 word24_67 word23_67 R_wl
Cwl_24_67 word24_67 gnd C_wl
Rw25_67 word25_67 word24_67 R_wl
Cwl_25_67 word25_67 gnd C_wl
Rw26_67 word26_67 word25_67 R_wl
Cwl_26_67 word26_67 gnd C_wl
Rw27_67 word27_67 word26_67 R_wl
Cwl_27_67 word27_67 gnd C_wl
Rw28_67 word28_67 word27_67 R_wl
Cwl_28_67 word28_67 gnd C_wl
Rw29_67 word29_67 word28_67 R_wl
Cwl_29_67 word29_67 gnd C_wl
Rw30_67 word30_67 word29_67 R_wl
Cwl_30_67 word30_67 gnd C_wl
Rw31_67 word31_67 word30_67 R_wl
Cwl_31_67 word31_67 gnd C_wl
Rw32_67 word32_67 word31_67 R_wl
Cwl_32_67 word32_67 gnd C_wl
Rw33_67 word33_67 word32_67 R_wl
Cwl_33_67 word33_67 gnd C_wl
Rw34_67 word34_67 word33_67 R_wl
Cwl_34_67 word34_67 gnd C_wl
Rw35_67 word35_67 word34_67 R_wl
Cwl_35_67 word35_67 gnd C_wl
Rw36_67 word36_67 word35_67 R_wl
Cwl_36_67 word36_67 gnd C_wl
Rw37_67 word37_67 word36_67 R_wl
Cwl_37_67 word37_67 gnd C_wl
Rw38_67 word38_67 word37_67 R_wl
Cwl_38_67 word38_67 gnd C_wl
Rw39_67 word39_67 word38_67 R_wl
Cwl_39_67 word39_67 gnd C_wl
Rw40_67 word40_67 word39_67 R_wl
Cwl_40_67 word40_67 gnd C_wl
Rw41_67 word41_67 word40_67 R_wl
Cwl_41_67 word41_67 gnd C_wl
Rw42_67 word42_67 word41_67 R_wl
Cwl_42_67 word42_67 gnd C_wl
Rw43_67 word43_67 word42_67 R_wl
Cwl_43_67 word43_67 gnd C_wl
Rw44_67 word44_67 word43_67 R_wl
Cwl_44_67 word44_67 gnd C_wl
Rw45_67 word45_67 word44_67 R_wl
Cwl_45_67 word45_67 gnd C_wl
Rw46_67 word46_67 word45_67 R_wl
Cwl_46_67 word46_67 gnd C_wl
Rw47_67 word47_67 word46_67 R_wl
Cwl_47_67 word47_67 gnd C_wl
Rw48_67 word48_67 word47_67 R_wl
Cwl_48_67 word48_67 gnd C_wl
Rw49_67 word49_67 word48_67 R_wl
Cwl_49_67 word49_67 gnd C_wl
Rw50_67 word50_67 word49_67 R_wl
Cwl_50_67 word50_67 gnd C_wl
Rw51_67 word51_67 word50_67 R_wl
Cwl_51_67 word51_67 gnd C_wl
Rw52_67 word52_67 word51_67 R_wl
Cwl_52_67 word52_67 gnd C_wl
Rw53_67 word53_67 word52_67 R_wl
Cwl_53_67 word53_67 gnd C_wl
Rw54_67 word54_67 word53_67 R_wl
Cwl_54_67 word54_67 gnd C_wl
Rw55_67 word55_67 word54_67 R_wl
Cwl_55_67 word55_67 gnd C_wl
Rw56_67 word56_67 word55_67 R_wl
Cwl_56_67 word56_67 gnd C_wl
Rw57_67 word57_67 word56_67 R_wl
Cwl_57_67 word57_67 gnd C_wl
Rw58_67 word58_67 word57_67 R_wl
Cwl_58_67 word58_67 gnd C_wl
Rw59_67 word59_67 word58_67 R_wl
Cwl_59_67 word59_67 gnd C_wl
Rw60_67 word60_67 word59_67 R_wl
Cwl_60_67 word60_67 gnd C_wl
Rw61_67 word61_67 word60_67 R_wl
Cwl_61_67 word61_67 gnd C_wl
Rw62_67 word62_67 word61_67 R_wl
Cwl_62_67 word62_67 gnd C_wl
Rw63_67 word63_67 word62_67 R_wl
Cwl_63_67 word63_67 gnd C_wl
Rw64_67 word64_67 word63_67 R_wl
Cwl_64_67 word64_67 gnd C_wl
Rw65_67 word65_67 word64_67 R_wl
Cwl_65_67 word65_67 gnd C_wl
Rw66_67 word66_67 word65_67 R_wl
Cwl_66_67 word66_67 gnd C_wl
Rw67_67 word67_67 word66_67 R_wl
Cwl_67_67 word67_67 gnd C_wl
Rw68_67 word68_67 word67_67 R_wl
Cwl_68_67 word68_67 gnd C_wl
Rw69_67 word69_67 word68_67 R_wl
Cwl_69_67 word69_67 gnd C_wl
Rw70_67 word70_67 word69_67 R_wl
Cwl_70_67 word70_67 gnd C_wl
Rw71_67 word71_67 word70_67 R_wl
Cwl_71_67 word71_67 gnd C_wl
Rw72_67 word72_67 word71_67 R_wl
Cwl_72_67 word72_67 gnd C_wl
Rw73_67 word73_67 word72_67 R_wl
Cwl_73_67 word73_67 gnd C_wl
Rw74_67 word74_67 word73_67 R_wl
Cwl_74_67 word74_67 gnd C_wl
Rw75_67 word75_67 word74_67 R_wl
Cwl_75_67 word75_67 gnd C_wl
Rw76_67 word76_67 word75_67 R_wl
Cwl_76_67 word76_67 gnd C_wl
Rw77_67 word77_67 word76_67 R_wl
Cwl_77_67 word77_67 gnd C_wl
Rw78_67 word78_67 word77_67 R_wl
Cwl_78_67 word78_67 gnd C_wl
Rw79_67 word79_67 word78_67 R_wl
Cwl_79_67 word79_67 gnd C_wl
Rw80_67 word80_67 word79_67 R_wl
Cwl_80_67 word80_67 gnd C_wl
Rw81_67 word81_67 word80_67 R_wl
Cwl_81_67 word81_67 gnd C_wl
Rw82_67 word82_67 word81_67 R_wl
Cwl_82_67 word82_67 gnd C_wl
Rw83_67 word83_67 word82_67 R_wl
Cwl_83_67 word83_67 gnd C_wl
Rw84_67 word84_67 word83_67 R_wl
Cwl_84_67 word84_67 gnd C_wl
Rw85_67 word85_67 word84_67 R_wl
Cwl_85_67 word85_67 gnd C_wl
Rw86_67 word86_67 word85_67 R_wl
Cwl_86_67 word86_67 gnd C_wl
Rw87_67 word87_67 word86_67 R_wl
Cwl_87_67 word87_67 gnd C_wl
Rw88_67 word88_67 word87_67 R_wl
Cwl_88_67 word88_67 gnd C_wl
Rw89_67 word89_67 word88_67 R_wl
Cwl_89_67 word89_67 gnd C_wl
Rw90_67 word90_67 word89_67 R_wl
Cwl_90_67 word90_67 gnd C_wl
Rw91_67 word91_67 word90_67 R_wl
Cwl_91_67 word91_67 gnd C_wl
Rw92_67 word92_67 word91_67 R_wl
Cwl_92_67 word92_67 gnd C_wl
Rw93_67 word93_67 word92_67 R_wl
Cwl_93_67 word93_67 gnd C_wl
Rw94_67 word94_67 word93_67 R_wl
Cwl_94_67 word94_67 gnd C_wl
Rw95_67 word95_67 word94_67 R_wl
Cwl_95_67 word95_67 gnd C_wl
Rw96_67 word96_67 word95_67 R_wl
Cwl_96_67 word96_67 gnd C_wl
Rw97_67 word97_67 word96_67 R_wl
Cwl_97_67 word97_67 gnd C_wl
Rw98_67 word98_67 word97_67 R_wl
Cwl_98_67 word98_67 gnd C_wl
Rw99_67 word99_67 word98_67 R_wl
Cwl_99_67 word99_67 gnd C_wl
Vwl_68 word_68 0 0
Rw0_68 word_68 word0_68 R_wl
Cwl_0_68 word0_68 gnd C_wl
Rw1_68 word1_68 word0_68 R_wl
Cwl_1_68 word1_68 gnd C_wl
Rw2_68 word2_68 word1_68 R_wl
Cwl_2_68 word2_68 gnd C_wl
Rw3_68 word3_68 word2_68 R_wl
Cwl_3_68 word3_68 gnd C_wl
Rw4_68 word4_68 word3_68 R_wl
Cwl_4_68 word4_68 gnd C_wl
Rw5_68 word5_68 word4_68 R_wl
Cwl_5_68 word5_68 gnd C_wl
Rw6_68 word6_68 word5_68 R_wl
Cwl_6_68 word6_68 gnd C_wl
Rw7_68 word7_68 word6_68 R_wl
Cwl_7_68 word7_68 gnd C_wl
Rw8_68 word8_68 word7_68 R_wl
Cwl_8_68 word8_68 gnd C_wl
Rw9_68 word9_68 word8_68 R_wl
Cwl_9_68 word9_68 gnd C_wl
Rw10_68 word10_68 word9_68 R_wl
Cwl_10_68 word10_68 gnd C_wl
Rw11_68 word11_68 word10_68 R_wl
Cwl_11_68 word11_68 gnd C_wl
Rw12_68 word12_68 word11_68 R_wl
Cwl_12_68 word12_68 gnd C_wl
Rw13_68 word13_68 word12_68 R_wl
Cwl_13_68 word13_68 gnd C_wl
Rw14_68 word14_68 word13_68 R_wl
Cwl_14_68 word14_68 gnd C_wl
Rw15_68 word15_68 word14_68 R_wl
Cwl_15_68 word15_68 gnd C_wl
Rw16_68 word16_68 word15_68 R_wl
Cwl_16_68 word16_68 gnd C_wl
Rw17_68 word17_68 word16_68 R_wl
Cwl_17_68 word17_68 gnd C_wl
Rw18_68 word18_68 word17_68 R_wl
Cwl_18_68 word18_68 gnd C_wl
Rw19_68 word19_68 word18_68 R_wl
Cwl_19_68 word19_68 gnd C_wl
Rw20_68 word20_68 word19_68 R_wl
Cwl_20_68 word20_68 gnd C_wl
Rw21_68 word21_68 word20_68 R_wl
Cwl_21_68 word21_68 gnd C_wl
Rw22_68 word22_68 word21_68 R_wl
Cwl_22_68 word22_68 gnd C_wl
Rw23_68 word23_68 word22_68 R_wl
Cwl_23_68 word23_68 gnd C_wl
Rw24_68 word24_68 word23_68 R_wl
Cwl_24_68 word24_68 gnd C_wl
Rw25_68 word25_68 word24_68 R_wl
Cwl_25_68 word25_68 gnd C_wl
Rw26_68 word26_68 word25_68 R_wl
Cwl_26_68 word26_68 gnd C_wl
Rw27_68 word27_68 word26_68 R_wl
Cwl_27_68 word27_68 gnd C_wl
Rw28_68 word28_68 word27_68 R_wl
Cwl_28_68 word28_68 gnd C_wl
Rw29_68 word29_68 word28_68 R_wl
Cwl_29_68 word29_68 gnd C_wl
Rw30_68 word30_68 word29_68 R_wl
Cwl_30_68 word30_68 gnd C_wl
Rw31_68 word31_68 word30_68 R_wl
Cwl_31_68 word31_68 gnd C_wl
Rw32_68 word32_68 word31_68 R_wl
Cwl_32_68 word32_68 gnd C_wl
Rw33_68 word33_68 word32_68 R_wl
Cwl_33_68 word33_68 gnd C_wl
Rw34_68 word34_68 word33_68 R_wl
Cwl_34_68 word34_68 gnd C_wl
Rw35_68 word35_68 word34_68 R_wl
Cwl_35_68 word35_68 gnd C_wl
Rw36_68 word36_68 word35_68 R_wl
Cwl_36_68 word36_68 gnd C_wl
Rw37_68 word37_68 word36_68 R_wl
Cwl_37_68 word37_68 gnd C_wl
Rw38_68 word38_68 word37_68 R_wl
Cwl_38_68 word38_68 gnd C_wl
Rw39_68 word39_68 word38_68 R_wl
Cwl_39_68 word39_68 gnd C_wl
Rw40_68 word40_68 word39_68 R_wl
Cwl_40_68 word40_68 gnd C_wl
Rw41_68 word41_68 word40_68 R_wl
Cwl_41_68 word41_68 gnd C_wl
Rw42_68 word42_68 word41_68 R_wl
Cwl_42_68 word42_68 gnd C_wl
Rw43_68 word43_68 word42_68 R_wl
Cwl_43_68 word43_68 gnd C_wl
Rw44_68 word44_68 word43_68 R_wl
Cwl_44_68 word44_68 gnd C_wl
Rw45_68 word45_68 word44_68 R_wl
Cwl_45_68 word45_68 gnd C_wl
Rw46_68 word46_68 word45_68 R_wl
Cwl_46_68 word46_68 gnd C_wl
Rw47_68 word47_68 word46_68 R_wl
Cwl_47_68 word47_68 gnd C_wl
Rw48_68 word48_68 word47_68 R_wl
Cwl_48_68 word48_68 gnd C_wl
Rw49_68 word49_68 word48_68 R_wl
Cwl_49_68 word49_68 gnd C_wl
Rw50_68 word50_68 word49_68 R_wl
Cwl_50_68 word50_68 gnd C_wl
Rw51_68 word51_68 word50_68 R_wl
Cwl_51_68 word51_68 gnd C_wl
Rw52_68 word52_68 word51_68 R_wl
Cwl_52_68 word52_68 gnd C_wl
Rw53_68 word53_68 word52_68 R_wl
Cwl_53_68 word53_68 gnd C_wl
Rw54_68 word54_68 word53_68 R_wl
Cwl_54_68 word54_68 gnd C_wl
Rw55_68 word55_68 word54_68 R_wl
Cwl_55_68 word55_68 gnd C_wl
Rw56_68 word56_68 word55_68 R_wl
Cwl_56_68 word56_68 gnd C_wl
Rw57_68 word57_68 word56_68 R_wl
Cwl_57_68 word57_68 gnd C_wl
Rw58_68 word58_68 word57_68 R_wl
Cwl_58_68 word58_68 gnd C_wl
Rw59_68 word59_68 word58_68 R_wl
Cwl_59_68 word59_68 gnd C_wl
Rw60_68 word60_68 word59_68 R_wl
Cwl_60_68 word60_68 gnd C_wl
Rw61_68 word61_68 word60_68 R_wl
Cwl_61_68 word61_68 gnd C_wl
Rw62_68 word62_68 word61_68 R_wl
Cwl_62_68 word62_68 gnd C_wl
Rw63_68 word63_68 word62_68 R_wl
Cwl_63_68 word63_68 gnd C_wl
Rw64_68 word64_68 word63_68 R_wl
Cwl_64_68 word64_68 gnd C_wl
Rw65_68 word65_68 word64_68 R_wl
Cwl_65_68 word65_68 gnd C_wl
Rw66_68 word66_68 word65_68 R_wl
Cwl_66_68 word66_68 gnd C_wl
Rw67_68 word67_68 word66_68 R_wl
Cwl_67_68 word67_68 gnd C_wl
Rw68_68 word68_68 word67_68 R_wl
Cwl_68_68 word68_68 gnd C_wl
Rw69_68 word69_68 word68_68 R_wl
Cwl_69_68 word69_68 gnd C_wl
Rw70_68 word70_68 word69_68 R_wl
Cwl_70_68 word70_68 gnd C_wl
Rw71_68 word71_68 word70_68 R_wl
Cwl_71_68 word71_68 gnd C_wl
Rw72_68 word72_68 word71_68 R_wl
Cwl_72_68 word72_68 gnd C_wl
Rw73_68 word73_68 word72_68 R_wl
Cwl_73_68 word73_68 gnd C_wl
Rw74_68 word74_68 word73_68 R_wl
Cwl_74_68 word74_68 gnd C_wl
Rw75_68 word75_68 word74_68 R_wl
Cwl_75_68 word75_68 gnd C_wl
Rw76_68 word76_68 word75_68 R_wl
Cwl_76_68 word76_68 gnd C_wl
Rw77_68 word77_68 word76_68 R_wl
Cwl_77_68 word77_68 gnd C_wl
Rw78_68 word78_68 word77_68 R_wl
Cwl_78_68 word78_68 gnd C_wl
Rw79_68 word79_68 word78_68 R_wl
Cwl_79_68 word79_68 gnd C_wl
Rw80_68 word80_68 word79_68 R_wl
Cwl_80_68 word80_68 gnd C_wl
Rw81_68 word81_68 word80_68 R_wl
Cwl_81_68 word81_68 gnd C_wl
Rw82_68 word82_68 word81_68 R_wl
Cwl_82_68 word82_68 gnd C_wl
Rw83_68 word83_68 word82_68 R_wl
Cwl_83_68 word83_68 gnd C_wl
Rw84_68 word84_68 word83_68 R_wl
Cwl_84_68 word84_68 gnd C_wl
Rw85_68 word85_68 word84_68 R_wl
Cwl_85_68 word85_68 gnd C_wl
Rw86_68 word86_68 word85_68 R_wl
Cwl_86_68 word86_68 gnd C_wl
Rw87_68 word87_68 word86_68 R_wl
Cwl_87_68 word87_68 gnd C_wl
Rw88_68 word88_68 word87_68 R_wl
Cwl_88_68 word88_68 gnd C_wl
Rw89_68 word89_68 word88_68 R_wl
Cwl_89_68 word89_68 gnd C_wl
Rw90_68 word90_68 word89_68 R_wl
Cwl_90_68 word90_68 gnd C_wl
Rw91_68 word91_68 word90_68 R_wl
Cwl_91_68 word91_68 gnd C_wl
Rw92_68 word92_68 word91_68 R_wl
Cwl_92_68 word92_68 gnd C_wl
Rw93_68 word93_68 word92_68 R_wl
Cwl_93_68 word93_68 gnd C_wl
Rw94_68 word94_68 word93_68 R_wl
Cwl_94_68 word94_68 gnd C_wl
Rw95_68 word95_68 word94_68 R_wl
Cwl_95_68 word95_68 gnd C_wl
Rw96_68 word96_68 word95_68 R_wl
Cwl_96_68 word96_68 gnd C_wl
Rw97_68 word97_68 word96_68 R_wl
Cwl_97_68 word97_68 gnd C_wl
Rw98_68 word98_68 word97_68 R_wl
Cwl_98_68 word98_68 gnd C_wl
Rw99_68 word99_68 word98_68 R_wl
Cwl_99_68 word99_68 gnd C_wl
Vwl_69 word_69 0 0
Rw0_69 word_69 word0_69 R_wl
Cwl_0_69 word0_69 gnd C_wl
Rw1_69 word1_69 word0_69 R_wl
Cwl_1_69 word1_69 gnd C_wl
Rw2_69 word2_69 word1_69 R_wl
Cwl_2_69 word2_69 gnd C_wl
Rw3_69 word3_69 word2_69 R_wl
Cwl_3_69 word3_69 gnd C_wl
Rw4_69 word4_69 word3_69 R_wl
Cwl_4_69 word4_69 gnd C_wl
Rw5_69 word5_69 word4_69 R_wl
Cwl_5_69 word5_69 gnd C_wl
Rw6_69 word6_69 word5_69 R_wl
Cwl_6_69 word6_69 gnd C_wl
Rw7_69 word7_69 word6_69 R_wl
Cwl_7_69 word7_69 gnd C_wl
Rw8_69 word8_69 word7_69 R_wl
Cwl_8_69 word8_69 gnd C_wl
Rw9_69 word9_69 word8_69 R_wl
Cwl_9_69 word9_69 gnd C_wl
Rw10_69 word10_69 word9_69 R_wl
Cwl_10_69 word10_69 gnd C_wl
Rw11_69 word11_69 word10_69 R_wl
Cwl_11_69 word11_69 gnd C_wl
Rw12_69 word12_69 word11_69 R_wl
Cwl_12_69 word12_69 gnd C_wl
Rw13_69 word13_69 word12_69 R_wl
Cwl_13_69 word13_69 gnd C_wl
Rw14_69 word14_69 word13_69 R_wl
Cwl_14_69 word14_69 gnd C_wl
Rw15_69 word15_69 word14_69 R_wl
Cwl_15_69 word15_69 gnd C_wl
Rw16_69 word16_69 word15_69 R_wl
Cwl_16_69 word16_69 gnd C_wl
Rw17_69 word17_69 word16_69 R_wl
Cwl_17_69 word17_69 gnd C_wl
Rw18_69 word18_69 word17_69 R_wl
Cwl_18_69 word18_69 gnd C_wl
Rw19_69 word19_69 word18_69 R_wl
Cwl_19_69 word19_69 gnd C_wl
Rw20_69 word20_69 word19_69 R_wl
Cwl_20_69 word20_69 gnd C_wl
Rw21_69 word21_69 word20_69 R_wl
Cwl_21_69 word21_69 gnd C_wl
Rw22_69 word22_69 word21_69 R_wl
Cwl_22_69 word22_69 gnd C_wl
Rw23_69 word23_69 word22_69 R_wl
Cwl_23_69 word23_69 gnd C_wl
Rw24_69 word24_69 word23_69 R_wl
Cwl_24_69 word24_69 gnd C_wl
Rw25_69 word25_69 word24_69 R_wl
Cwl_25_69 word25_69 gnd C_wl
Rw26_69 word26_69 word25_69 R_wl
Cwl_26_69 word26_69 gnd C_wl
Rw27_69 word27_69 word26_69 R_wl
Cwl_27_69 word27_69 gnd C_wl
Rw28_69 word28_69 word27_69 R_wl
Cwl_28_69 word28_69 gnd C_wl
Rw29_69 word29_69 word28_69 R_wl
Cwl_29_69 word29_69 gnd C_wl
Rw30_69 word30_69 word29_69 R_wl
Cwl_30_69 word30_69 gnd C_wl
Rw31_69 word31_69 word30_69 R_wl
Cwl_31_69 word31_69 gnd C_wl
Rw32_69 word32_69 word31_69 R_wl
Cwl_32_69 word32_69 gnd C_wl
Rw33_69 word33_69 word32_69 R_wl
Cwl_33_69 word33_69 gnd C_wl
Rw34_69 word34_69 word33_69 R_wl
Cwl_34_69 word34_69 gnd C_wl
Rw35_69 word35_69 word34_69 R_wl
Cwl_35_69 word35_69 gnd C_wl
Rw36_69 word36_69 word35_69 R_wl
Cwl_36_69 word36_69 gnd C_wl
Rw37_69 word37_69 word36_69 R_wl
Cwl_37_69 word37_69 gnd C_wl
Rw38_69 word38_69 word37_69 R_wl
Cwl_38_69 word38_69 gnd C_wl
Rw39_69 word39_69 word38_69 R_wl
Cwl_39_69 word39_69 gnd C_wl
Rw40_69 word40_69 word39_69 R_wl
Cwl_40_69 word40_69 gnd C_wl
Rw41_69 word41_69 word40_69 R_wl
Cwl_41_69 word41_69 gnd C_wl
Rw42_69 word42_69 word41_69 R_wl
Cwl_42_69 word42_69 gnd C_wl
Rw43_69 word43_69 word42_69 R_wl
Cwl_43_69 word43_69 gnd C_wl
Rw44_69 word44_69 word43_69 R_wl
Cwl_44_69 word44_69 gnd C_wl
Rw45_69 word45_69 word44_69 R_wl
Cwl_45_69 word45_69 gnd C_wl
Rw46_69 word46_69 word45_69 R_wl
Cwl_46_69 word46_69 gnd C_wl
Rw47_69 word47_69 word46_69 R_wl
Cwl_47_69 word47_69 gnd C_wl
Rw48_69 word48_69 word47_69 R_wl
Cwl_48_69 word48_69 gnd C_wl
Rw49_69 word49_69 word48_69 R_wl
Cwl_49_69 word49_69 gnd C_wl
Rw50_69 word50_69 word49_69 R_wl
Cwl_50_69 word50_69 gnd C_wl
Rw51_69 word51_69 word50_69 R_wl
Cwl_51_69 word51_69 gnd C_wl
Rw52_69 word52_69 word51_69 R_wl
Cwl_52_69 word52_69 gnd C_wl
Rw53_69 word53_69 word52_69 R_wl
Cwl_53_69 word53_69 gnd C_wl
Rw54_69 word54_69 word53_69 R_wl
Cwl_54_69 word54_69 gnd C_wl
Rw55_69 word55_69 word54_69 R_wl
Cwl_55_69 word55_69 gnd C_wl
Rw56_69 word56_69 word55_69 R_wl
Cwl_56_69 word56_69 gnd C_wl
Rw57_69 word57_69 word56_69 R_wl
Cwl_57_69 word57_69 gnd C_wl
Rw58_69 word58_69 word57_69 R_wl
Cwl_58_69 word58_69 gnd C_wl
Rw59_69 word59_69 word58_69 R_wl
Cwl_59_69 word59_69 gnd C_wl
Rw60_69 word60_69 word59_69 R_wl
Cwl_60_69 word60_69 gnd C_wl
Rw61_69 word61_69 word60_69 R_wl
Cwl_61_69 word61_69 gnd C_wl
Rw62_69 word62_69 word61_69 R_wl
Cwl_62_69 word62_69 gnd C_wl
Rw63_69 word63_69 word62_69 R_wl
Cwl_63_69 word63_69 gnd C_wl
Rw64_69 word64_69 word63_69 R_wl
Cwl_64_69 word64_69 gnd C_wl
Rw65_69 word65_69 word64_69 R_wl
Cwl_65_69 word65_69 gnd C_wl
Rw66_69 word66_69 word65_69 R_wl
Cwl_66_69 word66_69 gnd C_wl
Rw67_69 word67_69 word66_69 R_wl
Cwl_67_69 word67_69 gnd C_wl
Rw68_69 word68_69 word67_69 R_wl
Cwl_68_69 word68_69 gnd C_wl
Rw69_69 word69_69 word68_69 R_wl
Cwl_69_69 word69_69 gnd C_wl
Rw70_69 word70_69 word69_69 R_wl
Cwl_70_69 word70_69 gnd C_wl
Rw71_69 word71_69 word70_69 R_wl
Cwl_71_69 word71_69 gnd C_wl
Rw72_69 word72_69 word71_69 R_wl
Cwl_72_69 word72_69 gnd C_wl
Rw73_69 word73_69 word72_69 R_wl
Cwl_73_69 word73_69 gnd C_wl
Rw74_69 word74_69 word73_69 R_wl
Cwl_74_69 word74_69 gnd C_wl
Rw75_69 word75_69 word74_69 R_wl
Cwl_75_69 word75_69 gnd C_wl
Rw76_69 word76_69 word75_69 R_wl
Cwl_76_69 word76_69 gnd C_wl
Rw77_69 word77_69 word76_69 R_wl
Cwl_77_69 word77_69 gnd C_wl
Rw78_69 word78_69 word77_69 R_wl
Cwl_78_69 word78_69 gnd C_wl
Rw79_69 word79_69 word78_69 R_wl
Cwl_79_69 word79_69 gnd C_wl
Rw80_69 word80_69 word79_69 R_wl
Cwl_80_69 word80_69 gnd C_wl
Rw81_69 word81_69 word80_69 R_wl
Cwl_81_69 word81_69 gnd C_wl
Rw82_69 word82_69 word81_69 R_wl
Cwl_82_69 word82_69 gnd C_wl
Rw83_69 word83_69 word82_69 R_wl
Cwl_83_69 word83_69 gnd C_wl
Rw84_69 word84_69 word83_69 R_wl
Cwl_84_69 word84_69 gnd C_wl
Rw85_69 word85_69 word84_69 R_wl
Cwl_85_69 word85_69 gnd C_wl
Rw86_69 word86_69 word85_69 R_wl
Cwl_86_69 word86_69 gnd C_wl
Rw87_69 word87_69 word86_69 R_wl
Cwl_87_69 word87_69 gnd C_wl
Rw88_69 word88_69 word87_69 R_wl
Cwl_88_69 word88_69 gnd C_wl
Rw89_69 word89_69 word88_69 R_wl
Cwl_89_69 word89_69 gnd C_wl
Rw90_69 word90_69 word89_69 R_wl
Cwl_90_69 word90_69 gnd C_wl
Rw91_69 word91_69 word90_69 R_wl
Cwl_91_69 word91_69 gnd C_wl
Rw92_69 word92_69 word91_69 R_wl
Cwl_92_69 word92_69 gnd C_wl
Rw93_69 word93_69 word92_69 R_wl
Cwl_93_69 word93_69 gnd C_wl
Rw94_69 word94_69 word93_69 R_wl
Cwl_94_69 word94_69 gnd C_wl
Rw95_69 word95_69 word94_69 R_wl
Cwl_95_69 word95_69 gnd C_wl
Rw96_69 word96_69 word95_69 R_wl
Cwl_96_69 word96_69 gnd C_wl
Rw97_69 word97_69 word96_69 R_wl
Cwl_97_69 word97_69 gnd C_wl
Rw98_69 word98_69 word97_69 R_wl
Cwl_98_69 word98_69 gnd C_wl
Rw99_69 word99_69 word98_69 R_wl
Cwl_99_69 word99_69 gnd C_wl
Vwl_70 word_70 0 0
Rw0_70 word_70 word0_70 R_wl
Cwl_0_70 word0_70 gnd C_wl
Rw1_70 word1_70 word0_70 R_wl
Cwl_1_70 word1_70 gnd C_wl
Rw2_70 word2_70 word1_70 R_wl
Cwl_2_70 word2_70 gnd C_wl
Rw3_70 word3_70 word2_70 R_wl
Cwl_3_70 word3_70 gnd C_wl
Rw4_70 word4_70 word3_70 R_wl
Cwl_4_70 word4_70 gnd C_wl
Rw5_70 word5_70 word4_70 R_wl
Cwl_5_70 word5_70 gnd C_wl
Rw6_70 word6_70 word5_70 R_wl
Cwl_6_70 word6_70 gnd C_wl
Rw7_70 word7_70 word6_70 R_wl
Cwl_7_70 word7_70 gnd C_wl
Rw8_70 word8_70 word7_70 R_wl
Cwl_8_70 word8_70 gnd C_wl
Rw9_70 word9_70 word8_70 R_wl
Cwl_9_70 word9_70 gnd C_wl
Rw10_70 word10_70 word9_70 R_wl
Cwl_10_70 word10_70 gnd C_wl
Rw11_70 word11_70 word10_70 R_wl
Cwl_11_70 word11_70 gnd C_wl
Rw12_70 word12_70 word11_70 R_wl
Cwl_12_70 word12_70 gnd C_wl
Rw13_70 word13_70 word12_70 R_wl
Cwl_13_70 word13_70 gnd C_wl
Rw14_70 word14_70 word13_70 R_wl
Cwl_14_70 word14_70 gnd C_wl
Rw15_70 word15_70 word14_70 R_wl
Cwl_15_70 word15_70 gnd C_wl
Rw16_70 word16_70 word15_70 R_wl
Cwl_16_70 word16_70 gnd C_wl
Rw17_70 word17_70 word16_70 R_wl
Cwl_17_70 word17_70 gnd C_wl
Rw18_70 word18_70 word17_70 R_wl
Cwl_18_70 word18_70 gnd C_wl
Rw19_70 word19_70 word18_70 R_wl
Cwl_19_70 word19_70 gnd C_wl
Rw20_70 word20_70 word19_70 R_wl
Cwl_20_70 word20_70 gnd C_wl
Rw21_70 word21_70 word20_70 R_wl
Cwl_21_70 word21_70 gnd C_wl
Rw22_70 word22_70 word21_70 R_wl
Cwl_22_70 word22_70 gnd C_wl
Rw23_70 word23_70 word22_70 R_wl
Cwl_23_70 word23_70 gnd C_wl
Rw24_70 word24_70 word23_70 R_wl
Cwl_24_70 word24_70 gnd C_wl
Rw25_70 word25_70 word24_70 R_wl
Cwl_25_70 word25_70 gnd C_wl
Rw26_70 word26_70 word25_70 R_wl
Cwl_26_70 word26_70 gnd C_wl
Rw27_70 word27_70 word26_70 R_wl
Cwl_27_70 word27_70 gnd C_wl
Rw28_70 word28_70 word27_70 R_wl
Cwl_28_70 word28_70 gnd C_wl
Rw29_70 word29_70 word28_70 R_wl
Cwl_29_70 word29_70 gnd C_wl
Rw30_70 word30_70 word29_70 R_wl
Cwl_30_70 word30_70 gnd C_wl
Rw31_70 word31_70 word30_70 R_wl
Cwl_31_70 word31_70 gnd C_wl
Rw32_70 word32_70 word31_70 R_wl
Cwl_32_70 word32_70 gnd C_wl
Rw33_70 word33_70 word32_70 R_wl
Cwl_33_70 word33_70 gnd C_wl
Rw34_70 word34_70 word33_70 R_wl
Cwl_34_70 word34_70 gnd C_wl
Rw35_70 word35_70 word34_70 R_wl
Cwl_35_70 word35_70 gnd C_wl
Rw36_70 word36_70 word35_70 R_wl
Cwl_36_70 word36_70 gnd C_wl
Rw37_70 word37_70 word36_70 R_wl
Cwl_37_70 word37_70 gnd C_wl
Rw38_70 word38_70 word37_70 R_wl
Cwl_38_70 word38_70 gnd C_wl
Rw39_70 word39_70 word38_70 R_wl
Cwl_39_70 word39_70 gnd C_wl
Rw40_70 word40_70 word39_70 R_wl
Cwl_40_70 word40_70 gnd C_wl
Rw41_70 word41_70 word40_70 R_wl
Cwl_41_70 word41_70 gnd C_wl
Rw42_70 word42_70 word41_70 R_wl
Cwl_42_70 word42_70 gnd C_wl
Rw43_70 word43_70 word42_70 R_wl
Cwl_43_70 word43_70 gnd C_wl
Rw44_70 word44_70 word43_70 R_wl
Cwl_44_70 word44_70 gnd C_wl
Rw45_70 word45_70 word44_70 R_wl
Cwl_45_70 word45_70 gnd C_wl
Rw46_70 word46_70 word45_70 R_wl
Cwl_46_70 word46_70 gnd C_wl
Rw47_70 word47_70 word46_70 R_wl
Cwl_47_70 word47_70 gnd C_wl
Rw48_70 word48_70 word47_70 R_wl
Cwl_48_70 word48_70 gnd C_wl
Rw49_70 word49_70 word48_70 R_wl
Cwl_49_70 word49_70 gnd C_wl
Rw50_70 word50_70 word49_70 R_wl
Cwl_50_70 word50_70 gnd C_wl
Rw51_70 word51_70 word50_70 R_wl
Cwl_51_70 word51_70 gnd C_wl
Rw52_70 word52_70 word51_70 R_wl
Cwl_52_70 word52_70 gnd C_wl
Rw53_70 word53_70 word52_70 R_wl
Cwl_53_70 word53_70 gnd C_wl
Rw54_70 word54_70 word53_70 R_wl
Cwl_54_70 word54_70 gnd C_wl
Rw55_70 word55_70 word54_70 R_wl
Cwl_55_70 word55_70 gnd C_wl
Rw56_70 word56_70 word55_70 R_wl
Cwl_56_70 word56_70 gnd C_wl
Rw57_70 word57_70 word56_70 R_wl
Cwl_57_70 word57_70 gnd C_wl
Rw58_70 word58_70 word57_70 R_wl
Cwl_58_70 word58_70 gnd C_wl
Rw59_70 word59_70 word58_70 R_wl
Cwl_59_70 word59_70 gnd C_wl
Rw60_70 word60_70 word59_70 R_wl
Cwl_60_70 word60_70 gnd C_wl
Rw61_70 word61_70 word60_70 R_wl
Cwl_61_70 word61_70 gnd C_wl
Rw62_70 word62_70 word61_70 R_wl
Cwl_62_70 word62_70 gnd C_wl
Rw63_70 word63_70 word62_70 R_wl
Cwl_63_70 word63_70 gnd C_wl
Rw64_70 word64_70 word63_70 R_wl
Cwl_64_70 word64_70 gnd C_wl
Rw65_70 word65_70 word64_70 R_wl
Cwl_65_70 word65_70 gnd C_wl
Rw66_70 word66_70 word65_70 R_wl
Cwl_66_70 word66_70 gnd C_wl
Rw67_70 word67_70 word66_70 R_wl
Cwl_67_70 word67_70 gnd C_wl
Rw68_70 word68_70 word67_70 R_wl
Cwl_68_70 word68_70 gnd C_wl
Rw69_70 word69_70 word68_70 R_wl
Cwl_69_70 word69_70 gnd C_wl
Rw70_70 word70_70 word69_70 R_wl
Cwl_70_70 word70_70 gnd C_wl
Rw71_70 word71_70 word70_70 R_wl
Cwl_71_70 word71_70 gnd C_wl
Rw72_70 word72_70 word71_70 R_wl
Cwl_72_70 word72_70 gnd C_wl
Rw73_70 word73_70 word72_70 R_wl
Cwl_73_70 word73_70 gnd C_wl
Rw74_70 word74_70 word73_70 R_wl
Cwl_74_70 word74_70 gnd C_wl
Rw75_70 word75_70 word74_70 R_wl
Cwl_75_70 word75_70 gnd C_wl
Rw76_70 word76_70 word75_70 R_wl
Cwl_76_70 word76_70 gnd C_wl
Rw77_70 word77_70 word76_70 R_wl
Cwl_77_70 word77_70 gnd C_wl
Rw78_70 word78_70 word77_70 R_wl
Cwl_78_70 word78_70 gnd C_wl
Rw79_70 word79_70 word78_70 R_wl
Cwl_79_70 word79_70 gnd C_wl
Rw80_70 word80_70 word79_70 R_wl
Cwl_80_70 word80_70 gnd C_wl
Rw81_70 word81_70 word80_70 R_wl
Cwl_81_70 word81_70 gnd C_wl
Rw82_70 word82_70 word81_70 R_wl
Cwl_82_70 word82_70 gnd C_wl
Rw83_70 word83_70 word82_70 R_wl
Cwl_83_70 word83_70 gnd C_wl
Rw84_70 word84_70 word83_70 R_wl
Cwl_84_70 word84_70 gnd C_wl
Rw85_70 word85_70 word84_70 R_wl
Cwl_85_70 word85_70 gnd C_wl
Rw86_70 word86_70 word85_70 R_wl
Cwl_86_70 word86_70 gnd C_wl
Rw87_70 word87_70 word86_70 R_wl
Cwl_87_70 word87_70 gnd C_wl
Rw88_70 word88_70 word87_70 R_wl
Cwl_88_70 word88_70 gnd C_wl
Rw89_70 word89_70 word88_70 R_wl
Cwl_89_70 word89_70 gnd C_wl
Rw90_70 word90_70 word89_70 R_wl
Cwl_90_70 word90_70 gnd C_wl
Rw91_70 word91_70 word90_70 R_wl
Cwl_91_70 word91_70 gnd C_wl
Rw92_70 word92_70 word91_70 R_wl
Cwl_92_70 word92_70 gnd C_wl
Rw93_70 word93_70 word92_70 R_wl
Cwl_93_70 word93_70 gnd C_wl
Rw94_70 word94_70 word93_70 R_wl
Cwl_94_70 word94_70 gnd C_wl
Rw95_70 word95_70 word94_70 R_wl
Cwl_95_70 word95_70 gnd C_wl
Rw96_70 word96_70 word95_70 R_wl
Cwl_96_70 word96_70 gnd C_wl
Rw97_70 word97_70 word96_70 R_wl
Cwl_97_70 word97_70 gnd C_wl
Rw98_70 word98_70 word97_70 R_wl
Cwl_98_70 word98_70 gnd C_wl
Rw99_70 word99_70 word98_70 R_wl
Cwl_99_70 word99_70 gnd C_wl
Vwl_71 word_71 0 0
Rw0_71 word_71 word0_71 R_wl
Cwl_0_71 word0_71 gnd C_wl
Rw1_71 word1_71 word0_71 R_wl
Cwl_1_71 word1_71 gnd C_wl
Rw2_71 word2_71 word1_71 R_wl
Cwl_2_71 word2_71 gnd C_wl
Rw3_71 word3_71 word2_71 R_wl
Cwl_3_71 word3_71 gnd C_wl
Rw4_71 word4_71 word3_71 R_wl
Cwl_4_71 word4_71 gnd C_wl
Rw5_71 word5_71 word4_71 R_wl
Cwl_5_71 word5_71 gnd C_wl
Rw6_71 word6_71 word5_71 R_wl
Cwl_6_71 word6_71 gnd C_wl
Rw7_71 word7_71 word6_71 R_wl
Cwl_7_71 word7_71 gnd C_wl
Rw8_71 word8_71 word7_71 R_wl
Cwl_8_71 word8_71 gnd C_wl
Rw9_71 word9_71 word8_71 R_wl
Cwl_9_71 word9_71 gnd C_wl
Rw10_71 word10_71 word9_71 R_wl
Cwl_10_71 word10_71 gnd C_wl
Rw11_71 word11_71 word10_71 R_wl
Cwl_11_71 word11_71 gnd C_wl
Rw12_71 word12_71 word11_71 R_wl
Cwl_12_71 word12_71 gnd C_wl
Rw13_71 word13_71 word12_71 R_wl
Cwl_13_71 word13_71 gnd C_wl
Rw14_71 word14_71 word13_71 R_wl
Cwl_14_71 word14_71 gnd C_wl
Rw15_71 word15_71 word14_71 R_wl
Cwl_15_71 word15_71 gnd C_wl
Rw16_71 word16_71 word15_71 R_wl
Cwl_16_71 word16_71 gnd C_wl
Rw17_71 word17_71 word16_71 R_wl
Cwl_17_71 word17_71 gnd C_wl
Rw18_71 word18_71 word17_71 R_wl
Cwl_18_71 word18_71 gnd C_wl
Rw19_71 word19_71 word18_71 R_wl
Cwl_19_71 word19_71 gnd C_wl
Rw20_71 word20_71 word19_71 R_wl
Cwl_20_71 word20_71 gnd C_wl
Rw21_71 word21_71 word20_71 R_wl
Cwl_21_71 word21_71 gnd C_wl
Rw22_71 word22_71 word21_71 R_wl
Cwl_22_71 word22_71 gnd C_wl
Rw23_71 word23_71 word22_71 R_wl
Cwl_23_71 word23_71 gnd C_wl
Rw24_71 word24_71 word23_71 R_wl
Cwl_24_71 word24_71 gnd C_wl
Rw25_71 word25_71 word24_71 R_wl
Cwl_25_71 word25_71 gnd C_wl
Rw26_71 word26_71 word25_71 R_wl
Cwl_26_71 word26_71 gnd C_wl
Rw27_71 word27_71 word26_71 R_wl
Cwl_27_71 word27_71 gnd C_wl
Rw28_71 word28_71 word27_71 R_wl
Cwl_28_71 word28_71 gnd C_wl
Rw29_71 word29_71 word28_71 R_wl
Cwl_29_71 word29_71 gnd C_wl
Rw30_71 word30_71 word29_71 R_wl
Cwl_30_71 word30_71 gnd C_wl
Rw31_71 word31_71 word30_71 R_wl
Cwl_31_71 word31_71 gnd C_wl
Rw32_71 word32_71 word31_71 R_wl
Cwl_32_71 word32_71 gnd C_wl
Rw33_71 word33_71 word32_71 R_wl
Cwl_33_71 word33_71 gnd C_wl
Rw34_71 word34_71 word33_71 R_wl
Cwl_34_71 word34_71 gnd C_wl
Rw35_71 word35_71 word34_71 R_wl
Cwl_35_71 word35_71 gnd C_wl
Rw36_71 word36_71 word35_71 R_wl
Cwl_36_71 word36_71 gnd C_wl
Rw37_71 word37_71 word36_71 R_wl
Cwl_37_71 word37_71 gnd C_wl
Rw38_71 word38_71 word37_71 R_wl
Cwl_38_71 word38_71 gnd C_wl
Rw39_71 word39_71 word38_71 R_wl
Cwl_39_71 word39_71 gnd C_wl
Rw40_71 word40_71 word39_71 R_wl
Cwl_40_71 word40_71 gnd C_wl
Rw41_71 word41_71 word40_71 R_wl
Cwl_41_71 word41_71 gnd C_wl
Rw42_71 word42_71 word41_71 R_wl
Cwl_42_71 word42_71 gnd C_wl
Rw43_71 word43_71 word42_71 R_wl
Cwl_43_71 word43_71 gnd C_wl
Rw44_71 word44_71 word43_71 R_wl
Cwl_44_71 word44_71 gnd C_wl
Rw45_71 word45_71 word44_71 R_wl
Cwl_45_71 word45_71 gnd C_wl
Rw46_71 word46_71 word45_71 R_wl
Cwl_46_71 word46_71 gnd C_wl
Rw47_71 word47_71 word46_71 R_wl
Cwl_47_71 word47_71 gnd C_wl
Rw48_71 word48_71 word47_71 R_wl
Cwl_48_71 word48_71 gnd C_wl
Rw49_71 word49_71 word48_71 R_wl
Cwl_49_71 word49_71 gnd C_wl
Rw50_71 word50_71 word49_71 R_wl
Cwl_50_71 word50_71 gnd C_wl
Rw51_71 word51_71 word50_71 R_wl
Cwl_51_71 word51_71 gnd C_wl
Rw52_71 word52_71 word51_71 R_wl
Cwl_52_71 word52_71 gnd C_wl
Rw53_71 word53_71 word52_71 R_wl
Cwl_53_71 word53_71 gnd C_wl
Rw54_71 word54_71 word53_71 R_wl
Cwl_54_71 word54_71 gnd C_wl
Rw55_71 word55_71 word54_71 R_wl
Cwl_55_71 word55_71 gnd C_wl
Rw56_71 word56_71 word55_71 R_wl
Cwl_56_71 word56_71 gnd C_wl
Rw57_71 word57_71 word56_71 R_wl
Cwl_57_71 word57_71 gnd C_wl
Rw58_71 word58_71 word57_71 R_wl
Cwl_58_71 word58_71 gnd C_wl
Rw59_71 word59_71 word58_71 R_wl
Cwl_59_71 word59_71 gnd C_wl
Rw60_71 word60_71 word59_71 R_wl
Cwl_60_71 word60_71 gnd C_wl
Rw61_71 word61_71 word60_71 R_wl
Cwl_61_71 word61_71 gnd C_wl
Rw62_71 word62_71 word61_71 R_wl
Cwl_62_71 word62_71 gnd C_wl
Rw63_71 word63_71 word62_71 R_wl
Cwl_63_71 word63_71 gnd C_wl
Rw64_71 word64_71 word63_71 R_wl
Cwl_64_71 word64_71 gnd C_wl
Rw65_71 word65_71 word64_71 R_wl
Cwl_65_71 word65_71 gnd C_wl
Rw66_71 word66_71 word65_71 R_wl
Cwl_66_71 word66_71 gnd C_wl
Rw67_71 word67_71 word66_71 R_wl
Cwl_67_71 word67_71 gnd C_wl
Rw68_71 word68_71 word67_71 R_wl
Cwl_68_71 word68_71 gnd C_wl
Rw69_71 word69_71 word68_71 R_wl
Cwl_69_71 word69_71 gnd C_wl
Rw70_71 word70_71 word69_71 R_wl
Cwl_70_71 word70_71 gnd C_wl
Rw71_71 word71_71 word70_71 R_wl
Cwl_71_71 word71_71 gnd C_wl
Rw72_71 word72_71 word71_71 R_wl
Cwl_72_71 word72_71 gnd C_wl
Rw73_71 word73_71 word72_71 R_wl
Cwl_73_71 word73_71 gnd C_wl
Rw74_71 word74_71 word73_71 R_wl
Cwl_74_71 word74_71 gnd C_wl
Rw75_71 word75_71 word74_71 R_wl
Cwl_75_71 word75_71 gnd C_wl
Rw76_71 word76_71 word75_71 R_wl
Cwl_76_71 word76_71 gnd C_wl
Rw77_71 word77_71 word76_71 R_wl
Cwl_77_71 word77_71 gnd C_wl
Rw78_71 word78_71 word77_71 R_wl
Cwl_78_71 word78_71 gnd C_wl
Rw79_71 word79_71 word78_71 R_wl
Cwl_79_71 word79_71 gnd C_wl
Rw80_71 word80_71 word79_71 R_wl
Cwl_80_71 word80_71 gnd C_wl
Rw81_71 word81_71 word80_71 R_wl
Cwl_81_71 word81_71 gnd C_wl
Rw82_71 word82_71 word81_71 R_wl
Cwl_82_71 word82_71 gnd C_wl
Rw83_71 word83_71 word82_71 R_wl
Cwl_83_71 word83_71 gnd C_wl
Rw84_71 word84_71 word83_71 R_wl
Cwl_84_71 word84_71 gnd C_wl
Rw85_71 word85_71 word84_71 R_wl
Cwl_85_71 word85_71 gnd C_wl
Rw86_71 word86_71 word85_71 R_wl
Cwl_86_71 word86_71 gnd C_wl
Rw87_71 word87_71 word86_71 R_wl
Cwl_87_71 word87_71 gnd C_wl
Rw88_71 word88_71 word87_71 R_wl
Cwl_88_71 word88_71 gnd C_wl
Rw89_71 word89_71 word88_71 R_wl
Cwl_89_71 word89_71 gnd C_wl
Rw90_71 word90_71 word89_71 R_wl
Cwl_90_71 word90_71 gnd C_wl
Rw91_71 word91_71 word90_71 R_wl
Cwl_91_71 word91_71 gnd C_wl
Rw92_71 word92_71 word91_71 R_wl
Cwl_92_71 word92_71 gnd C_wl
Rw93_71 word93_71 word92_71 R_wl
Cwl_93_71 word93_71 gnd C_wl
Rw94_71 word94_71 word93_71 R_wl
Cwl_94_71 word94_71 gnd C_wl
Rw95_71 word95_71 word94_71 R_wl
Cwl_95_71 word95_71 gnd C_wl
Rw96_71 word96_71 word95_71 R_wl
Cwl_96_71 word96_71 gnd C_wl
Rw97_71 word97_71 word96_71 R_wl
Cwl_97_71 word97_71 gnd C_wl
Rw98_71 word98_71 word97_71 R_wl
Cwl_98_71 word98_71 gnd C_wl
Rw99_71 word99_71 word98_71 R_wl
Cwl_99_71 word99_71 gnd C_wl
Vwl_72 word_72 0 0
Rw0_72 word_72 word0_72 R_wl
Cwl_0_72 word0_72 gnd C_wl
Rw1_72 word1_72 word0_72 R_wl
Cwl_1_72 word1_72 gnd C_wl
Rw2_72 word2_72 word1_72 R_wl
Cwl_2_72 word2_72 gnd C_wl
Rw3_72 word3_72 word2_72 R_wl
Cwl_3_72 word3_72 gnd C_wl
Rw4_72 word4_72 word3_72 R_wl
Cwl_4_72 word4_72 gnd C_wl
Rw5_72 word5_72 word4_72 R_wl
Cwl_5_72 word5_72 gnd C_wl
Rw6_72 word6_72 word5_72 R_wl
Cwl_6_72 word6_72 gnd C_wl
Rw7_72 word7_72 word6_72 R_wl
Cwl_7_72 word7_72 gnd C_wl
Rw8_72 word8_72 word7_72 R_wl
Cwl_8_72 word8_72 gnd C_wl
Rw9_72 word9_72 word8_72 R_wl
Cwl_9_72 word9_72 gnd C_wl
Rw10_72 word10_72 word9_72 R_wl
Cwl_10_72 word10_72 gnd C_wl
Rw11_72 word11_72 word10_72 R_wl
Cwl_11_72 word11_72 gnd C_wl
Rw12_72 word12_72 word11_72 R_wl
Cwl_12_72 word12_72 gnd C_wl
Rw13_72 word13_72 word12_72 R_wl
Cwl_13_72 word13_72 gnd C_wl
Rw14_72 word14_72 word13_72 R_wl
Cwl_14_72 word14_72 gnd C_wl
Rw15_72 word15_72 word14_72 R_wl
Cwl_15_72 word15_72 gnd C_wl
Rw16_72 word16_72 word15_72 R_wl
Cwl_16_72 word16_72 gnd C_wl
Rw17_72 word17_72 word16_72 R_wl
Cwl_17_72 word17_72 gnd C_wl
Rw18_72 word18_72 word17_72 R_wl
Cwl_18_72 word18_72 gnd C_wl
Rw19_72 word19_72 word18_72 R_wl
Cwl_19_72 word19_72 gnd C_wl
Rw20_72 word20_72 word19_72 R_wl
Cwl_20_72 word20_72 gnd C_wl
Rw21_72 word21_72 word20_72 R_wl
Cwl_21_72 word21_72 gnd C_wl
Rw22_72 word22_72 word21_72 R_wl
Cwl_22_72 word22_72 gnd C_wl
Rw23_72 word23_72 word22_72 R_wl
Cwl_23_72 word23_72 gnd C_wl
Rw24_72 word24_72 word23_72 R_wl
Cwl_24_72 word24_72 gnd C_wl
Rw25_72 word25_72 word24_72 R_wl
Cwl_25_72 word25_72 gnd C_wl
Rw26_72 word26_72 word25_72 R_wl
Cwl_26_72 word26_72 gnd C_wl
Rw27_72 word27_72 word26_72 R_wl
Cwl_27_72 word27_72 gnd C_wl
Rw28_72 word28_72 word27_72 R_wl
Cwl_28_72 word28_72 gnd C_wl
Rw29_72 word29_72 word28_72 R_wl
Cwl_29_72 word29_72 gnd C_wl
Rw30_72 word30_72 word29_72 R_wl
Cwl_30_72 word30_72 gnd C_wl
Rw31_72 word31_72 word30_72 R_wl
Cwl_31_72 word31_72 gnd C_wl
Rw32_72 word32_72 word31_72 R_wl
Cwl_32_72 word32_72 gnd C_wl
Rw33_72 word33_72 word32_72 R_wl
Cwl_33_72 word33_72 gnd C_wl
Rw34_72 word34_72 word33_72 R_wl
Cwl_34_72 word34_72 gnd C_wl
Rw35_72 word35_72 word34_72 R_wl
Cwl_35_72 word35_72 gnd C_wl
Rw36_72 word36_72 word35_72 R_wl
Cwl_36_72 word36_72 gnd C_wl
Rw37_72 word37_72 word36_72 R_wl
Cwl_37_72 word37_72 gnd C_wl
Rw38_72 word38_72 word37_72 R_wl
Cwl_38_72 word38_72 gnd C_wl
Rw39_72 word39_72 word38_72 R_wl
Cwl_39_72 word39_72 gnd C_wl
Rw40_72 word40_72 word39_72 R_wl
Cwl_40_72 word40_72 gnd C_wl
Rw41_72 word41_72 word40_72 R_wl
Cwl_41_72 word41_72 gnd C_wl
Rw42_72 word42_72 word41_72 R_wl
Cwl_42_72 word42_72 gnd C_wl
Rw43_72 word43_72 word42_72 R_wl
Cwl_43_72 word43_72 gnd C_wl
Rw44_72 word44_72 word43_72 R_wl
Cwl_44_72 word44_72 gnd C_wl
Rw45_72 word45_72 word44_72 R_wl
Cwl_45_72 word45_72 gnd C_wl
Rw46_72 word46_72 word45_72 R_wl
Cwl_46_72 word46_72 gnd C_wl
Rw47_72 word47_72 word46_72 R_wl
Cwl_47_72 word47_72 gnd C_wl
Rw48_72 word48_72 word47_72 R_wl
Cwl_48_72 word48_72 gnd C_wl
Rw49_72 word49_72 word48_72 R_wl
Cwl_49_72 word49_72 gnd C_wl
Rw50_72 word50_72 word49_72 R_wl
Cwl_50_72 word50_72 gnd C_wl
Rw51_72 word51_72 word50_72 R_wl
Cwl_51_72 word51_72 gnd C_wl
Rw52_72 word52_72 word51_72 R_wl
Cwl_52_72 word52_72 gnd C_wl
Rw53_72 word53_72 word52_72 R_wl
Cwl_53_72 word53_72 gnd C_wl
Rw54_72 word54_72 word53_72 R_wl
Cwl_54_72 word54_72 gnd C_wl
Rw55_72 word55_72 word54_72 R_wl
Cwl_55_72 word55_72 gnd C_wl
Rw56_72 word56_72 word55_72 R_wl
Cwl_56_72 word56_72 gnd C_wl
Rw57_72 word57_72 word56_72 R_wl
Cwl_57_72 word57_72 gnd C_wl
Rw58_72 word58_72 word57_72 R_wl
Cwl_58_72 word58_72 gnd C_wl
Rw59_72 word59_72 word58_72 R_wl
Cwl_59_72 word59_72 gnd C_wl
Rw60_72 word60_72 word59_72 R_wl
Cwl_60_72 word60_72 gnd C_wl
Rw61_72 word61_72 word60_72 R_wl
Cwl_61_72 word61_72 gnd C_wl
Rw62_72 word62_72 word61_72 R_wl
Cwl_62_72 word62_72 gnd C_wl
Rw63_72 word63_72 word62_72 R_wl
Cwl_63_72 word63_72 gnd C_wl
Rw64_72 word64_72 word63_72 R_wl
Cwl_64_72 word64_72 gnd C_wl
Rw65_72 word65_72 word64_72 R_wl
Cwl_65_72 word65_72 gnd C_wl
Rw66_72 word66_72 word65_72 R_wl
Cwl_66_72 word66_72 gnd C_wl
Rw67_72 word67_72 word66_72 R_wl
Cwl_67_72 word67_72 gnd C_wl
Rw68_72 word68_72 word67_72 R_wl
Cwl_68_72 word68_72 gnd C_wl
Rw69_72 word69_72 word68_72 R_wl
Cwl_69_72 word69_72 gnd C_wl
Rw70_72 word70_72 word69_72 R_wl
Cwl_70_72 word70_72 gnd C_wl
Rw71_72 word71_72 word70_72 R_wl
Cwl_71_72 word71_72 gnd C_wl
Rw72_72 word72_72 word71_72 R_wl
Cwl_72_72 word72_72 gnd C_wl
Rw73_72 word73_72 word72_72 R_wl
Cwl_73_72 word73_72 gnd C_wl
Rw74_72 word74_72 word73_72 R_wl
Cwl_74_72 word74_72 gnd C_wl
Rw75_72 word75_72 word74_72 R_wl
Cwl_75_72 word75_72 gnd C_wl
Rw76_72 word76_72 word75_72 R_wl
Cwl_76_72 word76_72 gnd C_wl
Rw77_72 word77_72 word76_72 R_wl
Cwl_77_72 word77_72 gnd C_wl
Rw78_72 word78_72 word77_72 R_wl
Cwl_78_72 word78_72 gnd C_wl
Rw79_72 word79_72 word78_72 R_wl
Cwl_79_72 word79_72 gnd C_wl
Rw80_72 word80_72 word79_72 R_wl
Cwl_80_72 word80_72 gnd C_wl
Rw81_72 word81_72 word80_72 R_wl
Cwl_81_72 word81_72 gnd C_wl
Rw82_72 word82_72 word81_72 R_wl
Cwl_82_72 word82_72 gnd C_wl
Rw83_72 word83_72 word82_72 R_wl
Cwl_83_72 word83_72 gnd C_wl
Rw84_72 word84_72 word83_72 R_wl
Cwl_84_72 word84_72 gnd C_wl
Rw85_72 word85_72 word84_72 R_wl
Cwl_85_72 word85_72 gnd C_wl
Rw86_72 word86_72 word85_72 R_wl
Cwl_86_72 word86_72 gnd C_wl
Rw87_72 word87_72 word86_72 R_wl
Cwl_87_72 word87_72 gnd C_wl
Rw88_72 word88_72 word87_72 R_wl
Cwl_88_72 word88_72 gnd C_wl
Rw89_72 word89_72 word88_72 R_wl
Cwl_89_72 word89_72 gnd C_wl
Rw90_72 word90_72 word89_72 R_wl
Cwl_90_72 word90_72 gnd C_wl
Rw91_72 word91_72 word90_72 R_wl
Cwl_91_72 word91_72 gnd C_wl
Rw92_72 word92_72 word91_72 R_wl
Cwl_92_72 word92_72 gnd C_wl
Rw93_72 word93_72 word92_72 R_wl
Cwl_93_72 word93_72 gnd C_wl
Rw94_72 word94_72 word93_72 R_wl
Cwl_94_72 word94_72 gnd C_wl
Rw95_72 word95_72 word94_72 R_wl
Cwl_95_72 word95_72 gnd C_wl
Rw96_72 word96_72 word95_72 R_wl
Cwl_96_72 word96_72 gnd C_wl
Rw97_72 word97_72 word96_72 R_wl
Cwl_97_72 word97_72 gnd C_wl
Rw98_72 word98_72 word97_72 R_wl
Cwl_98_72 word98_72 gnd C_wl
Rw99_72 word99_72 word98_72 R_wl
Cwl_99_72 word99_72 gnd C_wl
Vwl_73 word_73 0 0
Rw0_73 word_73 word0_73 R_wl
Cwl_0_73 word0_73 gnd C_wl
Rw1_73 word1_73 word0_73 R_wl
Cwl_1_73 word1_73 gnd C_wl
Rw2_73 word2_73 word1_73 R_wl
Cwl_2_73 word2_73 gnd C_wl
Rw3_73 word3_73 word2_73 R_wl
Cwl_3_73 word3_73 gnd C_wl
Rw4_73 word4_73 word3_73 R_wl
Cwl_4_73 word4_73 gnd C_wl
Rw5_73 word5_73 word4_73 R_wl
Cwl_5_73 word5_73 gnd C_wl
Rw6_73 word6_73 word5_73 R_wl
Cwl_6_73 word6_73 gnd C_wl
Rw7_73 word7_73 word6_73 R_wl
Cwl_7_73 word7_73 gnd C_wl
Rw8_73 word8_73 word7_73 R_wl
Cwl_8_73 word8_73 gnd C_wl
Rw9_73 word9_73 word8_73 R_wl
Cwl_9_73 word9_73 gnd C_wl
Rw10_73 word10_73 word9_73 R_wl
Cwl_10_73 word10_73 gnd C_wl
Rw11_73 word11_73 word10_73 R_wl
Cwl_11_73 word11_73 gnd C_wl
Rw12_73 word12_73 word11_73 R_wl
Cwl_12_73 word12_73 gnd C_wl
Rw13_73 word13_73 word12_73 R_wl
Cwl_13_73 word13_73 gnd C_wl
Rw14_73 word14_73 word13_73 R_wl
Cwl_14_73 word14_73 gnd C_wl
Rw15_73 word15_73 word14_73 R_wl
Cwl_15_73 word15_73 gnd C_wl
Rw16_73 word16_73 word15_73 R_wl
Cwl_16_73 word16_73 gnd C_wl
Rw17_73 word17_73 word16_73 R_wl
Cwl_17_73 word17_73 gnd C_wl
Rw18_73 word18_73 word17_73 R_wl
Cwl_18_73 word18_73 gnd C_wl
Rw19_73 word19_73 word18_73 R_wl
Cwl_19_73 word19_73 gnd C_wl
Rw20_73 word20_73 word19_73 R_wl
Cwl_20_73 word20_73 gnd C_wl
Rw21_73 word21_73 word20_73 R_wl
Cwl_21_73 word21_73 gnd C_wl
Rw22_73 word22_73 word21_73 R_wl
Cwl_22_73 word22_73 gnd C_wl
Rw23_73 word23_73 word22_73 R_wl
Cwl_23_73 word23_73 gnd C_wl
Rw24_73 word24_73 word23_73 R_wl
Cwl_24_73 word24_73 gnd C_wl
Rw25_73 word25_73 word24_73 R_wl
Cwl_25_73 word25_73 gnd C_wl
Rw26_73 word26_73 word25_73 R_wl
Cwl_26_73 word26_73 gnd C_wl
Rw27_73 word27_73 word26_73 R_wl
Cwl_27_73 word27_73 gnd C_wl
Rw28_73 word28_73 word27_73 R_wl
Cwl_28_73 word28_73 gnd C_wl
Rw29_73 word29_73 word28_73 R_wl
Cwl_29_73 word29_73 gnd C_wl
Rw30_73 word30_73 word29_73 R_wl
Cwl_30_73 word30_73 gnd C_wl
Rw31_73 word31_73 word30_73 R_wl
Cwl_31_73 word31_73 gnd C_wl
Rw32_73 word32_73 word31_73 R_wl
Cwl_32_73 word32_73 gnd C_wl
Rw33_73 word33_73 word32_73 R_wl
Cwl_33_73 word33_73 gnd C_wl
Rw34_73 word34_73 word33_73 R_wl
Cwl_34_73 word34_73 gnd C_wl
Rw35_73 word35_73 word34_73 R_wl
Cwl_35_73 word35_73 gnd C_wl
Rw36_73 word36_73 word35_73 R_wl
Cwl_36_73 word36_73 gnd C_wl
Rw37_73 word37_73 word36_73 R_wl
Cwl_37_73 word37_73 gnd C_wl
Rw38_73 word38_73 word37_73 R_wl
Cwl_38_73 word38_73 gnd C_wl
Rw39_73 word39_73 word38_73 R_wl
Cwl_39_73 word39_73 gnd C_wl
Rw40_73 word40_73 word39_73 R_wl
Cwl_40_73 word40_73 gnd C_wl
Rw41_73 word41_73 word40_73 R_wl
Cwl_41_73 word41_73 gnd C_wl
Rw42_73 word42_73 word41_73 R_wl
Cwl_42_73 word42_73 gnd C_wl
Rw43_73 word43_73 word42_73 R_wl
Cwl_43_73 word43_73 gnd C_wl
Rw44_73 word44_73 word43_73 R_wl
Cwl_44_73 word44_73 gnd C_wl
Rw45_73 word45_73 word44_73 R_wl
Cwl_45_73 word45_73 gnd C_wl
Rw46_73 word46_73 word45_73 R_wl
Cwl_46_73 word46_73 gnd C_wl
Rw47_73 word47_73 word46_73 R_wl
Cwl_47_73 word47_73 gnd C_wl
Rw48_73 word48_73 word47_73 R_wl
Cwl_48_73 word48_73 gnd C_wl
Rw49_73 word49_73 word48_73 R_wl
Cwl_49_73 word49_73 gnd C_wl
Rw50_73 word50_73 word49_73 R_wl
Cwl_50_73 word50_73 gnd C_wl
Rw51_73 word51_73 word50_73 R_wl
Cwl_51_73 word51_73 gnd C_wl
Rw52_73 word52_73 word51_73 R_wl
Cwl_52_73 word52_73 gnd C_wl
Rw53_73 word53_73 word52_73 R_wl
Cwl_53_73 word53_73 gnd C_wl
Rw54_73 word54_73 word53_73 R_wl
Cwl_54_73 word54_73 gnd C_wl
Rw55_73 word55_73 word54_73 R_wl
Cwl_55_73 word55_73 gnd C_wl
Rw56_73 word56_73 word55_73 R_wl
Cwl_56_73 word56_73 gnd C_wl
Rw57_73 word57_73 word56_73 R_wl
Cwl_57_73 word57_73 gnd C_wl
Rw58_73 word58_73 word57_73 R_wl
Cwl_58_73 word58_73 gnd C_wl
Rw59_73 word59_73 word58_73 R_wl
Cwl_59_73 word59_73 gnd C_wl
Rw60_73 word60_73 word59_73 R_wl
Cwl_60_73 word60_73 gnd C_wl
Rw61_73 word61_73 word60_73 R_wl
Cwl_61_73 word61_73 gnd C_wl
Rw62_73 word62_73 word61_73 R_wl
Cwl_62_73 word62_73 gnd C_wl
Rw63_73 word63_73 word62_73 R_wl
Cwl_63_73 word63_73 gnd C_wl
Rw64_73 word64_73 word63_73 R_wl
Cwl_64_73 word64_73 gnd C_wl
Rw65_73 word65_73 word64_73 R_wl
Cwl_65_73 word65_73 gnd C_wl
Rw66_73 word66_73 word65_73 R_wl
Cwl_66_73 word66_73 gnd C_wl
Rw67_73 word67_73 word66_73 R_wl
Cwl_67_73 word67_73 gnd C_wl
Rw68_73 word68_73 word67_73 R_wl
Cwl_68_73 word68_73 gnd C_wl
Rw69_73 word69_73 word68_73 R_wl
Cwl_69_73 word69_73 gnd C_wl
Rw70_73 word70_73 word69_73 R_wl
Cwl_70_73 word70_73 gnd C_wl
Rw71_73 word71_73 word70_73 R_wl
Cwl_71_73 word71_73 gnd C_wl
Rw72_73 word72_73 word71_73 R_wl
Cwl_72_73 word72_73 gnd C_wl
Rw73_73 word73_73 word72_73 R_wl
Cwl_73_73 word73_73 gnd C_wl
Rw74_73 word74_73 word73_73 R_wl
Cwl_74_73 word74_73 gnd C_wl
Rw75_73 word75_73 word74_73 R_wl
Cwl_75_73 word75_73 gnd C_wl
Rw76_73 word76_73 word75_73 R_wl
Cwl_76_73 word76_73 gnd C_wl
Rw77_73 word77_73 word76_73 R_wl
Cwl_77_73 word77_73 gnd C_wl
Rw78_73 word78_73 word77_73 R_wl
Cwl_78_73 word78_73 gnd C_wl
Rw79_73 word79_73 word78_73 R_wl
Cwl_79_73 word79_73 gnd C_wl
Rw80_73 word80_73 word79_73 R_wl
Cwl_80_73 word80_73 gnd C_wl
Rw81_73 word81_73 word80_73 R_wl
Cwl_81_73 word81_73 gnd C_wl
Rw82_73 word82_73 word81_73 R_wl
Cwl_82_73 word82_73 gnd C_wl
Rw83_73 word83_73 word82_73 R_wl
Cwl_83_73 word83_73 gnd C_wl
Rw84_73 word84_73 word83_73 R_wl
Cwl_84_73 word84_73 gnd C_wl
Rw85_73 word85_73 word84_73 R_wl
Cwl_85_73 word85_73 gnd C_wl
Rw86_73 word86_73 word85_73 R_wl
Cwl_86_73 word86_73 gnd C_wl
Rw87_73 word87_73 word86_73 R_wl
Cwl_87_73 word87_73 gnd C_wl
Rw88_73 word88_73 word87_73 R_wl
Cwl_88_73 word88_73 gnd C_wl
Rw89_73 word89_73 word88_73 R_wl
Cwl_89_73 word89_73 gnd C_wl
Rw90_73 word90_73 word89_73 R_wl
Cwl_90_73 word90_73 gnd C_wl
Rw91_73 word91_73 word90_73 R_wl
Cwl_91_73 word91_73 gnd C_wl
Rw92_73 word92_73 word91_73 R_wl
Cwl_92_73 word92_73 gnd C_wl
Rw93_73 word93_73 word92_73 R_wl
Cwl_93_73 word93_73 gnd C_wl
Rw94_73 word94_73 word93_73 R_wl
Cwl_94_73 word94_73 gnd C_wl
Rw95_73 word95_73 word94_73 R_wl
Cwl_95_73 word95_73 gnd C_wl
Rw96_73 word96_73 word95_73 R_wl
Cwl_96_73 word96_73 gnd C_wl
Rw97_73 word97_73 word96_73 R_wl
Cwl_97_73 word97_73 gnd C_wl
Rw98_73 word98_73 word97_73 R_wl
Cwl_98_73 word98_73 gnd C_wl
Rw99_73 word99_73 word98_73 R_wl
Cwl_99_73 word99_73 gnd C_wl
Vwl_74 word_74 0 0
Rw0_74 word_74 word0_74 R_wl
Cwl_0_74 word0_74 gnd C_wl
Rw1_74 word1_74 word0_74 R_wl
Cwl_1_74 word1_74 gnd C_wl
Rw2_74 word2_74 word1_74 R_wl
Cwl_2_74 word2_74 gnd C_wl
Rw3_74 word3_74 word2_74 R_wl
Cwl_3_74 word3_74 gnd C_wl
Rw4_74 word4_74 word3_74 R_wl
Cwl_4_74 word4_74 gnd C_wl
Rw5_74 word5_74 word4_74 R_wl
Cwl_5_74 word5_74 gnd C_wl
Rw6_74 word6_74 word5_74 R_wl
Cwl_6_74 word6_74 gnd C_wl
Rw7_74 word7_74 word6_74 R_wl
Cwl_7_74 word7_74 gnd C_wl
Rw8_74 word8_74 word7_74 R_wl
Cwl_8_74 word8_74 gnd C_wl
Rw9_74 word9_74 word8_74 R_wl
Cwl_9_74 word9_74 gnd C_wl
Rw10_74 word10_74 word9_74 R_wl
Cwl_10_74 word10_74 gnd C_wl
Rw11_74 word11_74 word10_74 R_wl
Cwl_11_74 word11_74 gnd C_wl
Rw12_74 word12_74 word11_74 R_wl
Cwl_12_74 word12_74 gnd C_wl
Rw13_74 word13_74 word12_74 R_wl
Cwl_13_74 word13_74 gnd C_wl
Rw14_74 word14_74 word13_74 R_wl
Cwl_14_74 word14_74 gnd C_wl
Rw15_74 word15_74 word14_74 R_wl
Cwl_15_74 word15_74 gnd C_wl
Rw16_74 word16_74 word15_74 R_wl
Cwl_16_74 word16_74 gnd C_wl
Rw17_74 word17_74 word16_74 R_wl
Cwl_17_74 word17_74 gnd C_wl
Rw18_74 word18_74 word17_74 R_wl
Cwl_18_74 word18_74 gnd C_wl
Rw19_74 word19_74 word18_74 R_wl
Cwl_19_74 word19_74 gnd C_wl
Rw20_74 word20_74 word19_74 R_wl
Cwl_20_74 word20_74 gnd C_wl
Rw21_74 word21_74 word20_74 R_wl
Cwl_21_74 word21_74 gnd C_wl
Rw22_74 word22_74 word21_74 R_wl
Cwl_22_74 word22_74 gnd C_wl
Rw23_74 word23_74 word22_74 R_wl
Cwl_23_74 word23_74 gnd C_wl
Rw24_74 word24_74 word23_74 R_wl
Cwl_24_74 word24_74 gnd C_wl
Rw25_74 word25_74 word24_74 R_wl
Cwl_25_74 word25_74 gnd C_wl
Rw26_74 word26_74 word25_74 R_wl
Cwl_26_74 word26_74 gnd C_wl
Rw27_74 word27_74 word26_74 R_wl
Cwl_27_74 word27_74 gnd C_wl
Rw28_74 word28_74 word27_74 R_wl
Cwl_28_74 word28_74 gnd C_wl
Rw29_74 word29_74 word28_74 R_wl
Cwl_29_74 word29_74 gnd C_wl
Rw30_74 word30_74 word29_74 R_wl
Cwl_30_74 word30_74 gnd C_wl
Rw31_74 word31_74 word30_74 R_wl
Cwl_31_74 word31_74 gnd C_wl
Rw32_74 word32_74 word31_74 R_wl
Cwl_32_74 word32_74 gnd C_wl
Rw33_74 word33_74 word32_74 R_wl
Cwl_33_74 word33_74 gnd C_wl
Rw34_74 word34_74 word33_74 R_wl
Cwl_34_74 word34_74 gnd C_wl
Rw35_74 word35_74 word34_74 R_wl
Cwl_35_74 word35_74 gnd C_wl
Rw36_74 word36_74 word35_74 R_wl
Cwl_36_74 word36_74 gnd C_wl
Rw37_74 word37_74 word36_74 R_wl
Cwl_37_74 word37_74 gnd C_wl
Rw38_74 word38_74 word37_74 R_wl
Cwl_38_74 word38_74 gnd C_wl
Rw39_74 word39_74 word38_74 R_wl
Cwl_39_74 word39_74 gnd C_wl
Rw40_74 word40_74 word39_74 R_wl
Cwl_40_74 word40_74 gnd C_wl
Rw41_74 word41_74 word40_74 R_wl
Cwl_41_74 word41_74 gnd C_wl
Rw42_74 word42_74 word41_74 R_wl
Cwl_42_74 word42_74 gnd C_wl
Rw43_74 word43_74 word42_74 R_wl
Cwl_43_74 word43_74 gnd C_wl
Rw44_74 word44_74 word43_74 R_wl
Cwl_44_74 word44_74 gnd C_wl
Rw45_74 word45_74 word44_74 R_wl
Cwl_45_74 word45_74 gnd C_wl
Rw46_74 word46_74 word45_74 R_wl
Cwl_46_74 word46_74 gnd C_wl
Rw47_74 word47_74 word46_74 R_wl
Cwl_47_74 word47_74 gnd C_wl
Rw48_74 word48_74 word47_74 R_wl
Cwl_48_74 word48_74 gnd C_wl
Rw49_74 word49_74 word48_74 R_wl
Cwl_49_74 word49_74 gnd C_wl
Rw50_74 word50_74 word49_74 R_wl
Cwl_50_74 word50_74 gnd C_wl
Rw51_74 word51_74 word50_74 R_wl
Cwl_51_74 word51_74 gnd C_wl
Rw52_74 word52_74 word51_74 R_wl
Cwl_52_74 word52_74 gnd C_wl
Rw53_74 word53_74 word52_74 R_wl
Cwl_53_74 word53_74 gnd C_wl
Rw54_74 word54_74 word53_74 R_wl
Cwl_54_74 word54_74 gnd C_wl
Rw55_74 word55_74 word54_74 R_wl
Cwl_55_74 word55_74 gnd C_wl
Rw56_74 word56_74 word55_74 R_wl
Cwl_56_74 word56_74 gnd C_wl
Rw57_74 word57_74 word56_74 R_wl
Cwl_57_74 word57_74 gnd C_wl
Rw58_74 word58_74 word57_74 R_wl
Cwl_58_74 word58_74 gnd C_wl
Rw59_74 word59_74 word58_74 R_wl
Cwl_59_74 word59_74 gnd C_wl
Rw60_74 word60_74 word59_74 R_wl
Cwl_60_74 word60_74 gnd C_wl
Rw61_74 word61_74 word60_74 R_wl
Cwl_61_74 word61_74 gnd C_wl
Rw62_74 word62_74 word61_74 R_wl
Cwl_62_74 word62_74 gnd C_wl
Rw63_74 word63_74 word62_74 R_wl
Cwl_63_74 word63_74 gnd C_wl
Rw64_74 word64_74 word63_74 R_wl
Cwl_64_74 word64_74 gnd C_wl
Rw65_74 word65_74 word64_74 R_wl
Cwl_65_74 word65_74 gnd C_wl
Rw66_74 word66_74 word65_74 R_wl
Cwl_66_74 word66_74 gnd C_wl
Rw67_74 word67_74 word66_74 R_wl
Cwl_67_74 word67_74 gnd C_wl
Rw68_74 word68_74 word67_74 R_wl
Cwl_68_74 word68_74 gnd C_wl
Rw69_74 word69_74 word68_74 R_wl
Cwl_69_74 word69_74 gnd C_wl
Rw70_74 word70_74 word69_74 R_wl
Cwl_70_74 word70_74 gnd C_wl
Rw71_74 word71_74 word70_74 R_wl
Cwl_71_74 word71_74 gnd C_wl
Rw72_74 word72_74 word71_74 R_wl
Cwl_72_74 word72_74 gnd C_wl
Rw73_74 word73_74 word72_74 R_wl
Cwl_73_74 word73_74 gnd C_wl
Rw74_74 word74_74 word73_74 R_wl
Cwl_74_74 word74_74 gnd C_wl
Rw75_74 word75_74 word74_74 R_wl
Cwl_75_74 word75_74 gnd C_wl
Rw76_74 word76_74 word75_74 R_wl
Cwl_76_74 word76_74 gnd C_wl
Rw77_74 word77_74 word76_74 R_wl
Cwl_77_74 word77_74 gnd C_wl
Rw78_74 word78_74 word77_74 R_wl
Cwl_78_74 word78_74 gnd C_wl
Rw79_74 word79_74 word78_74 R_wl
Cwl_79_74 word79_74 gnd C_wl
Rw80_74 word80_74 word79_74 R_wl
Cwl_80_74 word80_74 gnd C_wl
Rw81_74 word81_74 word80_74 R_wl
Cwl_81_74 word81_74 gnd C_wl
Rw82_74 word82_74 word81_74 R_wl
Cwl_82_74 word82_74 gnd C_wl
Rw83_74 word83_74 word82_74 R_wl
Cwl_83_74 word83_74 gnd C_wl
Rw84_74 word84_74 word83_74 R_wl
Cwl_84_74 word84_74 gnd C_wl
Rw85_74 word85_74 word84_74 R_wl
Cwl_85_74 word85_74 gnd C_wl
Rw86_74 word86_74 word85_74 R_wl
Cwl_86_74 word86_74 gnd C_wl
Rw87_74 word87_74 word86_74 R_wl
Cwl_87_74 word87_74 gnd C_wl
Rw88_74 word88_74 word87_74 R_wl
Cwl_88_74 word88_74 gnd C_wl
Rw89_74 word89_74 word88_74 R_wl
Cwl_89_74 word89_74 gnd C_wl
Rw90_74 word90_74 word89_74 R_wl
Cwl_90_74 word90_74 gnd C_wl
Rw91_74 word91_74 word90_74 R_wl
Cwl_91_74 word91_74 gnd C_wl
Rw92_74 word92_74 word91_74 R_wl
Cwl_92_74 word92_74 gnd C_wl
Rw93_74 word93_74 word92_74 R_wl
Cwl_93_74 word93_74 gnd C_wl
Rw94_74 word94_74 word93_74 R_wl
Cwl_94_74 word94_74 gnd C_wl
Rw95_74 word95_74 word94_74 R_wl
Cwl_95_74 word95_74 gnd C_wl
Rw96_74 word96_74 word95_74 R_wl
Cwl_96_74 word96_74 gnd C_wl
Rw97_74 word97_74 word96_74 R_wl
Cwl_97_74 word97_74 gnd C_wl
Rw98_74 word98_74 word97_74 R_wl
Cwl_98_74 word98_74 gnd C_wl
Rw99_74 word99_74 word98_74 R_wl
Cwl_99_74 word99_74 gnd C_wl
Vwl_75 word_75 0 0
Rw0_75 word_75 word0_75 R_wl
Cwl_0_75 word0_75 gnd C_wl
Rw1_75 word1_75 word0_75 R_wl
Cwl_1_75 word1_75 gnd C_wl
Rw2_75 word2_75 word1_75 R_wl
Cwl_2_75 word2_75 gnd C_wl
Rw3_75 word3_75 word2_75 R_wl
Cwl_3_75 word3_75 gnd C_wl
Rw4_75 word4_75 word3_75 R_wl
Cwl_4_75 word4_75 gnd C_wl
Rw5_75 word5_75 word4_75 R_wl
Cwl_5_75 word5_75 gnd C_wl
Rw6_75 word6_75 word5_75 R_wl
Cwl_6_75 word6_75 gnd C_wl
Rw7_75 word7_75 word6_75 R_wl
Cwl_7_75 word7_75 gnd C_wl
Rw8_75 word8_75 word7_75 R_wl
Cwl_8_75 word8_75 gnd C_wl
Rw9_75 word9_75 word8_75 R_wl
Cwl_9_75 word9_75 gnd C_wl
Rw10_75 word10_75 word9_75 R_wl
Cwl_10_75 word10_75 gnd C_wl
Rw11_75 word11_75 word10_75 R_wl
Cwl_11_75 word11_75 gnd C_wl
Rw12_75 word12_75 word11_75 R_wl
Cwl_12_75 word12_75 gnd C_wl
Rw13_75 word13_75 word12_75 R_wl
Cwl_13_75 word13_75 gnd C_wl
Rw14_75 word14_75 word13_75 R_wl
Cwl_14_75 word14_75 gnd C_wl
Rw15_75 word15_75 word14_75 R_wl
Cwl_15_75 word15_75 gnd C_wl
Rw16_75 word16_75 word15_75 R_wl
Cwl_16_75 word16_75 gnd C_wl
Rw17_75 word17_75 word16_75 R_wl
Cwl_17_75 word17_75 gnd C_wl
Rw18_75 word18_75 word17_75 R_wl
Cwl_18_75 word18_75 gnd C_wl
Rw19_75 word19_75 word18_75 R_wl
Cwl_19_75 word19_75 gnd C_wl
Rw20_75 word20_75 word19_75 R_wl
Cwl_20_75 word20_75 gnd C_wl
Rw21_75 word21_75 word20_75 R_wl
Cwl_21_75 word21_75 gnd C_wl
Rw22_75 word22_75 word21_75 R_wl
Cwl_22_75 word22_75 gnd C_wl
Rw23_75 word23_75 word22_75 R_wl
Cwl_23_75 word23_75 gnd C_wl
Rw24_75 word24_75 word23_75 R_wl
Cwl_24_75 word24_75 gnd C_wl
Rw25_75 word25_75 word24_75 R_wl
Cwl_25_75 word25_75 gnd C_wl
Rw26_75 word26_75 word25_75 R_wl
Cwl_26_75 word26_75 gnd C_wl
Rw27_75 word27_75 word26_75 R_wl
Cwl_27_75 word27_75 gnd C_wl
Rw28_75 word28_75 word27_75 R_wl
Cwl_28_75 word28_75 gnd C_wl
Rw29_75 word29_75 word28_75 R_wl
Cwl_29_75 word29_75 gnd C_wl
Rw30_75 word30_75 word29_75 R_wl
Cwl_30_75 word30_75 gnd C_wl
Rw31_75 word31_75 word30_75 R_wl
Cwl_31_75 word31_75 gnd C_wl
Rw32_75 word32_75 word31_75 R_wl
Cwl_32_75 word32_75 gnd C_wl
Rw33_75 word33_75 word32_75 R_wl
Cwl_33_75 word33_75 gnd C_wl
Rw34_75 word34_75 word33_75 R_wl
Cwl_34_75 word34_75 gnd C_wl
Rw35_75 word35_75 word34_75 R_wl
Cwl_35_75 word35_75 gnd C_wl
Rw36_75 word36_75 word35_75 R_wl
Cwl_36_75 word36_75 gnd C_wl
Rw37_75 word37_75 word36_75 R_wl
Cwl_37_75 word37_75 gnd C_wl
Rw38_75 word38_75 word37_75 R_wl
Cwl_38_75 word38_75 gnd C_wl
Rw39_75 word39_75 word38_75 R_wl
Cwl_39_75 word39_75 gnd C_wl
Rw40_75 word40_75 word39_75 R_wl
Cwl_40_75 word40_75 gnd C_wl
Rw41_75 word41_75 word40_75 R_wl
Cwl_41_75 word41_75 gnd C_wl
Rw42_75 word42_75 word41_75 R_wl
Cwl_42_75 word42_75 gnd C_wl
Rw43_75 word43_75 word42_75 R_wl
Cwl_43_75 word43_75 gnd C_wl
Rw44_75 word44_75 word43_75 R_wl
Cwl_44_75 word44_75 gnd C_wl
Rw45_75 word45_75 word44_75 R_wl
Cwl_45_75 word45_75 gnd C_wl
Rw46_75 word46_75 word45_75 R_wl
Cwl_46_75 word46_75 gnd C_wl
Rw47_75 word47_75 word46_75 R_wl
Cwl_47_75 word47_75 gnd C_wl
Rw48_75 word48_75 word47_75 R_wl
Cwl_48_75 word48_75 gnd C_wl
Rw49_75 word49_75 word48_75 R_wl
Cwl_49_75 word49_75 gnd C_wl
Rw50_75 word50_75 word49_75 R_wl
Cwl_50_75 word50_75 gnd C_wl
Rw51_75 word51_75 word50_75 R_wl
Cwl_51_75 word51_75 gnd C_wl
Rw52_75 word52_75 word51_75 R_wl
Cwl_52_75 word52_75 gnd C_wl
Rw53_75 word53_75 word52_75 R_wl
Cwl_53_75 word53_75 gnd C_wl
Rw54_75 word54_75 word53_75 R_wl
Cwl_54_75 word54_75 gnd C_wl
Rw55_75 word55_75 word54_75 R_wl
Cwl_55_75 word55_75 gnd C_wl
Rw56_75 word56_75 word55_75 R_wl
Cwl_56_75 word56_75 gnd C_wl
Rw57_75 word57_75 word56_75 R_wl
Cwl_57_75 word57_75 gnd C_wl
Rw58_75 word58_75 word57_75 R_wl
Cwl_58_75 word58_75 gnd C_wl
Rw59_75 word59_75 word58_75 R_wl
Cwl_59_75 word59_75 gnd C_wl
Rw60_75 word60_75 word59_75 R_wl
Cwl_60_75 word60_75 gnd C_wl
Rw61_75 word61_75 word60_75 R_wl
Cwl_61_75 word61_75 gnd C_wl
Rw62_75 word62_75 word61_75 R_wl
Cwl_62_75 word62_75 gnd C_wl
Rw63_75 word63_75 word62_75 R_wl
Cwl_63_75 word63_75 gnd C_wl
Rw64_75 word64_75 word63_75 R_wl
Cwl_64_75 word64_75 gnd C_wl
Rw65_75 word65_75 word64_75 R_wl
Cwl_65_75 word65_75 gnd C_wl
Rw66_75 word66_75 word65_75 R_wl
Cwl_66_75 word66_75 gnd C_wl
Rw67_75 word67_75 word66_75 R_wl
Cwl_67_75 word67_75 gnd C_wl
Rw68_75 word68_75 word67_75 R_wl
Cwl_68_75 word68_75 gnd C_wl
Rw69_75 word69_75 word68_75 R_wl
Cwl_69_75 word69_75 gnd C_wl
Rw70_75 word70_75 word69_75 R_wl
Cwl_70_75 word70_75 gnd C_wl
Rw71_75 word71_75 word70_75 R_wl
Cwl_71_75 word71_75 gnd C_wl
Rw72_75 word72_75 word71_75 R_wl
Cwl_72_75 word72_75 gnd C_wl
Rw73_75 word73_75 word72_75 R_wl
Cwl_73_75 word73_75 gnd C_wl
Rw74_75 word74_75 word73_75 R_wl
Cwl_74_75 word74_75 gnd C_wl
Rw75_75 word75_75 word74_75 R_wl
Cwl_75_75 word75_75 gnd C_wl
Rw76_75 word76_75 word75_75 R_wl
Cwl_76_75 word76_75 gnd C_wl
Rw77_75 word77_75 word76_75 R_wl
Cwl_77_75 word77_75 gnd C_wl
Rw78_75 word78_75 word77_75 R_wl
Cwl_78_75 word78_75 gnd C_wl
Rw79_75 word79_75 word78_75 R_wl
Cwl_79_75 word79_75 gnd C_wl
Rw80_75 word80_75 word79_75 R_wl
Cwl_80_75 word80_75 gnd C_wl
Rw81_75 word81_75 word80_75 R_wl
Cwl_81_75 word81_75 gnd C_wl
Rw82_75 word82_75 word81_75 R_wl
Cwl_82_75 word82_75 gnd C_wl
Rw83_75 word83_75 word82_75 R_wl
Cwl_83_75 word83_75 gnd C_wl
Rw84_75 word84_75 word83_75 R_wl
Cwl_84_75 word84_75 gnd C_wl
Rw85_75 word85_75 word84_75 R_wl
Cwl_85_75 word85_75 gnd C_wl
Rw86_75 word86_75 word85_75 R_wl
Cwl_86_75 word86_75 gnd C_wl
Rw87_75 word87_75 word86_75 R_wl
Cwl_87_75 word87_75 gnd C_wl
Rw88_75 word88_75 word87_75 R_wl
Cwl_88_75 word88_75 gnd C_wl
Rw89_75 word89_75 word88_75 R_wl
Cwl_89_75 word89_75 gnd C_wl
Rw90_75 word90_75 word89_75 R_wl
Cwl_90_75 word90_75 gnd C_wl
Rw91_75 word91_75 word90_75 R_wl
Cwl_91_75 word91_75 gnd C_wl
Rw92_75 word92_75 word91_75 R_wl
Cwl_92_75 word92_75 gnd C_wl
Rw93_75 word93_75 word92_75 R_wl
Cwl_93_75 word93_75 gnd C_wl
Rw94_75 word94_75 word93_75 R_wl
Cwl_94_75 word94_75 gnd C_wl
Rw95_75 word95_75 word94_75 R_wl
Cwl_95_75 word95_75 gnd C_wl
Rw96_75 word96_75 word95_75 R_wl
Cwl_96_75 word96_75 gnd C_wl
Rw97_75 word97_75 word96_75 R_wl
Cwl_97_75 word97_75 gnd C_wl
Rw98_75 word98_75 word97_75 R_wl
Cwl_98_75 word98_75 gnd C_wl
Rw99_75 word99_75 word98_75 R_wl
Cwl_99_75 word99_75 gnd C_wl
Vwl_76 word_76 0 0
Rw0_76 word_76 word0_76 R_wl
Cwl_0_76 word0_76 gnd C_wl
Rw1_76 word1_76 word0_76 R_wl
Cwl_1_76 word1_76 gnd C_wl
Rw2_76 word2_76 word1_76 R_wl
Cwl_2_76 word2_76 gnd C_wl
Rw3_76 word3_76 word2_76 R_wl
Cwl_3_76 word3_76 gnd C_wl
Rw4_76 word4_76 word3_76 R_wl
Cwl_4_76 word4_76 gnd C_wl
Rw5_76 word5_76 word4_76 R_wl
Cwl_5_76 word5_76 gnd C_wl
Rw6_76 word6_76 word5_76 R_wl
Cwl_6_76 word6_76 gnd C_wl
Rw7_76 word7_76 word6_76 R_wl
Cwl_7_76 word7_76 gnd C_wl
Rw8_76 word8_76 word7_76 R_wl
Cwl_8_76 word8_76 gnd C_wl
Rw9_76 word9_76 word8_76 R_wl
Cwl_9_76 word9_76 gnd C_wl
Rw10_76 word10_76 word9_76 R_wl
Cwl_10_76 word10_76 gnd C_wl
Rw11_76 word11_76 word10_76 R_wl
Cwl_11_76 word11_76 gnd C_wl
Rw12_76 word12_76 word11_76 R_wl
Cwl_12_76 word12_76 gnd C_wl
Rw13_76 word13_76 word12_76 R_wl
Cwl_13_76 word13_76 gnd C_wl
Rw14_76 word14_76 word13_76 R_wl
Cwl_14_76 word14_76 gnd C_wl
Rw15_76 word15_76 word14_76 R_wl
Cwl_15_76 word15_76 gnd C_wl
Rw16_76 word16_76 word15_76 R_wl
Cwl_16_76 word16_76 gnd C_wl
Rw17_76 word17_76 word16_76 R_wl
Cwl_17_76 word17_76 gnd C_wl
Rw18_76 word18_76 word17_76 R_wl
Cwl_18_76 word18_76 gnd C_wl
Rw19_76 word19_76 word18_76 R_wl
Cwl_19_76 word19_76 gnd C_wl
Rw20_76 word20_76 word19_76 R_wl
Cwl_20_76 word20_76 gnd C_wl
Rw21_76 word21_76 word20_76 R_wl
Cwl_21_76 word21_76 gnd C_wl
Rw22_76 word22_76 word21_76 R_wl
Cwl_22_76 word22_76 gnd C_wl
Rw23_76 word23_76 word22_76 R_wl
Cwl_23_76 word23_76 gnd C_wl
Rw24_76 word24_76 word23_76 R_wl
Cwl_24_76 word24_76 gnd C_wl
Rw25_76 word25_76 word24_76 R_wl
Cwl_25_76 word25_76 gnd C_wl
Rw26_76 word26_76 word25_76 R_wl
Cwl_26_76 word26_76 gnd C_wl
Rw27_76 word27_76 word26_76 R_wl
Cwl_27_76 word27_76 gnd C_wl
Rw28_76 word28_76 word27_76 R_wl
Cwl_28_76 word28_76 gnd C_wl
Rw29_76 word29_76 word28_76 R_wl
Cwl_29_76 word29_76 gnd C_wl
Rw30_76 word30_76 word29_76 R_wl
Cwl_30_76 word30_76 gnd C_wl
Rw31_76 word31_76 word30_76 R_wl
Cwl_31_76 word31_76 gnd C_wl
Rw32_76 word32_76 word31_76 R_wl
Cwl_32_76 word32_76 gnd C_wl
Rw33_76 word33_76 word32_76 R_wl
Cwl_33_76 word33_76 gnd C_wl
Rw34_76 word34_76 word33_76 R_wl
Cwl_34_76 word34_76 gnd C_wl
Rw35_76 word35_76 word34_76 R_wl
Cwl_35_76 word35_76 gnd C_wl
Rw36_76 word36_76 word35_76 R_wl
Cwl_36_76 word36_76 gnd C_wl
Rw37_76 word37_76 word36_76 R_wl
Cwl_37_76 word37_76 gnd C_wl
Rw38_76 word38_76 word37_76 R_wl
Cwl_38_76 word38_76 gnd C_wl
Rw39_76 word39_76 word38_76 R_wl
Cwl_39_76 word39_76 gnd C_wl
Rw40_76 word40_76 word39_76 R_wl
Cwl_40_76 word40_76 gnd C_wl
Rw41_76 word41_76 word40_76 R_wl
Cwl_41_76 word41_76 gnd C_wl
Rw42_76 word42_76 word41_76 R_wl
Cwl_42_76 word42_76 gnd C_wl
Rw43_76 word43_76 word42_76 R_wl
Cwl_43_76 word43_76 gnd C_wl
Rw44_76 word44_76 word43_76 R_wl
Cwl_44_76 word44_76 gnd C_wl
Rw45_76 word45_76 word44_76 R_wl
Cwl_45_76 word45_76 gnd C_wl
Rw46_76 word46_76 word45_76 R_wl
Cwl_46_76 word46_76 gnd C_wl
Rw47_76 word47_76 word46_76 R_wl
Cwl_47_76 word47_76 gnd C_wl
Rw48_76 word48_76 word47_76 R_wl
Cwl_48_76 word48_76 gnd C_wl
Rw49_76 word49_76 word48_76 R_wl
Cwl_49_76 word49_76 gnd C_wl
Rw50_76 word50_76 word49_76 R_wl
Cwl_50_76 word50_76 gnd C_wl
Rw51_76 word51_76 word50_76 R_wl
Cwl_51_76 word51_76 gnd C_wl
Rw52_76 word52_76 word51_76 R_wl
Cwl_52_76 word52_76 gnd C_wl
Rw53_76 word53_76 word52_76 R_wl
Cwl_53_76 word53_76 gnd C_wl
Rw54_76 word54_76 word53_76 R_wl
Cwl_54_76 word54_76 gnd C_wl
Rw55_76 word55_76 word54_76 R_wl
Cwl_55_76 word55_76 gnd C_wl
Rw56_76 word56_76 word55_76 R_wl
Cwl_56_76 word56_76 gnd C_wl
Rw57_76 word57_76 word56_76 R_wl
Cwl_57_76 word57_76 gnd C_wl
Rw58_76 word58_76 word57_76 R_wl
Cwl_58_76 word58_76 gnd C_wl
Rw59_76 word59_76 word58_76 R_wl
Cwl_59_76 word59_76 gnd C_wl
Rw60_76 word60_76 word59_76 R_wl
Cwl_60_76 word60_76 gnd C_wl
Rw61_76 word61_76 word60_76 R_wl
Cwl_61_76 word61_76 gnd C_wl
Rw62_76 word62_76 word61_76 R_wl
Cwl_62_76 word62_76 gnd C_wl
Rw63_76 word63_76 word62_76 R_wl
Cwl_63_76 word63_76 gnd C_wl
Rw64_76 word64_76 word63_76 R_wl
Cwl_64_76 word64_76 gnd C_wl
Rw65_76 word65_76 word64_76 R_wl
Cwl_65_76 word65_76 gnd C_wl
Rw66_76 word66_76 word65_76 R_wl
Cwl_66_76 word66_76 gnd C_wl
Rw67_76 word67_76 word66_76 R_wl
Cwl_67_76 word67_76 gnd C_wl
Rw68_76 word68_76 word67_76 R_wl
Cwl_68_76 word68_76 gnd C_wl
Rw69_76 word69_76 word68_76 R_wl
Cwl_69_76 word69_76 gnd C_wl
Rw70_76 word70_76 word69_76 R_wl
Cwl_70_76 word70_76 gnd C_wl
Rw71_76 word71_76 word70_76 R_wl
Cwl_71_76 word71_76 gnd C_wl
Rw72_76 word72_76 word71_76 R_wl
Cwl_72_76 word72_76 gnd C_wl
Rw73_76 word73_76 word72_76 R_wl
Cwl_73_76 word73_76 gnd C_wl
Rw74_76 word74_76 word73_76 R_wl
Cwl_74_76 word74_76 gnd C_wl
Rw75_76 word75_76 word74_76 R_wl
Cwl_75_76 word75_76 gnd C_wl
Rw76_76 word76_76 word75_76 R_wl
Cwl_76_76 word76_76 gnd C_wl
Rw77_76 word77_76 word76_76 R_wl
Cwl_77_76 word77_76 gnd C_wl
Rw78_76 word78_76 word77_76 R_wl
Cwl_78_76 word78_76 gnd C_wl
Rw79_76 word79_76 word78_76 R_wl
Cwl_79_76 word79_76 gnd C_wl
Rw80_76 word80_76 word79_76 R_wl
Cwl_80_76 word80_76 gnd C_wl
Rw81_76 word81_76 word80_76 R_wl
Cwl_81_76 word81_76 gnd C_wl
Rw82_76 word82_76 word81_76 R_wl
Cwl_82_76 word82_76 gnd C_wl
Rw83_76 word83_76 word82_76 R_wl
Cwl_83_76 word83_76 gnd C_wl
Rw84_76 word84_76 word83_76 R_wl
Cwl_84_76 word84_76 gnd C_wl
Rw85_76 word85_76 word84_76 R_wl
Cwl_85_76 word85_76 gnd C_wl
Rw86_76 word86_76 word85_76 R_wl
Cwl_86_76 word86_76 gnd C_wl
Rw87_76 word87_76 word86_76 R_wl
Cwl_87_76 word87_76 gnd C_wl
Rw88_76 word88_76 word87_76 R_wl
Cwl_88_76 word88_76 gnd C_wl
Rw89_76 word89_76 word88_76 R_wl
Cwl_89_76 word89_76 gnd C_wl
Rw90_76 word90_76 word89_76 R_wl
Cwl_90_76 word90_76 gnd C_wl
Rw91_76 word91_76 word90_76 R_wl
Cwl_91_76 word91_76 gnd C_wl
Rw92_76 word92_76 word91_76 R_wl
Cwl_92_76 word92_76 gnd C_wl
Rw93_76 word93_76 word92_76 R_wl
Cwl_93_76 word93_76 gnd C_wl
Rw94_76 word94_76 word93_76 R_wl
Cwl_94_76 word94_76 gnd C_wl
Rw95_76 word95_76 word94_76 R_wl
Cwl_95_76 word95_76 gnd C_wl
Rw96_76 word96_76 word95_76 R_wl
Cwl_96_76 word96_76 gnd C_wl
Rw97_76 word97_76 word96_76 R_wl
Cwl_97_76 word97_76 gnd C_wl
Rw98_76 word98_76 word97_76 R_wl
Cwl_98_76 word98_76 gnd C_wl
Rw99_76 word99_76 word98_76 R_wl
Cwl_99_76 word99_76 gnd C_wl
Vwl_77 word_77 0 0
Rw0_77 word_77 word0_77 R_wl
Cwl_0_77 word0_77 gnd C_wl
Rw1_77 word1_77 word0_77 R_wl
Cwl_1_77 word1_77 gnd C_wl
Rw2_77 word2_77 word1_77 R_wl
Cwl_2_77 word2_77 gnd C_wl
Rw3_77 word3_77 word2_77 R_wl
Cwl_3_77 word3_77 gnd C_wl
Rw4_77 word4_77 word3_77 R_wl
Cwl_4_77 word4_77 gnd C_wl
Rw5_77 word5_77 word4_77 R_wl
Cwl_5_77 word5_77 gnd C_wl
Rw6_77 word6_77 word5_77 R_wl
Cwl_6_77 word6_77 gnd C_wl
Rw7_77 word7_77 word6_77 R_wl
Cwl_7_77 word7_77 gnd C_wl
Rw8_77 word8_77 word7_77 R_wl
Cwl_8_77 word8_77 gnd C_wl
Rw9_77 word9_77 word8_77 R_wl
Cwl_9_77 word9_77 gnd C_wl
Rw10_77 word10_77 word9_77 R_wl
Cwl_10_77 word10_77 gnd C_wl
Rw11_77 word11_77 word10_77 R_wl
Cwl_11_77 word11_77 gnd C_wl
Rw12_77 word12_77 word11_77 R_wl
Cwl_12_77 word12_77 gnd C_wl
Rw13_77 word13_77 word12_77 R_wl
Cwl_13_77 word13_77 gnd C_wl
Rw14_77 word14_77 word13_77 R_wl
Cwl_14_77 word14_77 gnd C_wl
Rw15_77 word15_77 word14_77 R_wl
Cwl_15_77 word15_77 gnd C_wl
Rw16_77 word16_77 word15_77 R_wl
Cwl_16_77 word16_77 gnd C_wl
Rw17_77 word17_77 word16_77 R_wl
Cwl_17_77 word17_77 gnd C_wl
Rw18_77 word18_77 word17_77 R_wl
Cwl_18_77 word18_77 gnd C_wl
Rw19_77 word19_77 word18_77 R_wl
Cwl_19_77 word19_77 gnd C_wl
Rw20_77 word20_77 word19_77 R_wl
Cwl_20_77 word20_77 gnd C_wl
Rw21_77 word21_77 word20_77 R_wl
Cwl_21_77 word21_77 gnd C_wl
Rw22_77 word22_77 word21_77 R_wl
Cwl_22_77 word22_77 gnd C_wl
Rw23_77 word23_77 word22_77 R_wl
Cwl_23_77 word23_77 gnd C_wl
Rw24_77 word24_77 word23_77 R_wl
Cwl_24_77 word24_77 gnd C_wl
Rw25_77 word25_77 word24_77 R_wl
Cwl_25_77 word25_77 gnd C_wl
Rw26_77 word26_77 word25_77 R_wl
Cwl_26_77 word26_77 gnd C_wl
Rw27_77 word27_77 word26_77 R_wl
Cwl_27_77 word27_77 gnd C_wl
Rw28_77 word28_77 word27_77 R_wl
Cwl_28_77 word28_77 gnd C_wl
Rw29_77 word29_77 word28_77 R_wl
Cwl_29_77 word29_77 gnd C_wl
Rw30_77 word30_77 word29_77 R_wl
Cwl_30_77 word30_77 gnd C_wl
Rw31_77 word31_77 word30_77 R_wl
Cwl_31_77 word31_77 gnd C_wl
Rw32_77 word32_77 word31_77 R_wl
Cwl_32_77 word32_77 gnd C_wl
Rw33_77 word33_77 word32_77 R_wl
Cwl_33_77 word33_77 gnd C_wl
Rw34_77 word34_77 word33_77 R_wl
Cwl_34_77 word34_77 gnd C_wl
Rw35_77 word35_77 word34_77 R_wl
Cwl_35_77 word35_77 gnd C_wl
Rw36_77 word36_77 word35_77 R_wl
Cwl_36_77 word36_77 gnd C_wl
Rw37_77 word37_77 word36_77 R_wl
Cwl_37_77 word37_77 gnd C_wl
Rw38_77 word38_77 word37_77 R_wl
Cwl_38_77 word38_77 gnd C_wl
Rw39_77 word39_77 word38_77 R_wl
Cwl_39_77 word39_77 gnd C_wl
Rw40_77 word40_77 word39_77 R_wl
Cwl_40_77 word40_77 gnd C_wl
Rw41_77 word41_77 word40_77 R_wl
Cwl_41_77 word41_77 gnd C_wl
Rw42_77 word42_77 word41_77 R_wl
Cwl_42_77 word42_77 gnd C_wl
Rw43_77 word43_77 word42_77 R_wl
Cwl_43_77 word43_77 gnd C_wl
Rw44_77 word44_77 word43_77 R_wl
Cwl_44_77 word44_77 gnd C_wl
Rw45_77 word45_77 word44_77 R_wl
Cwl_45_77 word45_77 gnd C_wl
Rw46_77 word46_77 word45_77 R_wl
Cwl_46_77 word46_77 gnd C_wl
Rw47_77 word47_77 word46_77 R_wl
Cwl_47_77 word47_77 gnd C_wl
Rw48_77 word48_77 word47_77 R_wl
Cwl_48_77 word48_77 gnd C_wl
Rw49_77 word49_77 word48_77 R_wl
Cwl_49_77 word49_77 gnd C_wl
Rw50_77 word50_77 word49_77 R_wl
Cwl_50_77 word50_77 gnd C_wl
Rw51_77 word51_77 word50_77 R_wl
Cwl_51_77 word51_77 gnd C_wl
Rw52_77 word52_77 word51_77 R_wl
Cwl_52_77 word52_77 gnd C_wl
Rw53_77 word53_77 word52_77 R_wl
Cwl_53_77 word53_77 gnd C_wl
Rw54_77 word54_77 word53_77 R_wl
Cwl_54_77 word54_77 gnd C_wl
Rw55_77 word55_77 word54_77 R_wl
Cwl_55_77 word55_77 gnd C_wl
Rw56_77 word56_77 word55_77 R_wl
Cwl_56_77 word56_77 gnd C_wl
Rw57_77 word57_77 word56_77 R_wl
Cwl_57_77 word57_77 gnd C_wl
Rw58_77 word58_77 word57_77 R_wl
Cwl_58_77 word58_77 gnd C_wl
Rw59_77 word59_77 word58_77 R_wl
Cwl_59_77 word59_77 gnd C_wl
Rw60_77 word60_77 word59_77 R_wl
Cwl_60_77 word60_77 gnd C_wl
Rw61_77 word61_77 word60_77 R_wl
Cwl_61_77 word61_77 gnd C_wl
Rw62_77 word62_77 word61_77 R_wl
Cwl_62_77 word62_77 gnd C_wl
Rw63_77 word63_77 word62_77 R_wl
Cwl_63_77 word63_77 gnd C_wl
Rw64_77 word64_77 word63_77 R_wl
Cwl_64_77 word64_77 gnd C_wl
Rw65_77 word65_77 word64_77 R_wl
Cwl_65_77 word65_77 gnd C_wl
Rw66_77 word66_77 word65_77 R_wl
Cwl_66_77 word66_77 gnd C_wl
Rw67_77 word67_77 word66_77 R_wl
Cwl_67_77 word67_77 gnd C_wl
Rw68_77 word68_77 word67_77 R_wl
Cwl_68_77 word68_77 gnd C_wl
Rw69_77 word69_77 word68_77 R_wl
Cwl_69_77 word69_77 gnd C_wl
Rw70_77 word70_77 word69_77 R_wl
Cwl_70_77 word70_77 gnd C_wl
Rw71_77 word71_77 word70_77 R_wl
Cwl_71_77 word71_77 gnd C_wl
Rw72_77 word72_77 word71_77 R_wl
Cwl_72_77 word72_77 gnd C_wl
Rw73_77 word73_77 word72_77 R_wl
Cwl_73_77 word73_77 gnd C_wl
Rw74_77 word74_77 word73_77 R_wl
Cwl_74_77 word74_77 gnd C_wl
Rw75_77 word75_77 word74_77 R_wl
Cwl_75_77 word75_77 gnd C_wl
Rw76_77 word76_77 word75_77 R_wl
Cwl_76_77 word76_77 gnd C_wl
Rw77_77 word77_77 word76_77 R_wl
Cwl_77_77 word77_77 gnd C_wl
Rw78_77 word78_77 word77_77 R_wl
Cwl_78_77 word78_77 gnd C_wl
Rw79_77 word79_77 word78_77 R_wl
Cwl_79_77 word79_77 gnd C_wl
Rw80_77 word80_77 word79_77 R_wl
Cwl_80_77 word80_77 gnd C_wl
Rw81_77 word81_77 word80_77 R_wl
Cwl_81_77 word81_77 gnd C_wl
Rw82_77 word82_77 word81_77 R_wl
Cwl_82_77 word82_77 gnd C_wl
Rw83_77 word83_77 word82_77 R_wl
Cwl_83_77 word83_77 gnd C_wl
Rw84_77 word84_77 word83_77 R_wl
Cwl_84_77 word84_77 gnd C_wl
Rw85_77 word85_77 word84_77 R_wl
Cwl_85_77 word85_77 gnd C_wl
Rw86_77 word86_77 word85_77 R_wl
Cwl_86_77 word86_77 gnd C_wl
Rw87_77 word87_77 word86_77 R_wl
Cwl_87_77 word87_77 gnd C_wl
Rw88_77 word88_77 word87_77 R_wl
Cwl_88_77 word88_77 gnd C_wl
Rw89_77 word89_77 word88_77 R_wl
Cwl_89_77 word89_77 gnd C_wl
Rw90_77 word90_77 word89_77 R_wl
Cwl_90_77 word90_77 gnd C_wl
Rw91_77 word91_77 word90_77 R_wl
Cwl_91_77 word91_77 gnd C_wl
Rw92_77 word92_77 word91_77 R_wl
Cwl_92_77 word92_77 gnd C_wl
Rw93_77 word93_77 word92_77 R_wl
Cwl_93_77 word93_77 gnd C_wl
Rw94_77 word94_77 word93_77 R_wl
Cwl_94_77 word94_77 gnd C_wl
Rw95_77 word95_77 word94_77 R_wl
Cwl_95_77 word95_77 gnd C_wl
Rw96_77 word96_77 word95_77 R_wl
Cwl_96_77 word96_77 gnd C_wl
Rw97_77 word97_77 word96_77 R_wl
Cwl_97_77 word97_77 gnd C_wl
Rw98_77 word98_77 word97_77 R_wl
Cwl_98_77 word98_77 gnd C_wl
Rw99_77 word99_77 word98_77 R_wl
Cwl_99_77 word99_77 gnd C_wl
Vwl_78 word_78 0 0
Rw0_78 word_78 word0_78 R_wl
Cwl_0_78 word0_78 gnd C_wl
Rw1_78 word1_78 word0_78 R_wl
Cwl_1_78 word1_78 gnd C_wl
Rw2_78 word2_78 word1_78 R_wl
Cwl_2_78 word2_78 gnd C_wl
Rw3_78 word3_78 word2_78 R_wl
Cwl_3_78 word3_78 gnd C_wl
Rw4_78 word4_78 word3_78 R_wl
Cwl_4_78 word4_78 gnd C_wl
Rw5_78 word5_78 word4_78 R_wl
Cwl_5_78 word5_78 gnd C_wl
Rw6_78 word6_78 word5_78 R_wl
Cwl_6_78 word6_78 gnd C_wl
Rw7_78 word7_78 word6_78 R_wl
Cwl_7_78 word7_78 gnd C_wl
Rw8_78 word8_78 word7_78 R_wl
Cwl_8_78 word8_78 gnd C_wl
Rw9_78 word9_78 word8_78 R_wl
Cwl_9_78 word9_78 gnd C_wl
Rw10_78 word10_78 word9_78 R_wl
Cwl_10_78 word10_78 gnd C_wl
Rw11_78 word11_78 word10_78 R_wl
Cwl_11_78 word11_78 gnd C_wl
Rw12_78 word12_78 word11_78 R_wl
Cwl_12_78 word12_78 gnd C_wl
Rw13_78 word13_78 word12_78 R_wl
Cwl_13_78 word13_78 gnd C_wl
Rw14_78 word14_78 word13_78 R_wl
Cwl_14_78 word14_78 gnd C_wl
Rw15_78 word15_78 word14_78 R_wl
Cwl_15_78 word15_78 gnd C_wl
Rw16_78 word16_78 word15_78 R_wl
Cwl_16_78 word16_78 gnd C_wl
Rw17_78 word17_78 word16_78 R_wl
Cwl_17_78 word17_78 gnd C_wl
Rw18_78 word18_78 word17_78 R_wl
Cwl_18_78 word18_78 gnd C_wl
Rw19_78 word19_78 word18_78 R_wl
Cwl_19_78 word19_78 gnd C_wl
Rw20_78 word20_78 word19_78 R_wl
Cwl_20_78 word20_78 gnd C_wl
Rw21_78 word21_78 word20_78 R_wl
Cwl_21_78 word21_78 gnd C_wl
Rw22_78 word22_78 word21_78 R_wl
Cwl_22_78 word22_78 gnd C_wl
Rw23_78 word23_78 word22_78 R_wl
Cwl_23_78 word23_78 gnd C_wl
Rw24_78 word24_78 word23_78 R_wl
Cwl_24_78 word24_78 gnd C_wl
Rw25_78 word25_78 word24_78 R_wl
Cwl_25_78 word25_78 gnd C_wl
Rw26_78 word26_78 word25_78 R_wl
Cwl_26_78 word26_78 gnd C_wl
Rw27_78 word27_78 word26_78 R_wl
Cwl_27_78 word27_78 gnd C_wl
Rw28_78 word28_78 word27_78 R_wl
Cwl_28_78 word28_78 gnd C_wl
Rw29_78 word29_78 word28_78 R_wl
Cwl_29_78 word29_78 gnd C_wl
Rw30_78 word30_78 word29_78 R_wl
Cwl_30_78 word30_78 gnd C_wl
Rw31_78 word31_78 word30_78 R_wl
Cwl_31_78 word31_78 gnd C_wl
Rw32_78 word32_78 word31_78 R_wl
Cwl_32_78 word32_78 gnd C_wl
Rw33_78 word33_78 word32_78 R_wl
Cwl_33_78 word33_78 gnd C_wl
Rw34_78 word34_78 word33_78 R_wl
Cwl_34_78 word34_78 gnd C_wl
Rw35_78 word35_78 word34_78 R_wl
Cwl_35_78 word35_78 gnd C_wl
Rw36_78 word36_78 word35_78 R_wl
Cwl_36_78 word36_78 gnd C_wl
Rw37_78 word37_78 word36_78 R_wl
Cwl_37_78 word37_78 gnd C_wl
Rw38_78 word38_78 word37_78 R_wl
Cwl_38_78 word38_78 gnd C_wl
Rw39_78 word39_78 word38_78 R_wl
Cwl_39_78 word39_78 gnd C_wl
Rw40_78 word40_78 word39_78 R_wl
Cwl_40_78 word40_78 gnd C_wl
Rw41_78 word41_78 word40_78 R_wl
Cwl_41_78 word41_78 gnd C_wl
Rw42_78 word42_78 word41_78 R_wl
Cwl_42_78 word42_78 gnd C_wl
Rw43_78 word43_78 word42_78 R_wl
Cwl_43_78 word43_78 gnd C_wl
Rw44_78 word44_78 word43_78 R_wl
Cwl_44_78 word44_78 gnd C_wl
Rw45_78 word45_78 word44_78 R_wl
Cwl_45_78 word45_78 gnd C_wl
Rw46_78 word46_78 word45_78 R_wl
Cwl_46_78 word46_78 gnd C_wl
Rw47_78 word47_78 word46_78 R_wl
Cwl_47_78 word47_78 gnd C_wl
Rw48_78 word48_78 word47_78 R_wl
Cwl_48_78 word48_78 gnd C_wl
Rw49_78 word49_78 word48_78 R_wl
Cwl_49_78 word49_78 gnd C_wl
Rw50_78 word50_78 word49_78 R_wl
Cwl_50_78 word50_78 gnd C_wl
Rw51_78 word51_78 word50_78 R_wl
Cwl_51_78 word51_78 gnd C_wl
Rw52_78 word52_78 word51_78 R_wl
Cwl_52_78 word52_78 gnd C_wl
Rw53_78 word53_78 word52_78 R_wl
Cwl_53_78 word53_78 gnd C_wl
Rw54_78 word54_78 word53_78 R_wl
Cwl_54_78 word54_78 gnd C_wl
Rw55_78 word55_78 word54_78 R_wl
Cwl_55_78 word55_78 gnd C_wl
Rw56_78 word56_78 word55_78 R_wl
Cwl_56_78 word56_78 gnd C_wl
Rw57_78 word57_78 word56_78 R_wl
Cwl_57_78 word57_78 gnd C_wl
Rw58_78 word58_78 word57_78 R_wl
Cwl_58_78 word58_78 gnd C_wl
Rw59_78 word59_78 word58_78 R_wl
Cwl_59_78 word59_78 gnd C_wl
Rw60_78 word60_78 word59_78 R_wl
Cwl_60_78 word60_78 gnd C_wl
Rw61_78 word61_78 word60_78 R_wl
Cwl_61_78 word61_78 gnd C_wl
Rw62_78 word62_78 word61_78 R_wl
Cwl_62_78 word62_78 gnd C_wl
Rw63_78 word63_78 word62_78 R_wl
Cwl_63_78 word63_78 gnd C_wl
Rw64_78 word64_78 word63_78 R_wl
Cwl_64_78 word64_78 gnd C_wl
Rw65_78 word65_78 word64_78 R_wl
Cwl_65_78 word65_78 gnd C_wl
Rw66_78 word66_78 word65_78 R_wl
Cwl_66_78 word66_78 gnd C_wl
Rw67_78 word67_78 word66_78 R_wl
Cwl_67_78 word67_78 gnd C_wl
Rw68_78 word68_78 word67_78 R_wl
Cwl_68_78 word68_78 gnd C_wl
Rw69_78 word69_78 word68_78 R_wl
Cwl_69_78 word69_78 gnd C_wl
Rw70_78 word70_78 word69_78 R_wl
Cwl_70_78 word70_78 gnd C_wl
Rw71_78 word71_78 word70_78 R_wl
Cwl_71_78 word71_78 gnd C_wl
Rw72_78 word72_78 word71_78 R_wl
Cwl_72_78 word72_78 gnd C_wl
Rw73_78 word73_78 word72_78 R_wl
Cwl_73_78 word73_78 gnd C_wl
Rw74_78 word74_78 word73_78 R_wl
Cwl_74_78 word74_78 gnd C_wl
Rw75_78 word75_78 word74_78 R_wl
Cwl_75_78 word75_78 gnd C_wl
Rw76_78 word76_78 word75_78 R_wl
Cwl_76_78 word76_78 gnd C_wl
Rw77_78 word77_78 word76_78 R_wl
Cwl_77_78 word77_78 gnd C_wl
Rw78_78 word78_78 word77_78 R_wl
Cwl_78_78 word78_78 gnd C_wl
Rw79_78 word79_78 word78_78 R_wl
Cwl_79_78 word79_78 gnd C_wl
Rw80_78 word80_78 word79_78 R_wl
Cwl_80_78 word80_78 gnd C_wl
Rw81_78 word81_78 word80_78 R_wl
Cwl_81_78 word81_78 gnd C_wl
Rw82_78 word82_78 word81_78 R_wl
Cwl_82_78 word82_78 gnd C_wl
Rw83_78 word83_78 word82_78 R_wl
Cwl_83_78 word83_78 gnd C_wl
Rw84_78 word84_78 word83_78 R_wl
Cwl_84_78 word84_78 gnd C_wl
Rw85_78 word85_78 word84_78 R_wl
Cwl_85_78 word85_78 gnd C_wl
Rw86_78 word86_78 word85_78 R_wl
Cwl_86_78 word86_78 gnd C_wl
Rw87_78 word87_78 word86_78 R_wl
Cwl_87_78 word87_78 gnd C_wl
Rw88_78 word88_78 word87_78 R_wl
Cwl_88_78 word88_78 gnd C_wl
Rw89_78 word89_78 word88_78 R_wl
Cwl_89_78 word89_78 gnd C_wl
Rw90_78 word90_78 word89_78 R_wl
Cwl_90_78 word90_78 gnd C_wl
Rw91_78 word91_78 word90_78 R_wl
Cwl_91_78 word91_78 gnd C_wl
Rw92_78 word92_78 word91_78 R_wl
Cwl_92_78 word92_78 gnd C_wl
Rw93_78 word93_78 word92_78 R_wl
Cwl_93_78 word93_78 gnd C_wl
Rw94_78 word94_78 word93_78 R_wl
Cwl_94_78 word94_78 gnd C_wl
Rw95_78 word95_78 word94_78 R_wl
Cwl_95_78 word95_78 gnd C_wl
Rw96_78 word96_78 word95_78 R_wl
Cwl_96_78 word96_78 gnd C_wl
Rw97_78 word97_78 word96_78 R_wl
Cwl_97_78 word97_78 gnd C_wl
Rw98_78 word98_78 word97_78 R_wl
Cwl_98_78 word98_78 gnd C_wl
Rw99_78 word99_78 word98_78 R_wl
Cwl_99_78 word99_78 gnd C_wl
Vwl_79 word_79 0 0
Rw0_79 word_79 word0_79 R_wl
Cwl_0_79 word0_79 gnd C_wl
Rw1_79 word1_79 word0_79 R_wl
Cwl_1_79 word1_79 gnd C_wl
Rw2_79 word2_79 word1_79 R_wl
Cwl_2_79 word2_79 gnd C_wl
Rw3_79 word3_79 word2_79 R_wl
Cwl_3_79 word3_79 gnd C_wl
Rw4_79 word4_79 word3_79 R_wl
Cwl_4_79 word4_79 gnd C_wl
Rw5_79 word5_79 word4_79 R_wl
Cwl_5_79 word5_79 gnd C_wl
Rw6_79 word6_79 word5_79 R_wl
Cwl_6_79 word6_79 gnd C_wl
Rw7_79 word7_79 word6_79 R_wl
Cwl_7_79 word7_79 gnd C_wl
Rw8_79 word8_79 word7_79 R_wl
Cwl_8_79 word8_79 gnd C_wl
Rw9_79 word9_79 word8_79 R_wl
Cwl_9_79 word9_79 gnd C_wl
Rw10_79 word10_79 word9_79 R_wl
Cwl_10_79 word10_79 gnd C_wl
Rw11_79 word11_79 word10_79 R_wl
Cwl_11_79 word11_79 gnd C_wl
Rw12_79 word12_79 word11_79 R_wl
Cwl_12_79 word12_79 gnd C_wl
Rw13_79 word13_79 word12_79 R_wl
Cwl_13_79 word13_79 gnd C_wl
Rw14_79 word14_79 word13_79 R_wl
Cwl_14_79 word14_79 gnd C_wl
Rw15_79 word15_79 word14_79 R_wl
Cwl_15_79 word15_79 gnd C_wl
Rw16_79 word16_79 word15_79 R_wl
Cwl_16_79 word16_79 gnd C_wl
Rw17_79 word17_79 word16_79 R_wl
Cwl_17_79 word17_79 gnd C_wl
Rw18_79 word18_79 word17_79 R_wl
Cwl_18_79 word18_79 gnd C_wl
Rw19_79 word19_79 word18_79 R_wl
Cwl_19_79 word19_79 gnd C_wl
Rw20_79 word20_79 word19_79 R_wl
Cwl_20_79 word20_79 gnd C_wl
Rw21_79 word21_79 word20_79 R_wl
Cwl_21_79 word21_79 gnd C_wl
Rw22_79 word22_79 word21_79 R_wl
Cwl_22_79 word22_79 gnd C_wl
Rw23_79 word23_79 word22_79 R_wl
Cwl_23_79 word23_79 gnd C_wl
Rw24_79 word24_79 word23_79 R_wl
Cwl_24_79 word24_79 gnd C_wl
Rw25_79 word25_79 word24_79 R_wl
Cwl_25_79 word25_79 gnd C_wl
Rw26_79 word26_79 word25_79 R_wl
Cwl_26_79 word26_79 gnd C_wl
Rw27_79 word27_79 word26_79 R_wl
Cwl_27_79 word27_79 gnd C_wl
Rw28_79 word28_79 word27_79 R_wl
Cwl_28_79 word28_79 gnd C_wl
Rw29_79 word29_79 word28_79 R_wl
Cwl_29_79 word29_79 gnd C_wl
Rw30_79 word30_79 word29_79 R_wl
Cwl_30_79 word30_79 gnd C_wl
Rw31_79 word31_79 word30_79 R_wl
Cwl_31_79 word31_79 gnd C_wl
Rw32_79 word32_79 word31_79 R_wl
Cwl_32_79 word32_79 gnd C_wl
Rw33_79 word33_79 word32_79 R_wl
Cwl_33_79 word33_79 gnd C_wl
Rw34_79 word34_79 word33_79 R_wl
Cwl_34_79 word34_79 gnd C_wl
Rw35_79 word35_79 word34_79 R_wl
Cwl_35_79 word35_79 gnd C_wl
Rw36_79 word36_79 word35_79 R_wl
Cwl_36_79 word36_79 gnd C_wl
Rw37_79 word37_79 word36_79 R_wl
Cwl_37_79 word37_79 gnd C_wl
Rw38_79 word38_79 word37_79 R_wl
Cwl_38_79 word38_79 gnd C_wl
Rw39_79 word39_79 word38_79 R_wl
Cwl_39_79 word39_79 gnd C_wl
Rw40_79 word40_79 word39_79 R_wl
Cwl_40_79 word40_79 gnd C_wl
Rw41_79 word41_79 word40_79 R_wl
Cwl_41_79 word41_79 gnd C_wl
Rw42_79 word42_79 word41_79 R_wl
Cwl_42_79 word42_79 gnd C_wl
Rw43_79 word43_79 word42_79 R_wl
Cwl_43_79 word43_79 gnd C_wl
Rw44_79 word44_79 word43_79 R_wl
Cwl_44_79 word44_79 gnd C_wl
Rw45_79 word45_79 word44_79 R_wl
Cwl_45_79 word45_79 gnd C_wl
Rw46_79 word46_79 word45_79 R_wl
Cwl_46_79 word46_79 gnd C_wl
Rw47_79 word47_79 word46_79 R_wl
Cwl_47_79 word47_79 gnd C_wl
Rw48_79 word48_79 word47_79 R_wl
Cwl_48_79 word48_79 gnd C_wl
Rw49_79 word49_79 word48_79 R_wl
Cwl_49_79 word49_79 gnd C_wl
Rw50_79 word50_79 word49_79 R_wl
Cwl_50_79 word50_79 gnd C_wl
Rw51_79 word51_79 word50_79 R_wl
Cwl_51_79 word51_79 gnd C_wl
Rw52_79 word52_79 word51_79 R_wl
Cwl_52_79 word52_79 gnd C_wl
Rw53_79 word53_79 word52_79 R_wl
Cwl_53_79 word53_79 gnd C_wl
Rw54_79 word54_79 word53_79 R_wl
Cwl_54_79 word54_79 gnd C_wl
Rw55_79 word55_79 word54_79 R_wl
Cwl_55_79 word55_79 gnd C_wl
Rw56_79 word56_79 word55_79 R_wl
Cwl_56_79 word56_79 gnd C_wl
Rw57_79 word57_79 word56_79 R_wl
Cwl_57_79 word57_79 gnd C_wl
Rw58_79 word58_79 word57_79 R_wl
Cwl_58_79 word58_79 gnd C_wl
Rw59_79 word59_79 word58_79 R_wl
Cwl_59_79 word59_79 gnd C_wl
Rw60_79 word60_79 word59_79 R_wl
Cwl_60_79 word60_79 gnd C_wl
Rw61_79 word61_79 word60_79 R_wl
Cwl_61_79 word61_79 gnd C_wl
Rw62_79 word62_79 word61_79 R_wl
Cwl_62_79 word62_79 gnd C_wl
Rw63_79 word63_79 word62_79 R_wl
Cwl_63_79 word63_79 gnd C_wl
Rw64_79 word64_79 word63_79 R_wl
Cwl_64_79 word64_79 gnd C_wl
Rw65_79 word65_79 word64_79 R_wl
Cwl_65_79 word65_79 gnd C_wl
Rw66_79 word66_79 word65_79 R_wl
Cwl_66_79 word66_79 gnd C_wl
Rw67_79 word67_79 word66_79 R_wl
Cwl_67_79 word67_79 gnd C_wl
Rw68_79 word68_79 word67_79 R_wl
Cwl_68_79 word68_79 gnd C_wl
Rw69_79 word69_79 word68_79 R_wl
Cwl_69_79 word69_79 gnd C_wl
Rw70_79 word70_79 word69_79 R_wl
Cwl_70_79 word70_79 gnd C_wl
Rw71_79 word71_79 word70_79 R_wl
Cwl_71_79 word71_79 gnd C_wl
Rw72_79 word72_79 word71_79 R_wl
Cwl_72_79 word72_79 gnd C_wl
Rw73_79 word73_79 word72_79 R_wl
Cwl_73_79 word73_79 gnd C_wl
Rw74_79 word74_79 word73_79 R_wl
Cwl_74_79 word74_79 gnd C_wl
Rw75_79 word75_79 word74_79 R_wl
Cwl_75_79 word75_79 gnd C_wl
Rw76_79 word76_79 word75_79 R_wl
Cwl_76_79 word76_79 gnd C_wl
Rw77_79 word77_79 word76_79 R_wl
Cwl_77_79 word77_79 gnd C_wl
Rw78_79 word78_79 word77_79 R_wl
Cwl_78_79 word78_79 gnd C_wl
Rw79_79 word79_79 word78_79 R_wl
Cwl_79_79 word79_79 gnd C_wl
Rw80_79 word80_79 word79_79 R_wl
Cwl_80_79 word80_79 gnd C_wl
Rw81_79 word81_79 word80_79 R_wl
Cwl_81_79 word81_79 gnd C_wl
Rw82_79 word82_79 word81_79 R_wl
Cwl_82_79 word82_79 gnd C_wl
Rw83_79 word83_79 word82_79 R_wl
Cwl_83_79 word83_79 gnd C_wl
Rw84_79 word84_79 word83_79 R_wl
Cwl_84_79 word84_79 gnd C_wl
Rw85_79 word85_79 word84_79 R_wl
Cwl_85_79 word85_79 gnd C_wl
Rw86_79 word86_79 word85_79 R_wl
Cwl_86_79 word86_79 gnd C_wl
Rw87_79 word87_79 word86_79 R_wl
Cwl_87_79 word87_79 gnd C_wl
Rw88_79 word88_79 word87_79 R_wl
Cwl_88_79 word88_79 gnd C_wl
Rw89_79 word89_79 word88_79 R_wl
Cwl_89_79 word89_79 gnd C_wl
Rw90_79 word90_79 word89_79 R_wl
Cwl_90_79 word90_79 gnd C_wl
Rw91_79 word91_79 word90_79 R_wl
Cwl_91_79 word91_79 gnd C_wl
Rw92_79 word92_79 word91_79 R_wl
Cwl_92_79 word92_79 gnd C_wl
Rw93_79 word93_79 word92_79 R_wl
Cwl_93_79 word93_79 gnd C_wl
Rw94_79 word94_79 word93_79 R_wl
Cwl_94_79 word94_79 gnd C_wl
Rw95_79 word95_79 word94_79 R_wl
Cwl_95_79 word95_79 gnd C_wl
Rw96_79 word96_79 word95_79 R_wl
Cwl_96_79 word96_79 gnd C_wl
Rw97_79 word97_79 word96_79 R_wl
Cwl_97_79 word97_79 gnd C_wl
Rw98_79 word98_79 word97_79 R_wl
Cwl_98_79 word98_79 gnd C_wl
Rw99_79 word99_79 word98_79 R_wl
Cwl_99_79 word99_79 gnd C_wl
Vwl_80 word_80 0 0
Rw0_80 word_80 word0_80 R_wl
Cwl_0_80 word0_80 gnd C_wl
Rw1_80 word1_80 word0_80 R_wl
Cwl_1_80 word1_80 gnd C_wl
Rw2_80 word2_80 word1_80 R_wl
Cwl_2_80 word2_80 gnd C_wl
Rw3_80 word3_80 word2_80 R_wl
Cwl_3_80 word3_80 gnd C_wl
Rw4_80 word4_80 word3_80 R_wl
Cwl_4_80 word4_80 gnd C_wl
Rw5_80 word5_80 word4_80 R_wl
Cwl_5_80 word5_80 gnd C_wl
Rw6_80 word6_80 word5_80 R_wl
Cwl_6_80 word6_80 gnd C_wl
Rw7_80 word7_80 word6_80 R_wl
Cwl_7_80 word7_80 gnd C_wl
Rw8_80 word8_80 word7_80 R_wl
Cwl_8_80 word8_80 gnd C_wl
Rw9_80 word9_80 word8_80 R_wl
Cwl_9_80 word9_80 gnd C_wl
Rw10_80 word10_80 word9_80 R_wl
Cwl_10_80 word10_80 gnd C_wl
Rw11_80 word11_80 word10_80 R_wl
Cwl_11_80 word11_80 gnd C_wl
Rw12_80 word12_80 word11_80 R_wl
Cwl_12_80 word12_80 gnd C_wl
Rw13_80 word13_80 word12_80 R_wl
Cwl_13_80 word13_80 gnd C_wl
Rw14_80 word14_80 word13_80 R_wl
Cwl_14_80 word14_80 gnd C_wl
Rw15_80 word15_80 word14_80 R_wl
Cwl_15_80 word15_80 gnd C_wl
Rw16_80 word16_80 word15_80 R_wl
Cwl_16_80 word16_80 gnd C_wl
Rw17_80 word17_80 word16_80 R_wl
Cwl_17_80 word17_80 gnd C_wl
Rw18_80 word18_80 word17_80 R_wl
Cwl_18_80 word18_80 gnd C_wl
Rw19_80 word19_80 word18_80 R_wl
Cwl_19_80 word19_80 gnd C_wl
Rw20_80 word20_80 word19_80 R_wl
Cwl_20_80 word20_80 gnd C_wl
Rw21_80 word21_80 word20_80 R_wl
Cwl_21_80 word21_80 gnd C_wl
Rw22_80 word22_80 word21_80 R_wl
Cwl_22_80 word22_80 gnd C_wl
Rw23_80 word23_80 word22_80 R_wl
Cwl_23_80 word23_80 gnd C_wl
Rw24_80 word24_80 word23_80 R_wl
Cwl_24_80 word24_80 gnd C_wl
Rw25_80 word25_80 word24_80 R_wl
Cwl_25_80 word25_80 gnd C_wl
Rw26_80 word26_80 word25_80 R_wl
Cwl_26_80 word26_80 gnd C_wl
Rw27_80 word27_80 word26_80 R_wl
Cwl_27_80 word27_80 gnd C_wl
Rw28_80 word28_80 word27_80 R_wl
Cwl_28_80 word28_80 gnd C_wl
Rw29_80 word29_80 word28_80 R_wl
Cwl_29_80 word29_80 gnd C_wl
Rw30_80 word30_80 word29_80 R_wl
Cwl_30_80 word30_80 gnd C_wl
Rw31_80 word31_80 word30_80 R_wl
Cwl_31_80 word31_80 gnd C_wl
Rw32_80 word32_80 word31_80 R_wl
Cwl_32_80 word32_80 gnd C_wl
Rw33_80 word33_80 word32_80 R_wl
Cwl_33_80 word33_80 gnd C_wl
Rw34_80 word34_80 word33_80 R_wl
Cwl_34_80 word34_80 gnd C_wl
Rw35_80 word35_80 word34_80 R_wl
Cwl_35_80 word35_80 gnd C_wl
Rw36_80 word36_80 word35_80 R_wl
Cwl_36_80 word36_80 gnd C_wl
Rw37_80 word37_80 word36_80 R_wl
Cwl_37_80 word37_80 gnd C_wl
Rw38_80 word38_80 word37_80 R_wl
Cwl_38_80 word38_80 gnd C_wl
Rw39_80 word39_80 word38_80 R_wl
Cwl_39_80 word39_80 gnd C_wl
Rw40_80 word40_80 word39_80 R_wl
Cwl_40_80 word40_80 gnd C_wl
Rw41_80 word41_80 word40_80 R_wl
Cwl_41_80 word41_80 gnd C_wl
Rw42_80 word42_80 word41_80 R_wl
Cwl_42_80 word42_80 gnd C_wl
Rw43_80 word43_80 word42_80 R_wl
Cwl_43_80 word43_80 gnd C_wl
Rw44_80 word44_80 word43_80 R_wl
Cwl_44_80 word44_80 gnd C_wl
Rw45_80 word45_80 word44_80 R_wl
Cwl_45_80 word45_80 gnd C_wl
Rw46_80 word46_80 word45_80 R_wl
Cwl_46_80 word46_80 gnd C_wl
Rw47_80 word47_80 word46_80 R_wl
Cwl_47_80 word47_80 gnd C_wl
Rw48_80 word48_80 word47_80 R_wl
Cwl_48_80 word48_80 gnd C_wl
Rw49_80 word49_80 word48_80 R_wl
Cwl_49_80 word49_80 gnd C_wl
Rw50_80 word50_80 word49_80 R_wl
Cwl_50_80 word50_80 gnd C_wl
Rw51_80 word51_80 word50_80 R_wl
Cwl_51_80 word51_80 gnd C_wl
Rw52_80 word52_80 word51_80 R_wl
Cwl_52_80 word52_80 gnd C_wl
Rw53_80 word53_80 word52_80 R_wl
Cwl_53_80 word53_80 gnd C_wl
Rw54_80 word54_80 word53_80 R_wl
Cwl_54_80 word54_80 gnd C_wl
Rw55_80 word55_80 word54_80 R_wl
Cwl_55_80 word55_80 gnd C_wl
Rw56_80 word56_80 word55_80 R_wl
Cwl_56_80 word56_80 gnd C_wl
Rw57_80 word57_80 word56_80 R_wl
Cwl_57_80 word57_80 gnd C_wl
Rw58_80 word58_80 word57_80 R_wl
Cwl_58_80 word58_80 gnd C_wl
Rw59_80 word59_80 word58_80 R_wl
Cwl_59_80 word59_80 gnd C_wl
Rw60_80 word60_80 word59_80 R_wl
Cwl_60_80 word60_80 gnd C_wl
Rw61_80 word61_80 word60_80 R_wl
Cwl_61_80 word61_80 gnd C_wl
Rw62_80 word62_80 word61_80 R_wl
Cwl_62_80 word62_80 gnd C_wl
Rw63_80 word63_80 word62_80 R_wl
Cwl_63_80 word63_80 gnd C_wl
Rw64_80 word64_80 word63_80 R_wl
Cwl_64_80 word64_80 gnd C_wl
Rw65_80 word65_80 word64_80 R_wl
Cwl_65_80 word65_80 gnd C_wl
Rw66_80 word66_80 word65_80 R_wl
Cwl_66_80 word66_80 gnd C_wl
Rw67_80 word67_80 word66_80 R_wl
Cwl_67_80 word67_80 gnd C_wl
Rw68_80 word68_80 word67_80 R_wl
Cwl_68_80 word68_80 gnd C_wl
Rw69_80 word69_80 word68_80 R_wl
Cwl_69_80 word69_80 gnd C_wl
Rw70_80 word70_80 word69_80 R_wl
Cwl_70_80 word70_80 gnd C_wl
Rw71_80 word71_80 word70_80 R_wl
Cwl_71_80 word71_80 gnd C_wl
Rw72_80 word72_80 word71_80 R_wl
Cwl_72_80 word72_80 gnd C_wl
Rw73_80 word73_80 word72_80 R_wl
Cwl_73_80 word73_80 gnd C_wl
Rw74_80 word74_80 word73_80 R_wl
Cwl_74_80 word74_80 gnd C_wl
Rw75_80 word75_80 word74_80 R_wl
Cwl_75_80 word75_80 gnd C_wl
Rw76_80 word76_80 word75_80 R_wl
Cwl_76_80 word76_80 gnd C_wl
Rw77_80 word77_80 word76_80 R_wl
Cwl_77_80 word77_80 gnd C_wl
Rw78_80 word78_80 word77_80 R_wl
Cwl_78_80 word78_80 gnd C_wl
Rw79_80 word79_80 word78_80 R_wl
Cwl_79_80 word79_80 gnd C_wl
Rw80_80 word80_80 word79_80 R_wl
Cwl_80_80 word80_80 gnd C_wl
Rw81_80 word81_80 word80_80 R_wl
Cwl_81_80 word81_80 gnd C_wl
Rw82_80 word82_80 word81_80 R_wl
Cwl_82_80 word82_80 gnd C_wl
Rw83_80 word83_80 word82_80 R_wl
Cwl_83_80 word83_80 gnd C_wl
Rw84_80 word84_80 word83_80 R_wl
Cwl_84_80 word84_80 gnd C_wl
Rw85_80 word85_80 word84_80 R_wl
Cwl_85_80 word85_80 gnd C_wl
Rw86_80 word86_80 word85_80 R_wl
Cwl_86_80 word86_80 gnd C_wl
Rw87_80 word87_80 word86_80 R_wl
Cwl_87_80 word87_80 gnd C_wl
Rw88_80 word88_80 word87_80 R_wl
Cwl_88_80 word88_80 gnd C_wl
Rw89_80 word89_80 word88_80 R_wl
Cwl_89_80 word89_80 gnd C_wl
Rw90_80 word90_80 word89_80 R_wl
Cwl_90_80 word90_80 gnd C_wl
Rw91_80 word91_80 word90_80 R_wl
Cwl_91_80 word91_80 gnd C_wl
Rw92_80 word92_80 word91_80 R_wl
Cwl_92_80 word92_80 gnd C_wl
Rw93_80 word93_80 word92_80 R_wl
Cwl_93_80 word93_80 gnd C_wl
Rw94_80 word94_80 word93_80 R_wl
Cwl_94_80 word94_80 gnd C_wl
Rw95_80 word95_80 word94_80 R_wl
Cwl_95_80 word95_80 gnd C_wl
Rw96_80 word96_80 word95_80 R_wl
Cwl_96_80 word96_80 gnd C_wl
Rw97_80 word97_80 word96_80 R_wl
Cwl_97_80 word97_80 gnd C_wl
Rw98_80 word98_80 word97_80 R_wl
Cwl_98_80 word98_80 gnd C_wl
Rw99_80 word99_80 word98_80 R_wl
Cwl_99_80 word99_80 gnd C_wl
Vwl_81 word_81 0 0
Rw0_81 word_81 word0_81 R_wl
Cwl_0_81 word0_81 gnd C_wl
Rw1_81 word1_81 word0_81 R_wl
Cwl_1_81 word1_81 gnd C_wl
Rw2_81 word2_81 word1_81 R_wl
Cwl_2_81 word2_81 gnd C_wl
Rw3_81 word3_81 word2_81 R_wl
Cwl_3_81 word3_81 gnd C_wl
Rw4_81 word4_81 word3_81 R_wl
Cwl_4_81 word4_81 gnd C_wl
Rw5_81 word5_81 word4_81 R_wl
Cwl_5_81 word5_81 gnd C_wl
Rw6_81 word6_81 word5_81 R_wl
Cwl_6_81 word6_81 gnd C_wl
Rw7_81 word7_81 word6_81 R_wl
Cwl_7_81 word7_81 gnd C_wl
Rw8_81 word8_81 word7_81 R_wl
Cwl_8_81 word8_81 gnd C_wl
Rw9_81 word9_81 word8_81 R_wl
Cwl_9_81 word9_81 gnd C_wl
Rw10_81 word10_81 word9_81 R_wl
Cwl_10_81 word10_81 gnd C_wl
Rw11_81 word11_81 word10_81 R_wl
Cwl_11_81 word11_81 gnd C_wl
Rw12_81 word12_81 word11_81 R_wl
Cwl_12_81 word12_81 gnd C_wl
Rw13_81 word13_81 word12_81 R_wl
Cwl_13_81 word13_81 gnd C_wl
Rw14_81 word14_81 word13_81 R_wl
Cwl_14_81 word14_81 gnd C_wl
Rw15_81 word15_81 word14_81 R_wl
Cwl_15_81 word15_81 gnd C_wl
Rw16_81 word16_81 word15_81 R_wl
Cwl_16_81 word16_81 gnd C_wl
Rw17_81 word17_81 word16_81 R_wl
Cwl_17_81 word17_81 gnd C_wl
Rw18_81 word18_81 word17_81 R_wl
Cwl_18_81 word18_81 gnd C_wl
Rw19_81 word19_81 word18_81 R_wl
Cwl_19_81 word19_81 gnd C_wl
Rw20_81 word20_81 word19_81 R_wl
Cwl_20_81 word20_81 gnd C_wl
Rw21_81 word21_81 word20_81 R_wl
Cwl_21_81 word21_81 gnd C_wl
Rw22_81 word22_81 word21_81 R_wl
Cwl_22_81 word22_81 gnd C_wl
Rw23_81 word23_81 word22_81 R_wl
Cwl_23_81 word23_81 gnd C_wl
Rw24_81 word24_81 word23_81 R_wl
Cwl_24_81 word24_81 gnd C_wl
Rw25_81 word25_81 word24_81 R_wl
Cwl_25_81 word25_81 gnd C_wl
Rw26_81 word26_81 word25_81 R_wl
Cwl_26_81 word26_81 gnd C_wl
Rw27_81 word27_81 word26_81 R_wl
Cwl_27_81 word27_81 gnd C_wl
Rw28_81 word28_81 word27_81 R_wl
Cwl_28_81 word28_81 gnd C_wl
Rw29_81 word29_81 word28_81 R_wl
Cwl_29_81 word29_81 gnd C_wl
Rw30_81 word30_81 word29_81 R_wl
Cwl_30_81 word30_81 gnd C_wl
Rw31_81 word31_81 word30_81 R_wl
Cwl_31_81 word31_81 gnd C_wl
Rw32_81 word32_81 word31_81 R_wl
Cwl_32_81 word32_81 gnd C_wl
Rw33_81 word33_81 word32_81 R_wl
Cwl_33_81 word33_81 gnd C_wl
Rw34_81 word34_81 word33_81 R_wl
Cwl_34_81 word34_81 gnd C_wl
Rw35_81 word35_81 word34_81 R_wl
Cwl_35_81 word35_81 gnd C_wl
Rw36_81 word36_81 word35_81 R_wl
Cwl_36_81 word36_81 gnd C_wl
Rw37_81 word37_81 word36_81 R_wl
Cwl_37_81 word37_81 gnd C_wl
Rw38_81 word38_81 word37_81 R_wl
Cwl_38_81 word38_81 gnd C_wl
Rw39_81 word39_81 word38_81 R_wl
Cwl_39_81 word39_81 gnd C_wl
Rw40_81 word40_81 word39_81 R_wl
Cwl_40_81 word40_81 gnd C_wl
Rw41_81 word41_81 word40_81 R_wl
Cwl_41_81 word41_81 gnd C_wl
Rw42_81 word42_81 word41_81 R_wl
Cwl_42_81 word42_81 gnd C_wl
Rw43_81 word43_81 word42_81 R_wl
Cwl_43_81 word43_81 gnd C_wl
Rw44_81 word44_81 word43_81 R_wl
Cwl_44_81 word44_81 gnd C_wl
Rw45_81 word45_81 word44_81 R_wl
Cwl_45_81 word45_81 gnd C_wl
Rw46_81 word46_81 word45_81 R_wl
Cwl_46_81 word46_81 gnd C_wl
Rw47_81 word47_81 word46_81 R_wl
Cwl_47_81 word47_81 gnd C_wl
Rw48_81 word48_81 word47_81 R_wl
Cwl_48_81 word48_81 gnd C_wl
Rw49_81 word49_81 word48_81 R_wl
Cwl_49_81 word49_81 gnd C_wl
Rw50_81 word50_81 word49_81 R_wl
Cwl_50_81 word50_81 gnd C_wl
Rw51_81 word51_81 word50_81 R_wl
Cwl_51_81 word51_81 gnd C_wl
Rw52_81 word52_81 word51_81 R_wl
Cwl_52_81 word52_81 gnd C_wl
Rw53_81 word53_81 word52_81 R_wl
Cwl_53_81 word53_81 gnd C_wl
Rw54_81 word54_81 word53_81 R_wl
Cwl_54_81 word54_81 gnd C_wl
Rw55_81 word55_81 word54_81 R_wl
Cwl_55_81 word55_81 gnd C_wl
Rw56_81 word56_81 word55_81 R_wl
Cwl_56_81 word56_81 gnd C_wl
Rw57_81 word57_81 word56_81 R_wl
Cwl_57_81 word57_81 gnd C_wl
Rw58_81 word58_81 word57_81 R_wl
Cwl_58_81 word58_81 gnd C_wl
Rw59_81 word59_81 word58_81 R_wl
Cwl_59_81 word59_81 gnd C_wl
Rw60_81 word60_81 word59_81 R_wl
Cwl_60_81 word60_81 gnd C_wl
Rw61_81 word61_81 word60_81 R_wl
Cwl_61_81 word61_81 gnd C_wl
Rw62_81 word62_81 word61_81 R_wl
Cwl_62_81 word62_81 gnd C_wl
Rw63_81 word63_81 word62_81 R_wl
Cwl_63_81 word63_81 gnd C_wl
Rw64_81 word64_81 word63_81 R_wl
Cwl_64_81 word64_81 gnd C_wl
Rw65_81 word65_81 word64_81 R_wl
Cwl_65_81 word65_81 gnd C_wl
Rw66_81 word66_81 word65_81 R_wl
Cwl_66_81 word66_81 gnd C_wl
Rw67_81 word67_81 word66_81 R_wl
Cwl_67_81 word67_81 gnd C_wl
Rw68_81 word68_81 word67_81 R_wl
Cwl_68_81 word68_81 gnd C_wl
Rw69_81 word69_81 word68_81 R_wl
Cwl_69_81 word69_81 gnd C_wl
Rw70_81 word70_81 word69_81 R_wl
Cwl_70_81 word70_81 gnd C_wl
Rw71_81 word71_81 word70_81 R_wl
Cwl_71_81 word71_81 gnd C_wl
Rw72_81 word72_81 word71_81 R_wl
Cwl_72_81 word72_81 gnd C_wl
Rw73_81 word73_81 word72_81 R_wl
Cwl_73_81 word73_81 gnd C_wl
Rw74_81 word74_81 word73_81 R_wl
Cwl_74_81 word74_81 gnd C_wl
Rw75_81 word75_81 word74_81 R_wl
Cwl_75_81 word75_81 gnd C_wl
Rw76_81 word76_81 word75_81 R_wl
Cwl_76_81 word76_81 gnd C_wl
Rw77_81 word77_81 word76_81 R_wl
Cwl_77_81 word77_81 gnd C_wl
Rw78_81 word78_81 word77_81 R_wl
Cwl_78_81 word78_81 gnd C_wl
Rw79_81 word79_81 word78_81 R_wl
Cwl_79_81 word79_81 gnd C_wl
Rw80_81 word80_81 word79_81 R_wl
Cwl_80_81 word80_81 gnd C_wl
Rw81_81 word81_81 word80_81 R_wl
Cwl_81_81 word81_81 gnd C_wl
Rw82_81 word82_81 word81_81 R_wl
Cwl_82_81 word82_81 gnd C_wl
Rw83_81 word83_81 word82_81 R_wl
Cwl_83_81 word83_81 gnd C_wl
Rw84_81 word84_81 word83_81 R_wl
Cwl_84_81 word84_81 gnd C_wl
Rw85_81 word85_81 word84_81 R_wl
Cwl_85_81 word85_81 gnd C_wl
Rw86_81 word86_81 word85_81 R_wl
Cwl_86_81 word86_81 gnd C_wl
Rw87_81 word87_81 word86_81 R_wl
Cwl_87_81 word87_81 gnd C_wl
Rw88_81 word88_81 word87_81 R_wl
Cwl_88_81 word88_81 gnd C_wl
Rw89_81 word89_81 word88_81 R_wl
Cwl_89_81 word89_81 gnd C_wl
Rw90_81 word90_81 word89_81 R_wl
Cwl_90_81 word90_81 gnd C_wl
Rw91_81 word91_81 word90_81 R_wl
Cwl_91_81 word91_81 gnd C_wl
Rw92_81 word92_81 word91_81 R_wl
Cwl_92_81 word92_81 gnd C_wl
Rw93_81 word93_81 word92_81 R_wl
Cwl_93_81 word93_81 gnd C_wl
Rw94_81 word94_81 word93_81 R_wl
Cwl_94_81 word94_81 gnd C_wl
Rw95_81 word95_81 word94_81 R_wl
Cwl_95_81 word95_81 gnd C_wl
Rw96_81 word96_81 word95_81 R_wl
Cwl_96_81 word96_81 gnd C_wl
Rw97_81 word97_81 word96_81 R_wl
Cwl_97_81 word97_81 gnd C_wl
Rw98_81 word98_81 word97_81 R_wl
Cwl_98_81 word98_81 gnd C_wl
Rw99_81 word99_81 word98_81 R_wl
Cwl_99_81 word99_81 gnd C_wl
Vwl_82 word_82 0 0
Rw0_82 word_82 word0_82 R_wl
Cwl_0_82 word0_82 gnd C_wl
Rw1_82 word1_82 word0_82 R_wl
Cwl_1_82 word1_82 gnd C_wl
Rw2_82 word2_82 word1_82 R_wl
Cwl_2_82 word2_82 gnd C_wl
Rw3_82 word3_82 word2_82 R_wl
Cwl_3_82 word3_82 gnd C_wl
Rw4_82 word4_82 word3_82 R_wl
Cwl_4_82 word4_82 gnd C_wl
Rw5_82 word5_82 word4_82 R_wl
Cwl_5_82 word5_82 gnd C_wl
Rw6_82 word6_82 word5_82 R_wl
Cwl_6_82 word6_82 gnd C_wl
Rw7_82 word7_82 word6_82 R_wl
Cwl_7_82 word7_82 gnd C_wl
Rw8_82 word8_82 word7_82 R_wl
Cwl_8_82 word8_82 gnd C_wl
Rw9_82 word9_82 word8_82 R_wl
Cwl_9_82 word9_82 gnd C_wl
Rw10_82 word10_82 word9_82 R_wl
Cwl_10_82 word10_82 gnd C_wl
Rw11_82 word11_82 word10_82 R_wl
Cwl_11_82 word11_82 gnd C_wl
Rw12_82 word12_82 word11_82 R_wl
Cwl_12_82 word12_82 gnd C_wl
Rw13_82 word13_82 word12_82 R_wl
Cwl_13_82 word13_82 gnd C_wl
Rw14_82 word14_82 word13_82 R_wl
Cwl_14_82 word14_82 gnd C_wl
Rw15_82 word15_82 word14_82 R_wl
Cwl_15_82 word15_82 gnd C_wl
Rw16_82 word16_82 word15_82 R_wl
Cwl_16_82 word16_82 gnd C_wl
Rw17_82 word17_82 word16_82 R_wl
Cwl_17_82 word17_82 gnd C_wl
Rw18_82 word18_82 word17_82 R_wl
Cwl_18_82 word18_82 gnd C_wl
Rw19_82 word19_82 word18_82 R_wl
Cwl_19_82 word19_82 gnd C_wl
Rw20_82 word20_82 word19_82 R_wl
Cwl_20_82 word20_82 gnd C_wl
Rw21_82 word21_82 word20_82 R_wl
Cwl_21_82 word21_82 gnd C_wl
Rw22_82 word22_82 word21_82 R_wl
Cwl_22_82 word22_82 gnd C_wl
Rw23_82 word23_82 word22_82 R_wl
Cwl_23_82 word23_82 gnd C_wl
Rw24_82 word24_82 word23_82 R_wl
Cwl_24_82 word24_82 gnd C_wl
Rw25_82 word25_82 word24_82 R_wl
Cwl_25_82 word25_82 gnd C_wl
Rw26_82 word26_82 word25_82 R_wl
Cwl_26_82 word26_82 gnd C_wl
Rw27_82 word27_82 word26_82 R_wl
Cwl_27_82 word27_82 gnd C_wl
Rw28_82 word28_82 word27_82 R_wl
Cwl_28_82 word28_82 gnd C_wl
Rw29_82 word29_82 word28_82 R_wl
Cwl_29_82 word29_82 gnd C_wl
Rw30_82 word30_82 word29_82 R_wl
Cwl_30_82 word30_82 gnd C_wl
Rw31_82 word31_82 word30_82 R_wl
Cwl_31_82 word31_82 gnd C_wl
Rw32_82 word32_82 word31_82 R_wl
Cwl_32_82 word32_82 gnd C_wl
Rw33_82 word33_82 word32_82 R_wl
Cwl_33_82 word33_82 gnd C_wl
Rw34_82 word34_82 word33_82 R_wl
Cwl_34_82 word34_82 gnd C_wl
Rw35_82 word35_82 word34_82 R_wl
Cwl_35_82 word35_82 gnd C_wl
Rw36_82 word36_82 word35_82 R_wl
Cwl_36_82 word36_82 gnd C_wl
Rw37_82 word37_82 word36_82 R_wl
Cwl_37_82 word37_82 gnd C_wl
Rw38_82 word38_82 word37_82 R_wl
Cwl_38_82 word38_82 gnd C_wl
Rw39_82 word39_82 word38_82 R_wl
Cwl_39_82 word39_82 gnd C_wl
Rw40_82 word40_82 word39_82 R_wl
Cwl_40_82 word40_82 gnd C_wl
Rw41_82 word41_82 word40_82 R_wl
Cwl_41_82 word41_82 gnd C_wl
Rw42_82 word42_82 word41_82 R_wl
Cwl_42_82 word42_82 gnd C_wl
Rw43_82 word43_82 word42_82 R_wl
Cwl_43_82 word43_82 gnd C_wl
Rw44_82 word44_82 word43_82 R_wl
Cwl_44_82 word44_82 gnd C_wl
Rw45_82 word45_82 word44_82 R_wl
Cwl_45_82 word45_82 gnd C_wl
Rw46_82 word46_82 word45_82 R_wl
Cwl_46_82 word46_82 gnd C_wl
Rw47_82 word47_82 word46_82 R_wl
Cwl_47_82 word47_82 gnd C_wl
Rw48_82 word48_82 word47_82 R_wl
Cwl_48_82 word48_82 gnd C_wl
Rw49_82 word49_82 word48_82 R_wl
Cwl_49_82 word49_82 gnd C_wl
Rw50_82 word50_82 word49_82 R_wl
Cwl_50_82 word50_82 gnd C_wl
Rw51_82 word51_82 word50_82 R_wl
Cwl_51_82 word51_82 gnd C_wl
Rw52_82 word52_82 word51_82 R_wl
Cwl_52_82 word52_82 gnd C_wl
Rw53_82 word53_82 word52_82 R_wl
Cwl_53_82 word53_82 gnd C_wl
Rw54_82 word54_82 word53_82 R_wl
Cwl_54_82 word54_82 gnd C_wl
Rw55_82 word55_82 word54_82 R_wl
Cwl_55_82 word55_82 gnd C_wl
Rw56_82 word56_82 word55_82 R_wl
Cwl_56_82 word56_82 gnd C_wl
Rw57_82 word57_82 word56_82 R_wl
Cwl_57_82 word57_82 gnd C_wl
Rw58_82 word58_82 word57_82 R_wl
Cwl_58_82 word58_82 gnd C_wl
Rw59_82 word59_82 word58_82 R_wl
Cwl_59_82 word59_82 gnd C_wl
Rw60_82 word60_82 word59_82 R_wl
Cwl_60_82 word60_82 gnd C_wl
Rw61_82 word61_82 word60_82 R_wl
Cwl_61_82 word61_82 gnd C_wl
Rw62_82 word62_82 word61_82 R_wl
Cwl_62_82 word62_82 gnd C_wl
Rw63_82 word63_82 word62_82 R_wl
Cwl_63_82 word63_82 gnd C_wl
Rw64_82 word64_82 word63_82 R_wl
Cwl_64_82 word64_82 gnd C_wl
Rw65_82 word65_82 word64_82 R_wl
Cwl_65_82 word65_82 gnd C_wl
Rw66_82 word66_82 word65_82 R_wl
Cwl_66_82 word66_82 gnd C_wl
Rw67_82 word67_82 word66_82 R_wl
Cwl_67_82 word67_82 gnd C_wl
Rw68_82 word68_82 word67_82 R_wl
Cwl_68_82 word68_82 gnd C_wl
Rw69_82 word69_82 word68_82 R_wl
Cwl_69_82 word69_82 gnd C_wl
Rw70_82 word70_82 word69_82 R_wl
Cwl_70_82 word70_82 gnd C_wl
Rw71_82 word71_82 word70_82 R_wl
Cwl_71_82 word71_82 gnd C_wl
Rw72_82 word72_82 word71_82 R_wl
Cwl_72_82 word72_82 gnd C_wl
Rw73_82 word73_82 word72_82 R_wl
Cwl_73_82 word73_82 gnd C_wl
Rw74_82 word74_82 word73_82 R_wl
Cwl_74_82 word74_82 gnd C_wl
Rw75_82 word75_82 word74_82 R_wl
Cwl_75_82 word75_82 gnd C_wl
Rw76_82 word76_82 word75_82 R_wl
Cwl_76_82 word76_82 gnd C_wl
Rw77_82 word77_82 word76_82 R_wl
Cwl_77_82 word77_82 gnd C_wl
Rw78_82 word78_82 word77_82 R_wl
Cwl_78_82 word78_82 gnd C_wl
Rw79_82 word79_82 word78_82 R_wl
Cwl_79_82 word79_82 gnd C_wl
Rw80_82 word80_82 word79_82 R_wl
Cwl_80_82 word80_82 gnd C_wl
Rw81_82 word81_82 word80_82 R_wl
Cwl_81_82 word81_82 gnd C_wl
Rw82_82 word82_82 word81_82 R_wl
Cwl_82_82 word82_82 gnd C_wl
Rw83_82 word83_82 word82_82 R_wl
Cwl_83_82 word83_82 gnd C_wl
Rw84_82 word84_82 word83_82 R_wl
Cwl_84_82 word84_82 gnd C_wl
Rw85_82 word85_82 word84_82 R_wl
Cwl_85_82 word85_82 gnd C_wl
Rw86_82 word86_82 word85_82 R_wl
Cwl_86_82 word86_82 gnd C_wl
Rw87_82 word87_82 word86_82 R_wl
Cwl_87_82 word87_82 gnd C_wl
Rw88_82 word88_82 word87_82 R_wl
Cwl_88_82 word88_82 gnd C_wl
Rw89_82 word89_82 word88_82 R_wl
Cwl_89_82 word89_82 gnd C_wl
Rw90_82 word90_82 word89_82 R_wl
Cwl_90_82 word90_82 gnd C_wl
Rw91_82 word91_82 word90_82 R_wl
Cwl_91_82 word91_82 gnd C_wl
Rw92_82 word92_82 word91_82 R_wl
Cwl_92_82 word92_82 gnd C_wl
Rw93_82 word93_82 word92_82 R_wl
Cwl_93_82 word93_82 gnd C_wl
Rw94_82 word94_82 word93_82 R_wl
Cwl_94_82 word94_82 gnd C_wl
Rw95_82 word95_82 word94_82 R_wl
Cwl_95_82 word95_82 gnd C_wl
Rw96_82 word96_82 word95_82 R_wl
Cwl_96_82 word96_82 gnd C_wl
Rw97_82 word97_82 word96_82 R_wl
Cwl_97_82 word97_82 gnd C_wl
Rw98_82 word98_82 word97_82 R_wl
Cwl_98_82 word98_82 gnd C_wl
Rw99_82 word99_82 word98_82 R_wl
Cwl_99_82 word99_82 gnd C_wl
Vwl_83 word_83 0 0
Rw0_83 word_83 word0_83 R_wl
Cwl_0_83 word0_83 gnd C_wl
Rw1_83 word1_83 word0_83 R_wl
Cwl_1_83 word1_83 gnd C_wl
Rw2_83 word2_83 word1_83 R_wl
Cwl_2_83 word2_83 gnd C_wl
Rw3_83 word3_83 word2_83 R_wl
Cwl_3_83 word3_83 gnd C_wl
Rw4_83 word4_83 word3_83 R_wl
Cwl_4_83 word4_83 gnd C_wl
Rw5_83 word5_83 word4_83 R_wl
Cwl_5_83 word5_83 gnd C_wl
Rw6_83 word6_83 word5_83 R_wl
Cwl_6_83 word6_83 gnd C_wl
Rw7_83 word7_83 word6_83 R_wl
Cwl_7_83 word7_83 gnd C_wl
Rw8_83 word8_83 word7_83 R_wl
Cwl_8_83 word8_83 gnd C_wl
Rw9_83 word9_83 word8_83 R_wl
Cwl_9_83 word9_83 gnd C_wl
Rw10_83 word10_83 word9_83 R_wl
Cwl_10_83 word10_83 gnd C_wl
Rw11_83 word11_83 word10_83 R_wl
Cwl_11_83 word11_83 gnd C_wl
Rw12_83 word12_83 word11_83 R_wl
Cwl_12_83 word12_83 gnd C_wl
Rw13_83 word13_83 word12_83 R_wl
Cwl_13_83 word13_83 gnd C_wl
Rw14_83 word14_83 word13_83 R_wl
Cwl_14_83 word14_83 gnd C_wl
Rw15_83 word15_83 word14_83 R_wl
Cwl_15_83 word15_83 gnd C_wl
Rw16_83 word16_83 word15_83 R_wl
Cwl_16_83 word16_83 gnd C_wl
Rw17_83 word17_83 word16_83 R_wl
Cwl_17_83 word17_83 gnd C_wl
Rw18_83 word18_83 word17_83 R_wl
Cwl_18_83 word18_83 gnd C_wl
Rw19_83 word19_83 word18_83 R_wl
Cwl_19_83 word19_83 gnd C_wl
Rw20_83 word20_83 word19_83 R_wl
Cwl_20_83 word20_83 gnd C_wl
Rw21_83 word21_83 word20_83 R_wl
Cwl_21_83 word21_83 gnd C_wl
Rw22_83 word22_83 word21_83 R_wl
Cwl_22_83 word22_83 gnd C_wl
Rw23_83 word23_83 word22_83 R_wl
Cwl_23_83 word23_83 gnd C_wl
Rw24_83 word24_83 word23_83 R_wl
Cwl_24_83 word24_83 gnd C_wl
Rw25_83 word25_83 word24_83 R_wl
Cwl_25_83 word25_83 gnd C_wl
Rw26_83 word26_83 word25_83 R_wl
Cwl_26_83 word26_83 gnd C_wl
Rw27_83 word27_83 word26_83 R_wl
Cwl_27_83 word27_83 gnd C_wl
Rw28_83 word28_83 word27_83 R_wl
Cwl_28_83 word28_83 gnd C_wl
Rw29_83 word29_83 word28_83 R_wl
Cwl_29_83 word29_83 gnd C_wl
Rw30_83 word30_83 word29_83 R_wl
Cwl_30_83 word30_83 gnd C_wl
Rw31_83 word31_83 word30_83 R_wl
Cwl_31_83 word31_83 gnd C_wl
Rw32_83 word32_83 word31_83 R_wl
Cwl_32_83 word32_83 gnd C_wl
Rw33_83 word33_83 word32_83 R_wl
Cwl_33_83 word33_83 gnd C_wl
Rw34_83 word34_83 word33_83 R_wl
Cwl_34_83 word34_83 gnd C_wl
Rw35_83 word35_83 word34_83 R_wl
Cwl_35_83 word35_83 gnd C_wl
Rw36_83 word36_83 word35_83 R_wl
Cwl_36_83 word36_83 gnd C_wl
Rw37_83 word37_83 word36_83 R_wl
Cwl_37_83 word37_83 gnd C_wl
Rw38_83 word38_83 word37_83 R_wl
Cwl_38_83 word38_83 gnd C_wl
Rw39_83 word39_83 word38_83 R_wl
Cwl_39_83 word39_83 gnd C_wl
Rw40_83 word40_83 word39_83 R_wl
Cwl_40_83 word40_83 gnd C_wl
Rw41_83 word41_83 word40_83 R_wl
Cwl_41_83 word41_83 gnd C_wl
Rw42_83 word42_83 word41_83 R_wl
Cwl_42_83 word42_83 gnd C_wl
Rw43_83 word43_83 word42_83 R_wl
Cwl_43_83 word43_83 gnd C_wl
Rw44_83 word44_83 word43_83 R_wl
Cwl_44_83 word44_83 gnd C_wl
Rw45_83 word45_83 word44_83 R_wl
Cwl_45_83 word45_83 gnd C_wl
Rw46_83 word46_83 word45_83 R_wl
Cwl_46_83 word46_83 gnd C_wl
Rw47_83 word47_83 word46_83 R_wl
Cwl_47_83 word47_83 gnd C_wl
Rw48_83 word48_83 word47_83 R_wl
Cwl_48_83 word48_83 gnd C_wl
Rw49_83 word49_83 word48_83 R_wl
Cwl_49_83 word49_83 gnd C_wl
Rw50_83 word50_83 word49_83 R_wl
Cwl_50_83 word50_83 gnd C_wl
Rw51_83 word51_83 word50_83 R_wl
Cwl_51_83 word51_83 gnd C_wl
Rw52_83 word52_83 word51_83 R_wl
Cwl_52_83 word52_83 gnd C_wl
Rw53_83 word53_83 word52_83 R_wl
Cwl_53_83 word53_83 gnd C_wl
Rw54_83 word54_83 word53_83 R_wl
Cwl_54_83 word54_83 gnd C_wl
Rw55_83 word55_83 word54_83 R_wl
Cwl_55_83 word55_83 gnd C_wl
Rw56_83 word56_83 word55_83 R_wl
Cwl_56_83 word56_83 gnd C_wl
Rw57_83 word57_83 word56_83 R_wl
Cwl_57_83 word57_83 gnd C_wl
Rw58_83 word58_83 word57_83 R_wl
Cwl_58_83 word58_83 gnd C_wl
Rw59_83 word59_83 word58_83 R_wl
Cwl_59_83 word59_83 gnd C_wl
Rw60_83 word60_83 word59_83 R_wl
Cwl_60_83 word60_83 gnd C_wl
Rw61_83 word61_83 word60_83 R_wl
Cwl_61_83 word61_83 gnd C_wl
Rw62_83 word62_83 word61_83 R_wl
Cwl_62_83 word62_83 gnd C_wl
Rw63_83 word63_83 word62_83 R_wl
Cwl_63_83 word63_83 gnd C_wl
Rw64_83 word64_83 word63_83 R_wl
Cwl_64_83 word64_83 gnd C_wl
Rw65_83 word65_83 word64_83 R_wl
Cwl_65_83 word65_83 gnd C_wl
Rw66_83 word66_83 word65_83 R_wl
Cwl_66_83 word66_83 gnd C_wl
Rw67_83 word67_83 word66_83 R_wl
Cwl_67_83 word67_83 gnd C_wl
Rw68_83 word68_83 word67_83 R_wl
Cwl_68_83 word68_83 gnd C_wl
Rw69_83 word69_83 word68_83 R_wl
Cwl_69_83 word69_83 gnd C_wl
Rw70_83 word70_83 word69_83 R_wl
Cwl_70_83 word70_83 gnd C_wl
Rw71_83 word71_83 word70_83 R_wl
Cwl_71_83 word71_83 gnd C_wl
Rw72_83 word72_83 word71_83 R_wl
Cwl_72_83 word72_83 gnd C_wl
Rw73_83 word73_83 word72_83 R_wl
Cwl_73_83 word73_83 gnd C_wl
Rw74_83 word74_83 word73_83 R_wl
Cwl_74_83 word74_83 gnd C_wl
Rw75_83 word75_83 word74_83 R_wl
Cwl_75_83 word75_83 gnd C_wl
Rw76_83 word76_83 word75_83 R_wl
Cwl_76_83 word76_83 gnd C_wl
Rw77_83 word77_83 word76_83 R_wl
Cwl_77_83 word77_83 gnd C_wl
Rw78_83 word78_83 word77_83 R_wl
Cwl_78_83 word78_83 gnd C_wl
Rw79_83 word79_83 word78_83 R_wl
Cwl_79_83 word79_83 gnd C_wl
Rw80_83 word80_83 word79_83 R_wl
Cwl_80_83 word80_83 gnd C_wl
Rw81_83 word81_83 word80_83 R_wl
Cwl_81_83 word81_83 gnd C_wl
Rw82_83 word82_83 word81_83 R_wl
Cwl_82_83 word82_83 gnd C_wl
Rw83_83 word83_83 word82_83 R_wl
Cwl_83_83 word83_83 gnd C_wl
Rw84_83 word84_83 word83_83 R_wl
Cwl_84_83 word84_83 gnd C_wl
Rw85_83 word85_83 word84_83 R_wl
Cwl_85_83 word85_83 gnd C_wl
Rw86_83 word86_83 word85_83 R_wl
Cwl_86_83 word86_83 gnd C_wl
Rw87_83 word87_83 word86_83 R_wl
Cwl_87_83 word87_83 gnd C_wl
Rw88_83 word88_83 word87_83 R_wl
Cwl_88_83 word88_83 gnd C_wl
Rw89_83 word89_83 word88_83 R_wl
Cwl_89_83 word89_83 gnd C_wl
Rw90_83 word90_83 word89_83 R_wl
Cwl_90_83 word90_83 gnd C_wl
Rw91_83 word91_83 word90_83 R_wl
Cwl_91_83 word91_83 gnd C_wl
Rw92_83 word92_83 word91_83 R_wl
Cwl_92_83 word92_83 gnd C_wl
Rw93_83 word93_83 word92_83 R_wl
Cwl_93_83 word93_83 gnd C_wl
Rw94_83 word94_83 word93_83 R_wl
Cwl_94_83 word94_83 gnd C_wl
Rw95_83 word95_83 word94_83 R_wl
Cwl_95_83 word95_83 gnd C_wl
Rw96_83 word96_83 word95_83 R_wl
Cwl_96_83 word96_83 gnd C_wl
Rw97_83 word97_83 word96_83 R_wl
Cwl_97_83 word97_83 gnd C_wl
Rw98_83 word98_83 word97_83 R_wl
Cwl_98_83 word98_83 gnd C_wl
Rw99_83 word99_83 word98_83 R_wl
Cwl_99_83 word99_83 gnd C_wl
Vwl_84 word_84 0 0
Rw0_84 word_84 word0_84 R_wl
Cwl_0_84 word0_84 gnd C_wl
Rw1_84 word1_84 word0_84 R_wl
Cwl_1_84 word1_84 gnd C_wl
Rw2_84 word2_84 word1_84 R_wl
Cwl_2_84 word2_84 gnd C_wl
Rw3_84 word3_84 word2_84 R_wl
Cwl_3_84 word3_84 gnd C_wl
Rw4_84 word4_84 word3_84 R_wl
Cwl_4_84 word4_84 gnd C_wl
Rw5_84 word5_84 word4_84 R_wl
Cwl_5_84 word5_84 gnd C_wl
Rw6_84 word6_84 word5_84 R_wl
Cwl_6_84 word6_84 gnd C_wl
Rw7_84 word7_84 word6_84 R_wl
Cwl_7_84 word7_84 gnd C_wl
Rw8_84 word8_84 word7_84 R_wl
Cwl_8_84 word8_84 gnd C_wl
Rw9_84 word9_84 word8_84 R_wl
Cwl_9_84 word9_84 gnd C_wl
Rw10_84 word10_84 word9_84 R_wl
Cwl_10_84 word10_84 gnd C_wl
Rw11_84 word11_84 word10_84 R_wl
Cwl_11_84 word11_84 gnd C_wl
Rw12_84 word12_84 word11_84 R_wl
Cwl_12_84 word12_84 gnd C_wl
Rw13_84 word13_84 word12_84 R_wl
Cwl_13_84 word13_84 gnd C_wl
Rw14_84 word14_84 word13_84 R_wl
Cwl_14_84 word14_84 gnd C_wl
Rw15_84 word15_84 word14_84 R_wl
Cwl_15_84 word15_84 gnd C_wl
Rw16_84 word16_84 word15_84 R_wl
Cwl_16_84 word16_84 gnd C_wl
Rw17_84 word17_84 word16_84 R_wl
Cwl_17_84 word17_84 gnd C_wl
Rw18_84 word18_84 word17_84 R_wl
Cwl_18_84 word18_84 gnd C_wl
Rw19_84 word19_84 word18_84 R_wl
Cwl_19_84 word19_84 gnd C_wl
Rw20_84 word20_84 word19_84 R_wl
Cwl_20_84 word20_84 gnd C_wl
Rw21_84 word21_84 word20_84 R_wl
Cwl_21_84 word21_84 gnd C_wl
Rw22_84 word22_84 word21_84 R_wl
Cwl_22_84 word22_84 gnd C_wl
Rw23_84 word23_84 word22_84 R_wl
Cwl_23_84 word23_84 gnd C_wl
Rw24_84 word24_84 word23_84 R_wl
Cwl_24_84 word24_84 gnd C_wl
Rw25_84 word25_84 word24_84 R_wl
Cwl_25_84 word25_84 gnd C_wl
Rw26_84 word26_84 word25_84 R_wl
Cwl_26_84 word26_84 gnd C_wl
Rw27_84 word27_84 word26_84 R_wl
Cwl_27_84 word27_84 gnd C_wl
Rw28_84 word28_84 word27_84 R_wl
Cwl_28_84 word28_84 gnd C_wl
Rw29_84 word29_84 word28_84 R_wl
Cwl_29_84 word29_84 gnd C_wl
Rw30_84 word30_84 word29_84 R_wl
Cwl_30_84 word30_84 gnd C_wl
Rw31_84 word31_84 word30_84 R_wl
Cwl_31_84 word31_84 gnd C_wl
Rw32_84 word32_84 word31_84 R_wl
Cwl_32_84 word32_84 gnd C_wl
Rw33_84 word33_84 word32_84 R_wl
Cwl_33_84 word33_84 gnd C_wl
Rw34_84 word34_84 word33_84 R_wl
Cwl_34_84 word34_84 gnd C_wl
Rw35_84 word35_84 word34_84 R_wl
Cwl_35_84 word35_84 gnd C_wl
Rw36_84 word36_84 word35_84 R_wl
Cwl_36_84 word36_84 gnd C_wl
Rw37_84 word37_84 word36_84 R_wl
Cwl_37_84 word37_84 gnd C_wl
Rw38_84 word38_84 word37_84 R_wl
Cwl_38_84 word38_84 gnd C_wl
Rw39_84 word39_84 word38_84 R_wl
Cwl_39_84 word39_84 gnd C_wl
Rw40_84 word40_84 word39_84 R_wl
Cwl_40_84 word40_84 gnd C_wl
Rw41_84 word41_84 word40_84 R_wl
Cwl_41_84 word41_84 gnd C_wl
Rw42_84 word42_84 word41_84 R_wl
Cwl_42_84 word42_84 gnd C_wl
Rw43_84 word43_84 word42_84 R_wl
Cwl_43_84 word43_84 gnd C_wl
Rw44_84 word44_84 word43_84 R_wl
Cwl_44_84 word44_84 gnd C_wl
Rw45_84 word45_84 word44_84 R_wl
Cwl_45_84 word45_84 gnd C_wl
Rw46_84 word46_84 word45_84 R_wl
Cwl_46_84 word46_84 gnd C_wl
Rw47_84 word47_84 word46_84 R_wl
Cwl_47_84 word47_84 gnd C_wl
Rw48_84 word48_84 word47_84 R_wl
Cwl_48_84 word48_84 gnd C_wl
Rw49_84 word49_84 word48_84 R_wl
Cwl_49_84 word49_84 gnd C_wl
Rw50_84 word50_84 word49_84 R_wl
Cwl_50_84 word50_84 gnd C_wl
Rw51_84 word51_84 word50_84 R_wl
Cwl_51_84 word51_84 gnd C_wl
Rw52_84 word52_84 word51_84 R_wl
Cwl_52_84 word52_84 gnd C_wl
Rw53_84 word53_84 word52_84 R_wl
Cwl_53_84 word53_84 gnd C_wl
Rw54_84 word54_84 word53_84 R_wl
Cwl_54_84 word54_84 gnd C_wl
Rw55_84 word55_84 word54_84 R_wl
Cwl_55_84 word55_84 gnd C_wl
Rw56_84 word56_84 word55_84 R_wl
Cwl_56_84 word56_84 gnd C_wl
Rw57_84 word57_84 word56_84 R_wl
Cwl_57_84 word57_84 gnd C_wl
Rw58_84 word58_84 word57_84 R_wl
Cwl_58_84 word58_84 gnd C_wl
Rw59_84 word59_84 word58_84 R_wl
Cwl_59_84 word59_84 gnd C_wl
Rw60_84 word60_84 word59_84 R_wl
Cwl_60_84 word60_84 gnd C_wl
Rw61_84 word61_84 word60_84 R_wl
Cwl_61_84 word61_84 gnd C_wl
Rw62_84 word62_84 word61_84 R_wl
Cwl_62_84 word62_84 gnd C_wl
Rw63_84 word63_84 word62_84 R_wl
Cwl_63_84 word63_84 gnd C_wl
Rw64_84 word64_84 word63_84 R_wl
Cwl_64_84 word64_84 gnd C_wl
Rw65_84 word65_84 word64_84 R_wl
Cwl_65_84 word65_84 gnd C_wl
Rw66_84 word66_84 word65_84 R_wl
Cwl_66_84 word66_84 gnd C_wl
Rw67_84 word67_84 word66_84 R_wl
Cwl_67_84 word67_84 gnd C_wl
Rw68_84 word68_84 word67_84 R_wl
Cwl_68_84 word68_84 gnd C_wl
Rw69_84 word69_84 word68_84 R_wl
Cwl_69_84 word69_84 gnd C_wl
Rw70_84 word70_84 word69_84 R_wl
Cwl_70_84 word70_84 gnd C_wl
Rw71_84 word71_84 word70_84 R_wl
Cwl_71_84 word71_84 gnd C_wl
Rw72_84 word72_84 word71_84 R_wl
Cwl_72_84 word72_84 gnd C_wl
Rw73_84 word73_84 word72_84 R_wl
Cwl_73_84 word73_84 gnd C_wl
Rw74_84 word74_84 word73_84 R_wl
Cwl_74_84 word74_84 gnd C_wl
Rw75_84 word75_84 word74_84 R_wl
Cwl_75_84 word75_84 gnd C_wl
Rw76_84 word76_84 word75_84 R_wl
Cwl_76_84 word76_84 gnd C_wl
Rw77_84 word77_84 word76_84 R_wl
Cwl_77_84 word77_84 gnd C_wl
Rw78_84 word78_84 word77_84 R_wl
Cwl_78_84 word78_84 gnd C_wl
Rw79_84 word79_84 word78_84 R_wl
Cwl_79_84 word79_84 gnd C_wl
Rw80_84 word80_84 word79_84 R_wl
Cwl_80_84 word80_84 gnd C_wl
Rw81_84 word81_84 word80_84 R_wl
Cwl_81_84 word81_84 gnd C_wl
Rw82_84 word82_84 word81_84 R_wl
Cwl_82_84 word82_84 gnd C_wl
Rw83_84 word83_84 word82_84 R_wl
Cwl_83_84 word83_84 gnd C_wl
Rw84_84 word84_84 word83_84 R_wl
Cwl_84_84 word84_84 gnd C_wl
Rw85_84 word85_84 word84_84 R_wl
Cwl_85_84 word85_84 gnd C_wl
Rw86_84 word86_84 word85_84 R_wl
Cwl_86_84 word86_84 gnd C_wl
Rw87_84 word87_84 word86_84 R_wl
Cwl_87_84 word87_84 gnd C_wl
Rw88_84 word88_84 word87_84 R_wl
Cwl_88_84 word88_84 gnd C_wl
Rw89_84 word89_84 word88_84 R_wl
Cwl_89_84 word89_84 gnd C_wl
Rw90_84 word90_84 word89_84 R_wl
Cwl_90_84 word90_84 gnd C_wl
Rw91_84 word91_84 word90_84 R_wl
Cwl_91_84 word91_84 gnd C_wl
Rw92_84 word92_84 word91_84 R_wl
Cwl_92_84 word92_84 gnd C_wl
Rw93_84 word93_84 word92_84 R_wl
Cwl_93_84 word93_84 gnd C_wl
Rw94_84 word94_84 word93_84 R_wl
Cwl_94_84 word94_84 gnd C_wl
Rw95_84 word95_84 word94_84 R_wl
Cwl_95_84 word95_84 gnd C_wl
Rw96_84 word96_84 word95_84 R_wl
Cwl_96_84 word96_84 gnd C_wl
Rw97_84 word97_84 word96_84 R_wl
Cwl_97_84 word97_84 gnd C_wl
Rw98_84 word98_84 word97_84 R_wl
Cwl_98_84 word98_84 gnd C_wl
Rw99_84 word99_84 word98_84 R_wl
Cwl_99_84 word99_84 gnd C_wl
Vwl_85 word_85 0 0
Rw0_85 word_85 word0_85 R_wl
Cwl_0_85 word0_85 gnd C_wl
Rw1_85 word1_85 word0_85 R_wl
Cwl_1_85 word1_85 gnd C_wl
Rw2_85 word2_85 word1_85 R_wl
Cwl_2_85 word2_85 gnd C_wl
Rw3_85 word3_85 word2_85 R_wl
Cwl_3_85 word3_85 gnd C_wl
Rw4_85 word4_85 word3_85 R_wl
Cwl_4_85 word4_85 gnd C_wl
Rw5_85 word5_85 word4_85 R_wl
Cwl_5_85 word5_85 gnd C_wl
Rw6_85 word6_85 word5_85 R_wl
Cwl_6_85 word6_85 gnd C_wl
Rw7_85 word7_85 word6_85 R_wl
Cwl_7_85 word7_85 gnd C_wl
Rw8_85 word8_85 word7_85 R_wl
Cwl_8_85 word8_85 gnd C_wl
Rw9_85 word9_85 word8_85 R_wl
Cwl_9_85 word9_85 gnd C_wl
Rw10_85 word10_85 word9_85 R_wl
Cwl_10_85 word10_85 gnd C_wl
Rw11_85 word11_85 word10_85 R_wl
Cwl_11_85 word11_85 gnd C_wl
Rw12_85 word12_85 word11_85 R_wl
Cwl_12_85 word12_85 gnd C_wl
Rw13_85 word13_85 word12_85 R_wl
Cwl_13_85 word13_85 gnd C_wl
Rw14_85 word14_85 word13_85 R_wl
Cwl_14_85 word14_85 gnd C_wl
Rw15_85 word15_85 word14_85 R_wl
Cwl_15_85 word15_85 gnd C_wl
Rw16_85 word16_85 word15_85 R_wl
Cwl_16_85 word16_85 gnd C_wl
Rw17_85 word17_85 word16_85 R_wl
Cwl_17_85 word17_85 gnd C_wl
Rw18_85 word18_85 word17_85 R_wl
Cwl_18_85 word18_85 gnd C_wl
Rw19_85 word19_85 word18_85 R_wl
Cwl_19_85 word19_85 gnd C_wl
Rw20_85 word20_85 word19_85 R_wl
Cwl_20_85 word20_85 gnd C_wl
Rw21_85 word21_85 word20_85 R_wl
Cwl_21_85 word21_85 gnd C_wl
Rw22_85 word22_85 word21_85 R_wl
Cwl_22_85 word22_85 gnd C_wl
Rw23_85 word23_85 word22_85 R_wl
Cwl_23_85 word23_85 gnd C_wl
Rw24_85 word24_85 word23_85 R_wl
Cwl_24_85 word24_85 gnd C_wl
Rw25_85 word25_85 word24_85 R_wl
Cwl_25_85 word25_85 gnd C_wl
Rw26_85 word26_85 word25_85 R_wl
Cwl_26_85 word26_85 gnd C_wl
Rw27_85 word27_85 word26_85 R_wl
Cwl_27_85 word27_85 gnd C_wl
Rw28_85 word28_85 word27_85 R_wl
Cwl_28_85 word28_85 gnd C_wl
Rw29_85 word29_85 word28_85 R_wl
Cwl_29_85 word29_85 gnd C_wl
Rw30_85 word30_85 word29_85 R_wl
Cwl_30_85 word30_85 gnd C_wl
Rw31_85 word31_85 word30_85 R_wl
Cwl_31_85 word31_85 gnd C_wl
Rw32_85 word32_85 word31_85 R_wl
Cwl_32_85 word32_85 gnd C_wl
Rw33_85 word33_85 word32_85 R_wl
Cwl_33_85 word33_85 gnd C_wl
Rw34_85 word34_85 word33_85 R_wl
Cwl_34_85 word34_85 gnd C_wl
Rw35_85 word35_85 word34_85 R_wl
Cwl_35_85 word35_85 gnd C_wl
Rw36_85 word36_85 word35_85 R_wl
Cwl_36_85 word36_85 gnd C_wl
Rw37_85 word37_85 word36_85 R_wl
Cwl_37_85 word37_85 gnd C_wl
Rw38_85 word38_85 word37_85 R_wl
Cwl_38_85 word38_85 gnd C_wl
Rw39_85 word39_85 word38_85 R_wl
Cwl_39_85 word39_85 gnd C_wl
Rw40_85 word40_85 word39_85 R_wl
Cwl_40_85 word40_85 gnd C_wl
Rw41_85 word41_85 word40_85 R_wl
Cwl_41_85 word41_85 gnd C_wl
Rw42_85 word42_85 word41_85 R_wl
Cwl_42_85 word42_85 gnd C_wl
Rw43_85 word43_85 word42_85 R_wl
Cwl_43_85 word43_85 gnd C_wl
Rw44_85 word44_85 word43_85 R_wl
Cwl_44_85 word44_85 gnd C_wl
Rw45_85 word45_85 word44_85 R_wl
Cwl_45_85 word45_85 gnd C_wl
Rw46_85 word46_85 word45_85 R_wl
Cwl_46_85 word46_85 gnd C_wl
Rw47_85 word47_85 word46_85 R_wl
Cwl_47_85 word47_85 gnd C_wl
Rw48_85 word48_85 word47_85 R_wl
Cwl_48_85 word48_85 gnd C_wl
Rw49_85 word49_85 word48_85 R_wl
Cwl_49_85 word49_85 gnd C_wl
Rw50_85 word50_85 word49_85 R_wl
Cwl_50_85 word50_85 gnd C_wl
Rw51_85 word51_85 word50_85 R_wl
Cwl_51_85 word51_85 gnd C_wl
Rw52_85 word52_85 word51_85 R_wl
Cwl_52_85 word52_85 gnd C_wl
Rw53_85 word53_85 word52_85 R_wl
Cwl_53_85 word53_85 gnd C_wl
Rw54_85 word54_85 word53_85 R_wl
Cwl_54_85 word54_85 gnd C_wl
Rw55_85 word55_85 word54_85 R_wl
Cwl_55_85 word55_85 gnd C_wl
Rw56_85 word56_85 word55_85 R_wl
Cwl_56_85 word56_85 gnd C_wl
Rw57_85 word57_85 word56_85 R_wl
Cwl_57_85 word57_85 gnd C_wl
Rw58_85 word58_85 word57_85 R_wl
Cwl_58_85 word58_85 gnd C_wl
Rw59_85 word59_85 word58_85 R_wl
Cwl_59_85 word59_85 gnd C_wl
Rw60_85 word60_85 word59_85 R_wl
Cwl_60_85 word60_85 gnd C_wl
Rw61_85 word61_85 word60_85 R_wl
Cwl_61_85 word61_85 gnd C_wl
Rw62_85 word62_85 word61_85 R_wl
Cwl_62_85 word62_85 gnd C_wl
Rw63_85 word63_85 word62_85 R_wl
Cwl_63_85 word63_85 gnd C_wl
Rw64_85 word64_85 word63_85 R_wl
Cwl_64_85 word64_85 gnd C_wl
Rw65_85 word65_85 word64_85 R_wl
Cwl_65_85 word65_85 gnd C_wl
Rw66_85 word66_85 word65_85 R_wl
Cwl_66_85 word66_85 gnd C_wl
Rw67_85 word67_85 word66_85 R_wl
Cwl_67_85 word67_85 gnd C_wl
Rw68_85 word68_85 word67_85 R_wl
Cwl_68_85 word68_85 gnd C_wl
Rw69_85 word69_85 word68_85 R_wl
Cwl_69_85 word69_85 gnd C_wl
Rw70_85 word70_85 word69_85 R_wl
Cwl_70_85 word70_85 gnd C_wl
Rw71_85 word71_85 word70_85 R_wl
Cwl_71_85 word71_85 gnd C_wl
Rw72_85 word72_85 word71_85 R_wl
Cwl_72_85 word72_85 gnd C_wl
Rw73_85 word73_85 word72_85 R_wl
Cwl_73_85 word73_85 gnd C_wl
Rw74_85 word74_85 word73_85 R_wl
Cwl_74_85 word74_85 gnd C_wl
Rw75_85 word75_85 word74_85 R_wl
Cwl_75_85 word75_85 gnd C_wl
Rw76_85 word76_85 word75_85 R_wl
Cwl_76_85 word76_85 gnd C_wl
Rw77_85 word77_85 word76_85 R_wl
Cwl_77_85 word77_85 gnd C_wl
Rw78_85 word78_85 word77_85 R_wl
Cwl_78_85 word78_85 gnd C_wl
Rw79_85 word79_85 word78_85 R_wl
Cwl_79_85 word79_85 gnd C_wl
Rw80_85 word80_85 word79_85 R_wl
Cwl_80_85 word80_85 gnd C_wl
Rw81_85 word81_85 word80_85 R_wl
Cwl_81_85 word81_85 gnd C_wl
Rw82_85 word82_85 word81_85 R_wl
Cwl_82_85 word82_85 gnd C_wl
Rw83_85 word83_85 word82_85 R_wl
Cwl_83_85 word83_85 gnd C_wl
Rw84_85 word84_85 word83_85 R_wl
Cwl_84_85 word84_85 gnd C_wl
Rw85_85 word85_85 word84_85 R_wl
Cwl_85_85 word85_85 gnd C_wl
Rw86_85 word86_85 word85_85 R_wl
Cwl_86_85 word86_85 gnd C_wl
Rw87_85 word87_85 word86_85 R_wl
Cwl_87_85 word87_85 gnd C_wl
Rw88_85 word88_85 word87_85 R_wl
Cwl_88_85 word88_85 gnd C_wl
Rw89_85 word89_85 word88_85 R_wl
Cwl_89_85 word89_85 gnd C_wl
Rw90_85 word90_85 word89_85 R_wl
Cwl_90_85 word90_85 gnd C_wl
Rw91_85 word91_85 word90_85 R_wl
Cwl_91_85 word91_85 gnd C_wl
Rw92_85 word92_85 word91_85 R_wl
Cwl_92_85 word92_85 gnd C_wl
Rw93_85 word93_85 word92_85 R_wl
Cwl_93_85 word93_85 gnd C_wl
Rw94_85 word94_85 word93_85 R_wl
Cwl_94_85 word94_85 gnd C_wl
Rw95_85 word95_85 word94_85 R_wl
Cwl_95_85 word95_85 gnd C_wl
Rw96_85 word96_85 word95_85 R_wl
Cwl_96_85 word96_85 gnd C_wl
Rw97_85 word97_85 word96_85 R_wl
Cwl_97_85 word97_85 gnd C_wl
Rw98_85 word98_85 word97_85 R_wl
Cwl_98_85 word98_85 gnd C_wl
Rw99_85 word99_85 word98_85 R_wl
Cwl_99_85 word99_85 gnd C_wl
Vwl_86 word_86 0 0
Rw0_86 word_86 word0_86 R_wl
Cwl_0_86 word0_86 gnd C_wl
Rw1_86 word1_86 word0_86 R_wl
Cwl_1_86 word1_86 gnd C_wl
Rw2_86 word2_86 word1_86 R_wl
Cwl_2_86 word2_86 gnd C_wl
Rw3_86 word3_86 word2_86 R_wl
Cwl_3_86 word3_86 gnd C_wl
Rw4_86 word4_86 word3_86 R_wl
Cwl_4_86 word4_86 gnd C_wl
Rw5_86 word5_86 word4_86 R_wl
Cwl_5_86 word5_86 gnd C_wl
Rw6_86 word6_86 word5_86 R_wl
Cwl_6_86 word6_86 gnd C_wl
Rw7_86 word7_86 word6_86 R_wl
Cwl_7_86 word7_86 gnd C_wl
Rw8_86 word8_86 word7_86 R_wl
Cwl_8_86 word8_86 gnd C_wl
Rw9_86 word9_86 word8_86 R_wl
Cwl_9_86 word9_86 gnd C_wl
Rw10_86 word10_86 word9_86 R_wl
Cwl_10_86 word10_86 gnd C_wl
Rw11_86 word11_86 word10_86 R_wl
Cwl_11_86 word11_86 gnd C_wl
Rw12_86 word12_86 word11_86 R_wl
Cwl_12_86 word12_86 gnd C_wl
Rw13_86 word13_86 word12_86 R_wl
Cwl_13_86 word13_86 gnd C_wl
Rw14_86 word14_86 word13_86 R_wl
Cwl_14_86 word14_86 gnd C_wl
Rw15_86 word15_86 word14_86 R_wl
Cwl_15_86 word15_86 gnd C_wl
Rw16_86 word16_86 word15_86 R_wl
Cwl_16_86 word16_86 gnd C_wl
Rw17_86 word17_86 word16_86 R_wl
Cwl_17_86 word17_86 gnd C_wl
Rw18_86 word18_86 word17_86 R_wl
Cwl_18_86 word18_86 gnd C_wl
Rw19_86 word19_86 word18_86 R_wl
Cwl_19_86 word19_86 gnd C_wl
Rw20_86 word20_86 word19_86 R_wl
Cwl_20_86 word20_86 gnd C_wl
Rw21_86 word21_86 word20_86 R_wl
Cwl_21_86 word21_86 gnd C_wl
Rw22_86 word22_86 word21_86 R_wl
Cwl_22_86 word22_86 gnd C_wl
Rw23_86 word23_86 word22_86 R_wl
Cwl_23_86 word23_86 gnd C_wl
Rw24_86 word24_86 word23_86 R_wl
Cwl_24_86 word24_86 gnd C_wl
Rw25_86 word25_86 word24_86 R_wl
Cwl_25_86 word25_86 gnd C_wl
Rw26_86 word26_86 word25_86 R_wl
Cwl_26_86 word26_86 gnd C_wl
Rw27_86 word27_86 word26_86 R_wl
Cwl_27_86 word27_86 gnd C_wl
Rw28_86 word28_86 word27_86 R_wl
Cwl_28_86 word28_86 gnd C_wl
Rw29_86 word29_86 word28_86 R_wl
Cwl_29_86 word29_86 gnd C_wl
Rw30_86 word30_86 word29_86 R_wl
Cwl_30_86 word30_86 gnd C_wl
Rw31_86 word31_86 word30_86 R_wl
Cwl_31_86 word31_86 gnd C_wl
Rw32_86 word32_86 word31_86 R_wl
Cwl_32_86 word32_86 gnd C_wl
Rw33_86 word33_86 word32_86 R_wl
Cwl_33_86 word33_86 gnd C_wl
Rw34_86 word34_86 word33_86 R_wl
Cwl_34_86 word34_86 gnd C_wl
Rw35_86 word35_86 word34_86 R_wl
Cwl_35_86 word35_86 gnd C_wl
Rw36_86 word36_86 word35_86 R_wl
Cwl_36_86 word36_86 gnd C_wl
Rw37_86 word37_86 word36_86 R_wl
Cwl_37_86 word37_86 gnd C_wl
Rw38_86 word38_86 word37_86 R_wl
Cwl_38_86 word38_86 gnd C_wl
Rw39_86 word39_86 word38_86 R_wl
Cwl_39_86 word39_86 gnd C_wl
Rw40_86 word40_86 word39_86 R_wl
Cwl_40_86 word40_86 gnd C_wl
Rw41_86 word41_86 word40_86 R_wl
Cwl_41_86 word41_86 gnd C_wl
Rw42_86 word42_86 word41_86 R_wl
Cwl_42_86 word42_86 gnd C_wl
Rw43_86 word43_86 word42_86 R_wl
Cwl_43_86 word43_86 gnd C_wl
Rw44_86 word44_86 word43_86 R_wl
Cwl_44_86 word44_86 gnd C_wl
Rw45_86 word45_86 word44_86 R_wl
Cwl_45_86 word45_86 gnd C_wl
Rw46_86 word46_86 word45_86 R_wl
Cwl_46_86 word46_86 gnd C_wl
Rw47_86 word47_86 word46_86 R_wl
Cwl_47_86 word47_86 gnd C_wl
Rw48_86 word48_86 word47_86 R_wl
Cwl_48_86 word48_86 gnd C_wl
Rw49_86 word49_86 word48_86 R_wl
Cwl_49_86 word49_86 gnd C_wl
Rw50_86 word50_86 word49_86 R_wl
Cwl_50_86 word50_86 gnd C_wl
Rw51_86 word51_86 word50_86 R_wl
Cwl_51_86 word51_86 gnd C_wl
Rw52_86 word52_86 word51_86 R_wl
Cwl_52_86 word52_86 gnd C_wl
Rw53_86 word53_86 word52_86 R_wl
Cwl_53_86 word53_86 gnd C_wl
Rw54_86 word54_86 word53_86 R_wl
Cwl_54_86 word54_86 gnd C_wl
Rw55_86 word55_86 word54_86 R_wl
Cwl_55_86 word55_86 gnd C_wl
Rw56_86 word56_86 word55_86 R_wl
Cwl_56_86 word56_86 gnd C_wl
Rw57_86 word57_86 word56_86 R_wl
Cwl_57_86 word57_86 gnd C_wl
Rw58_86 word58_86 word57_86 R_wl
Cwl_58_86 word58_86 gnd C_wl
Rw59_86 word59_86 word58_86 R_wl
Cwl_59_86 word59_86 gnd C_wl
Rw60_86 word60_86 word59_86 R_wl
Cwl_60_86 word60_86 gnd C_wl
Rw61_86 word61_86 word60_86 R_wl
Cwl_61_86 word61_86 gnd C_wl
Rw62_86 word62_86 word61_86 R_wl
Cwl_62_86 word62_86 gnd C_wl
Rw63_86 word63_86 word62_86 R_wl
Cwl_63_86 word63_86 gnd C_wl
Rw64_86 word64_86 word63_86 R_wl
Cwl_64_86 word64_86 gnd C_wl
Rw65_86 word65_86 word64_86 R_wl
Cwl_65_86 word65_86 gnd C_wl
Rw66_86 word66_86 word65_86 R_wl
Cwl_66_86 word66_86 gnd C_wl
Rw67_86 word67_86 word66_86 R_wl
Cwl_67_86 word67_86 gnd C_wl
Rw68_86 word68_86 word67_86 R_wl
Cwl_68_86 word68_86 gnd C_wl
Rw69_86 word69_86 word68_86 R_wl
Cwl_69_86 word69_86 gnd C_wl
Rw70_86 word70_86 word69_86 R_wl
Cwl_70_86 word70_86 gnd C_wl
Rw71_86 word71_86 word70_86 R_wl
Cwl_71_86 word71_86 gnd C_wl
Rw72_86 word72_86 word71_86 R_wl
Cwl_72_86 word72_86 gnd C_wl
Rw73_86 word73_86 word72_86 R_wl
Cwl_73_86 word73_86 gnd C_wl
Rw74_86 word74_86 word73_86 R_wl
Cwl_74_86 word74_86 gnd C_wl
Rw75_86 word75_86 word74_86 R_wl
Cwl_75_86 word75_86 gnd C_wl
Rw76_86 word76_86 word75_86 R_wl
Cwl_76_86 word76_86 gnd C_wl
Rw77_86 word77_86 word76_86 R_wl
Cwl_77_86 word77_86 gnd C_wl
Rw78_86 word78_86 word77_86 R_wl
Cwl_78_86 word78_86 gnd C_wl
Rw79_86 word79_86 word78_86 R_wl
Cwl_79_86 word79_86 gnd C_wl
Rw80_86 word80_86 word79_86 R_wl
Cwl_80_86 word80_86 gnd C_wl
Rw81_86 word81_86 word80_86 R_wl
Cwl_81_86 word81_86 gnd C_wl
Rw82_86 word82_86 word81_86 R_wl
Cwl_82_86 word82_86 gnd C_wl
Rw83_86 word83_86 word82_86 R_wl
Cwl_83_86 word83_86 gnd C_wl
Rw84_86 word84_86 word83_86 R_wl
Cwl_84_86 word84_86 gnd C_wl
Rw85_86 word85_86 word84_86 R_wl
Cwl_85_86 word85_86 gnd C_wl
Rw86_86 word86_86 word85_86 R_wl
Cwl_86_86 word86_86 gnd C_wl
Rw87_86 word87_86 word86_86 R_wl
Cwl_87_86 word87_86 gnd C_wl
Rw88_86 word88_86 word87_86 R_wl
Cwl_88_86 word88_86 gnd C_wl
Rw89_86 word89_86 word88_86 R_wl
Cwl_89_86 word89_86 gnd C_wl
Rw90_86 word90_86 word89_86 R_wl
Cwl_90_86 word90_86 gnd C_wl
Rw91_86 word91_86 word90_86 R_wl
Cwl_91_86 word91_86 gnd C_wl
Rw92_86 word92_86 word91_86 R_wl
Cwl_92_86 word92_86 gnd C_wl
Rw93_86 word93_86 word92_86 R_wl
Cwl_93_86 word93_86 gnd C_wl
Rw94_86 word94_86 word93_86 R_wl
Cwl_94_86 word94_86 gnd C_wl
Rw95_86 word95_86 word94_86 R_wl
Cwl_95_86 word95_86 gnd C_wl
Rw96_86 word96_86 word95_86 R_wl
Cwl_96_86 word96_86 gnd C_wl
Rw97_86 word97_86 word96_86 R_wl
Cwl_97_86 word97_86 gnd C_wl
Rw98_86 word98_86 word97_86 R_wl
Cwl_98_86 word98_86 gnd C_wl
Rw99_86 word99_86 word98_86 R_wl
Cwl_99_86 word99_86 gnd C_wl
Vwl_87 word_87 0 0
Rw0_87 word_87 word0_87 R_wl
Cwl_0_87 word0_87 gnd C_wl
Rw1_87 word1_87 word0_87 R_wl
Cwl_1_87 word1_87 gnd C_wl
Rw2_87 word2_87 word1_87 R_wl
Cwl_2_87 word2_87 gnd C_wl
Rw3_87 word3_87 word2_87 R_wl
Cwl_3_87 word3_87 gnd C_wl
Rw4_87 word4_87 word3_87 R_wl
Cwl_4_87 word4_87 gnd C_wl
Rw5_87 word5_87 word4_87 R_wl
Cwl_5_87 word5_87 gnd C_wl
Rw6_87 word6_87 word5_87 R_wl
Cwl_6_87 word6_87 gnd C_wl
Rw7_87 word7_87 word6_87 R_wl
Cwl_7_87 word7_87 gnd C_wl
Rw8_87 word8_87 word7_87 R_wl
Cwl_8_87 word8_87 gnd C_wl
Rw9_87 word9_87 word8_87 R_wl
Cwl_9_87 word9_87 gnd C_wl
Rw10_87 word10_87 word9_87 R_wl
Cwl_10_87 word10_87 gnd C_wl
Rw11_87 word11_87 word10_87 R_wl
Cwl_11_87 word11_87 gnd C_wl
Rw12_87 word12_87 word11_87 R_wl
Cwl_12_87 word12_87 gnd C_wl
Rw13_87 word13_87 word12_87 R_wl
Cwl_13_87 word13_87 gnd C_wl
Rw14_87 word14_87 word13_87 R_wl
Cwl_14_87 word14_87 gnd C_wl
Rw15_87 word15_87 word14_87 R_wl
Cwl_15_87 word15_87 gnd C_wl
Rw16_87 word16_87 word15_87 R_wl
Cwl_16_87 word16_87 gnd C_wl
Rw17_87 word17_87 word16_87 R_wl
Cwl_17_87 word17_87 gnd C_wl
Rw18_87 word18_87 word17_87 R_wl
Cwl_18_87 word18_87 gnd C_wl
Rw19_87 word19_87 word18_87 R_wl
Cwl_19_87 word19_87 gnd C_wl
Rw20_87 word20_87 word19_87 R_wl
Cwl_20_87 word20_87 gnd C_wl
Rw21_87 word21_87 word20_87 R_wl
Cwl_21_87 word21_87 gnd C_wl
Rw22_87 word22_87 word21_87 R_wl
Cwl_22_87 word22_87 gnd C_wl
Rw23_87 word23_87 word22_87 R_wl
Cwl_23_87 word23_87 gnd C_wl
Rw24_87 word24_87 word23_87 R_wl
Cwl_24_87 word24_87 gnd C_wl
Rw25_87 word25_87 word24_87 R_wl
Cwl_25_87 word25_87 gnd C_wl
Rw26_87 word26_87 word25_87 R_wl
Cwl_26_87 word26_87 gnd C_wl
Rw27_87 word27_87 word26_87 R_wl
Cwl_27_87 word27_87 gnd C_wl
Rw28_87 word28_87 word27_87 R_wl
Cwl_28_87 word28_87 gnd C_wl
Rw29_87 word29_87 word28_87 R_wl
Cwl_29_87 word29_87 gnd C_wl
Rw30_87 word30_87 word29_87 R_wl
Cwl_30_87 word30_87 gnd C_wl
Rw31_87 word31_87 word30_87 R_wl
Cwl_31_87 word31_87 gnd C_wl
Rw32_87 word32_87 word31_87 R_wl
Cwl_32_87 word32_87 gnd C_wl
Rw33_87 word33_87 word32_87 R_wl
Cwl_33_87 word33_87 gnd C_wl
Rw34_87 word34_87 word33_87 R_wl
Cwl_34_87 word34_87 gnd C_wl
Rw35_87 word35_87 word34_87 R_wl
Cwl_35_87 word35_87 gnd C_wl
Rw36_87 word36_87 word35_87 R_wl
Cwl_36_87 word36_87 gnd C_wl
Rw37_87 word37_87 word36_87 R_wl
Cwl_37_87 word37_87 gnd C_wl
Rw38_87 word38_87 word37_87 R_wl
Cwl_38_87 word38_87 gnd C_wl
Rw39_87 word39_87 word38_87 R_wl
Cwl_39_87 word39_87 gnd C_wl
Rw40_87 word40_87 word39_87 R_wl
Cwl_40_87 word40_87 gnd C_wl
Rw41_87 word41_87 word40_87 R_wl
Cwl_41_87 word41_87 gnd C_wl
Rw42_87 word42_87 word41_87 R_wl
Cwl_42_87 word42_87 gnd C_wl
Rw43_87 word43_87 word42_87 R_wl
Cwl_43_87 word43_87 gnd C_wl
Rw44_87 word44_87 word43_87 R_wl
Cwl_44_87 word44_87 gnd C_wl
Rw45_87 word45_87 word44_87 R_wl
Cwl_45_87 word45_87 gnd C_wl
Rw46_87 word46_87 word45_87 R_wl
Cwl_46_87 word46_87 gnd C_wl
Rw47_87 word47_87 word46_87 R_wl
Cwl_47_87 word47_87 gnd C_wl
Rw48_87 word48_87 word47_87 R_wl
Cwl_48_87 word48_87 gnd C_wl
Rw49_87 word49_87 word48_87 R_wl
Cwl_49_87 word49_87 gnd C_wl
Rw50_87 word50_87 word49_87 R_wl
Cwl_50_87 word50_87 gnd C_wl
Rw51_87 word51_87 word50_87 R_wl
Cwl_51_87 word51_87 gnd C_wl
Rw52_87 word52_87 word51_87 R_wl
Cwl_52_87 word52_87 gnd C_wl
Rw53_87 word53_87 word52_87 R_wl
Cwl_53_87 word53_87 gnd C_wl
Rw54_87 word54_87 word53_87 R_wl
Cwl_54_87 word54_87 gnd C_wl
Rw55_87 word55_87 word54_87 R_wl
Cwl_55_87 word55_87 gnd C_wl
Rw56_87 word56_87 word55_87 R_wl
Cwl_56_87 word56_87 gnd C_wl
Rw57_87 word57_87 word56_87 R_wl
Cwl_57_87 word57_87 gnd C_wl
Rw58_87 word58_87 word57_87 R_wl
Cwl_58_87 word58_87 gnd C_wl
Rw59_87 word59_87 word58_87 R_wl
Cwl_59_87 word59_87 gnd C_wl
Rw60_87 word60_87 word59_87 R_wl
Cwl_60_87 word60_87 gnd C_wl
Rw61_87 word61_87 word60_87 R_wl
Cwl_61_87 word61_87 gnd C_wl
Rw62_87 word62_87 word61_87 R_wl
Cwl_62_87 word62_87 gnd C_wl
Rw63_87 word63_87 word62_87 R_wl
Cwl_63_87 word63_87 gnd C_wl
Rw64_87 word64_87 word63_87 R_wl
Cwl_64_87 word64_87 gnd C_wl
Rw65_87 word65_87 word64_87 R_wl
Cwl_65_87 word65_87 gnd C_wl
Rw66_87 word66_87 word65_87 R_wl
Cwl_66_87 word66_87 gnd C_wl
Rw67_87 word67_87 word66_87 R_wl
Cwl_67_87 word67_87 gnd C_wl
Rw68_87 word68_87 word67_87 R_wl
Cwl_68_87 word68_87 gnd C_wl
Rw69_87 word69_87 word68_87 R_wl
Cwl_69_87 word69_87 gnd C_wl
Rw70_87 word70_87 word69_87 R_wl
Cwl_70_87 word70_87 gnd C_wl
Rw71_87 word71_87 word70_87 R_wl
Cwl_71_87 word71_87 gnd C_wl
Rw72_87 word72_87 word71_87 R_wl
Cwl_72_87 word72_87 gnd C_wl
Rw73_87 word73_87 word72_87 R_wl
Cwl_73_87 word73_87 gnd C_wl
Rw74_87 word74_87 word73_87 R_wl
Cwl_74_87 word74_87 gnd C_wl
Rw75_87 word75_87 word74_87 R_wl
Cwl_75_87 word75_87 gnd C_wl
Rw76_87 word76_87 word75_87 R_wl
Cwl_76_87 word76_87 gnd C_wl
Rw77_87 word77_87 word76_87 R_wl
Cwl_77_87 word77_87 gnd C_wl
Rw78_87 word78_87 word77_87 R_wl
Cwl_78_87 word78_87 gnd C_wl
Rw79_87 word79_87 word78_87 R_wl
Cwl_79_87 word79_87 gnd C_wl
Rw80_87 word80_87 word79_87 R_wl
Cwl_80_87 word80_87 gnd C_wl
Rw81_87 word81_87 word80_87 R_wl
Cwl_81_87 word81_87 gnd C_wl
Rw82_87 word82_87 word81_87 R_wl
Cwl_82_87 word82_87 gnd C_wl
Rw83_87 word83_87 word82_87 R_wl
Cwl_83_87 word83_87 gnd C_wl
Rw84_87 word84_87 word83_87 R_wl
Cwl_84_87 word84_87 gnd C_wl
Rw85_87 word85_87 word84_87 R_wl
Cwl_85_87 word85_87 gnd C_wl
Rw86_87 word86_87 word85_87 R_wl
Cwl_86_87 word86_87 gnd C_wl
Rw87_87 word87_87 word86_87 R_wl
Cwl_87_87 word87_87 gnd C_wl
Rw88_87 word88_87 word87_87 R_wl
Cwl_88_87 word88_87 gnd C_wl
Rw89_87 word89_87 word88_87 R_wl
Cwl_89_87 word89_87 gnd C_wl
Rw90_87 word90_87 word89_87 R_wl
Cwl_90_87 word90_87 gnd C_wl
Rw91_87 word91_87 word90_87 R_wl
Cwl_91_87 word91_87 gnd C_wl
Rw92_87 word92_87 word91_87 R_wl
Cwl_92_87 word92_87 gnd C_wl
Rw93_87 word93_87 word92_87 R_wl
Cwl_93_87 word93_87 gnd C_wl
Rw94_87 word94_87 word93_87 R_wl
Cwl_94_87 word94_87 gnd C_wl
Rw95_87 word95_87 word94_87 R_wl
Cwl_95_87 word95_87 gnd C_wl
Rw96_87 word96_87 word95_87 R_wl
Cwl_96_87 word96_87 gnd C_wl
Rw97_87 word97_87 word96_87 R_wl
Cwl_97_87 word97_87 gnd C_wl
Rw98_87 word98_87 word97_87 R_wl
Cwl_98_87 word98_87 gnd C_wl
Rw99_87 word99_87 word98_87 R_wl
Cwl_99_87 word99_87 gnd C_wl
Vwl_88 word_88 0 0
Rw0_88 word_88 word0_88 R_wl
Cwl_0_88 word0_88 gnd C_wl
Rw1_88 word1_88 word0_88 R_wl
Cwl_1_88 word1_88 gnd C_wl
Rw2_88 word2_88 word1_88 R_wl
Cwl_2_88 word2_88 gnd C_wl
Rw3_88 word3_88 word2_88 R_wl
Cwl_3_88 word3_88 gnd C_wl
Rw4_88 word4_88 word3_88 R_wl
Cwl_4_88 word4_88 gnd C_wl
Rw5_88 word5_88 word4_88 R_wl
Cwl_5_88 word5_88 gnd C_wl
Rw6_88 word6_88 word5_88 R_wl
Cwl_6_88 word6_88 gnd C_wl
Rw7_88 word7_88 word6_88 R_wl
Cwl_7_88 word7_88 gnd C_wl
Rw8_88 word8_88 word7_88 R_wl
Cwl_8_88 word8_88 gnd C_wl
Rw9_88 word9_88 word8_88 R_wl
Cwl_9_88 word9_88 gnd C_wl
Rw10_88 word10_88 word9_88 R_wl
Cwl_10_88 word10_88 gnd C_wl
Rw11_88 word11_88 word10_88 R_wl
Cwl_11_88 word11_88 gnd C_wl
Rw12_88 word12_88 word11_88 R_wl
Cwl_12_88 word12_88 gnd C_wl
Rw13_88 word13_88 word12_88 R_wl
Cwl_13_88 word13_88 gnd C_wl
Rw14_88 word14_88 word13_88 R_wl
Cwl_14_88 word14_88 gnd C_wl
Rw15_88 word15_88 word14_88 R_wl
Cwl_15_88 word15_88 gnd C_wl
Rw16_88 word16_88 word15_88 R_wl
Cwl_16_88 word16_88 gnd C_wl
Rw17_88 word17_88 word16_88 R_wl
Cwl_17_88 word17_88 gnd C_wl
Rw18_88 word18_88 word17_88 R_wl
Cwl_18_88 word18_88 gnd C_wl
Rw19_88 word19_88 word18_88 R_wl
Cwl_19_88 word19_88 gnd C_wl
Rw20_88 word20_88 word19_88 R_wl
Cwl_20_88 word20_88 gnd C_wl
Rw21_88 word21_88 word20_88 R_wl
Cwl_21_88 word21_88 gnd C_wl
Rw22_88 word22_88 word21_88 R_wl
Cwl_22_88 word22_88 gnd C_wl
Rw23_88 word23_88 word22_88 R_wl
Cwl_23_88 word23_88 gnd C_wl
Rw24_88 word24_88 word23_88 R_wl
Cwl_24_88 word24_88 gnd C_wl
Rw25_88 word25_88 word24_88 R_wl
Cwl_25_88 word25_88 gnd C_wl
Rw26_88 word26_88 word25_88 R_wl
Cwl_26_88 word26_88 gnd C_wl
Rw27_88 word27_88 word26_88 R_wl
Cwl_27_88 word27_88 gnd C_wl
Rw28_88 word28_88 word27_88 R_wl
Cwl_28_88 word28_88 gnd C_wl
Rw29_88 word29_88 word28_88 R_wl
Cwl_29_88 word29_88 gnd C_wl
Rw30_88 word30_88 word29_88 R_wl
Cwl_30_88 word30_88 gnd C_wl
Rw31_88 word31_88 word30_88 R_wl
Cwl_31_88 word31_88 gnd C_wl
Rw32_88 word32_88 word31_88 R_wl
Cwl_32_88 word32_88 gnd C_wl
Rw33_88 word33_88 word32_88 R_wl
Cwl_33_88 word33_88 gnd C_wl
Rw34_88 word34_88 word33_88 R_wl
Cwl_34_88 word34_88 gnd C_wl
Rw35_88 word35_88 word34_88 R_wl
Cwl_35_88 word35_88 gnd C_wl
Rw36_88 word36_88 word35_88 R_wl
Cwl_36_88 word36_88 gnd C_wl
Rw37_88 word37_88 word36_88 R_wl
Cwl_37_88 word37_88 gnd C_wl
Rw38_88 word38_88 word37_88 R_wl
Cwl_38_88 word38_88 gnd C_wl
Rw39_88 word39_88 word38_88 R_wl
Cwl_39_88 word39_88 gnd C_wl
Rw40_88 word40_88 word39_88 R_wl
Cwl_40_88 word40_88 gnd C_wl
Rw41_88 word41_88 word40_88 R_wl
Cwl_41_88 word41_88 gnd C_wl
Rw42_88 word42_88 word41_88 R_wl
Cwl_42_88 word42_88 gnd C_wl
Rw43_88 word43_88 word42_88 R_wl
Cwl_43_88 word43_88 gnd C_wl
Rw44_88 word44_88 word43_88 R_wl
Cwl_44_88 word44_88 gnd C_wl
Rw45_88 word45_88 word44_88 R_wl
Cwl_45_88 word45_88 gnd C_wl
Rw46_88 word46_88 word45_88 R_wl
Cwl_46_88 word46_88 gnd C_wl
Rw47_88 word47_88 word46_88 R_wl
Cwl_47_88 word47_88 gnd C_wl
Rw48_88 word48_88 word47_88 R_wl
Cwl_48_88 word48_88 gnd C_wl
Rw49_88 word49_88 word48_88 R_wl
Cwl_49_88 word49_88 gnd C_wl
Rw50_88 word50_88 word49_88 R_wl
Cwl_50_88 word50_88 gnd C_wl
Rw51_88 word51_88 word50_88 R_wl
Cwl_51_88 word51_88 gnd C_wl
Rw52_88 word52_88 word51_88 R_wl
Cwl_52_88 word52_88 gnd C_wl
Rw53_88 word53_88 word52_88 R_wl
Cwl_53_88 word53_88 gnd C_wl
Rw54_88 word54_88 word53_88 R_wl
Cwl_54_88 word54_88 gnd C_wl
Rw55_88 word55_88 word54_88 R_wl
Cwl_55_88 word55_88 gnd C_wl
Rw56_88 word56_88 word55_88 R_wl
Cwl_56_88 word56_88 gnd C_wl
Rw57_88 word57_88 word56_88 R_wl
Cwl_57_88 word57_88 gnd C_wl
Rw58_88 word58_88 word57_88 R_wl
Cwl_58_88 word58_88 gnd C_wl
Rw59_88 word59_88 word58_88 R_wl
Cwl_59_88 word59_88 gnd C_wl
Rw60_88 word60_88 word59_88 R_wl
Cwl_60_88 word60_88 gnd C_wl
Rw61_88 word61_88 word60_88 R_wl
Cwl_61_88 word61_88 gnd C_wl
Rw62_88 word62_88 word61_88 R_wl
Cwl_62_88 word62_88 gnd C_wl
Rw63_88 word63_88 word62_88 R_wl
Cwl_63_88 word63_88 gnd C_wl
Rw64_88 word64_88 word63_88 R_wl
Cwl_64_88 word64_88 gnd C_wl
Rw65_88 word65_88 word64_88 R_wl
Cwl_65_88 word65_88 gnd C_wl
Rw66_88 word66_88 word65_88 R_wl
Cwl_66_88 word66_88 gnd C_wl
Rw67_88 word67_88 word66_88 R_wl
Cwl_67_88 word67_88 gnd C_wl
Rw68_88 word68_88 word67_88 R_wl
Cwl_68_88 word68_88 gnd C_wl
Rw69_88 word69_88 word68_88 R_wl
Cwl_69_88 word69_88 gnd C_wl
Rw70_88 word70_88 word69_88 R_wl
Cwl_70_88 word70_88 gnd C_wl
Rw71_88 word71_88 word70_88 R_wl
Cwl_71_88 word71_88 gnd C_wl
Rw72_88 word72_88 word71_88 R_wl
Cwl_72_88 word72_88 gnd C_wl
Rw73_88 word73_88 word72_88 R_wl
Cwl_73_88 word73_88 gnd C_wl
Rw74_88 word74_88 word73_88 R_wl
Cwl_74_88 word74_88 gnd C_wl
Rw75_88 word75_88 word74_88 R_wl
Cwl_75_88 word75_88 gnd C_wl
Rw76_88 word76_88 word75_88 R_wl
Cwl_76_88 word76_88 gnd C_wl
Rw77_88 word77_88 word76_88 R_wl
Cwl_77_88 word77_88 gnd C_wl
Rw78_88 word78_88 word77_88 R_wl
Cwl_78_88 word78_88 gnd C_wl
Rw79_88 word79_88 word78_88 R_wl
Cwl_79_88 word79_88 gnd C_wl
Rw80_88 word80_88 word79_88 R_wl
Cwl_80_88 word80_88 gnd C_wl
Rw81_88 word81_88 word80_88 R_wl
Cwl_81_88 word81_88 gnd C_wl
Rw82_88 word82_88 word81_88 R_wl
Cwl_82_88 word82_88 gnd C_wl
Rw83_88 word83_88 word82_88 R_wl
Cwl_83_88 word83_88 gnd C_wl
Rw84_88 word84_88 word83_88 R_wl
Cwl_84_88 word84_88 gnd C_wl
Rw85_88 word85_88 word84_88 R_wl
Cwl_85_88 word85_88 gnd C_wl
Rw86_88 word86_88 word85_88 R_wl
Cwl_86_88 word86_88 gnd C_wl
Rw87_88 word87_88 word86_88 R_wl
Cwl_87_88 word87_88 gnd C_wl
Rw88_88 word88_88 word87_88 R_wl
Cwl_88_88 word88_88 gnd C_wl
Rw89_88 word89_88 word88_88 R_wl
Cwl_89_88 word89_88 gnd C_wl
Rw90_88 word90_88 word89_88 R_wl
Cwl_90_88 word90_88 gnd C_wl
Rw91_88 word91_88 word90_88 R_wl
Cwl_91_88 word91_88 gnd C_wl
Rw92_88 word92_88 word91_88 R_wl
Cwl_92_88 word92_88 gnd C_wl
Rw93_88 word93_88 word92_88 R_wl
Cwl_93_88 word93_88 gnd C_wl
Rw94_88 word94_88 word93_88 R_wl
Cwl_94_88 word94_88 gnd C_wl
Rw95_88 word95_88 word94_88 R_wl
Cwl_95_88 word95_88 gnd C_wl
Rw96_88 word96_88 word95_88 R_wl
Cwl_96_88 word96_88 gnd C_wl
Rw97_88 word97_88 word96_88 R_wl
Cwl_97_88 word97_88 gnd C_wl
Rw98_88 word98_88 word97_88 R_wl
Cwl_98_88 word98_88 gnd C_wl
Rw99_88 word99_88 word98_88 R_wl
Cwl_99_88 word99_88 gnd C_wl
Vwl_89 word_89 0 0
Rw0_89 word_89 word0_89 R_wl
Cwl_0_89 word0_89 gnd C_wl
Rw1_89 word1_89 word0_89 R_wl
Cwl_1_89 word1_89 gnd C_wl
Rw2_89 word2_89 word1_89 R_wl
Cwl_2_89 word2_89 gnd C_wl
Rw3_89 word3_89 word2_89 R_wl
Cwl_3_89 word3_89 gnd C_wl
Rw4_89 word4_89 word3_89 R_wl
Cwl_4_89 word4_89 gnd C_wl
Rw5_89 word5_89 word4_89 R_wl
Cwl_5_89 word5_89 gnd C_wl
Rw6_89 word6_89 word5_89 R_wl
Cwl_6_89 word6_89 gnd C_wl
Rw7_89 word7_89 word6_89 R_wl
Cwl_7_89 word7_89 gnd C_wl
Rw8_89 word8_89 word7_89 R_wl
Cwl_8_89 word8_89 gnd C_wl
Rw9_89 word9_89 word8_89 R_wl
Cwl_9_89 word9_89 gnd C_wl
Rw10_89 word10_89 word9_89 R_wl
Cwl_10_89 word10_89 gnd C_wl
Rw11_89 word11_89 word10_89 R_wl
Cwl_11_89 word11_89 gnd C_wl
Rw12_89 word12_89 word11_89 R_wl
Cwl_12_89 word12_89 gnd C_wl
Rw13_89 word13_89 word12_89 R_wl
Cwl_13_89 word13_89 gnd C_wl
Rw14_89 word14_89 word13_89 R_wl
Cwl_14_89 word14_89 gnd C_wl
Rw15_89 word15_89 word14_89 R_wl
Cwl_15_89 word15_89 gnd C_wl
Rw16_89 word16_89 word15_89 R_wl
Cwl_16_89 word16_89 gnd C_wl
Rw17_89 word17_89 word16_89 R_wl
Cwl_17_89 word17_89 gnd C_wl
Rw18_89 word18_89 word17_89 R_wl
Cwl_18_89 word18_89 gnd C_wl
Rw19_89 word19_89 word18_89 R_wl
Cwl_19_89 word19_89 gnd C_wl
Rw20_89 word20_89 word19_89 R_wl
Cwl_20_89 word20_89 gnd C_wl
Rw21_89 word21_89 word20_89 R_wl
Cwl_21_89 word21_89 gnd C_wl
Rw22_89 word22_89 word21_89 R_wl
Cwl_22_89 word22_89 gnd C_wl
Rw23_89 word23_89 word22_89 R_wl
Cwl_23_89 word23_89 gnd C_wl
Rw24_89 word24_89 word23_89 R_wl
Cwl_24_89 word24_89 gnd C_wl
Rw25_89 word25_89 word24_89 R_wl
Cwl_25_89 word25_89 gnd C_wl
Rw26_89 word26_89 word25_89 R_wl
Cwl_26_89 word26_89 gnd C_wl
Rw27_89 word27_89 word26_89 R_wl
Cwl_27_89 word27_89 gnd C_wl
Rw28_89 word28_89 word27_89 R_wl
Cwl_28_89 word28_89 gnd C_wl
Rw29_89 word29_89 word28_89 R_wl
Cwl_29_89 word29_89 gnd C_wl
Rw30_89 word30_89 word29_89 R_wl
Cwl_30_89 word30_89 gnd C_wl
Rw31_89 word31_89 word30_89 R_wl
Cwl_31_89 word31_89 gnd C_wl
Rw32_89 word32_89 word31_89 R_wl
Cwl_32_89 word32_89 gnd C_wl
Rw33_89 word33_89 word32_89 R_wl
Cwl_33_89 word33_89 gnd C_wl
Rw34_89 word34_89 word33_89 R_wl
Cwl_34_89 word34_89 gnd C_wl
Rw35_89 word35_89 word34_89 R_wl
Cwl_35_89 word35_89 gnd C_wl
Rw36_89 word36_89 word35_89 R_wl
Cwl_36_89 word36_89 gnd C_wl
Rw37_89 word37_89 word36_89 R_wl
Cwl_37_89 word37_89 gnd C_wl
Rw38_89 word38_89 word37_89 R_wl
Cwl_38_89 word38_89 gnd C_wl
Rw39_89 word39_89 word38_89 R_wl
Cwl_39_89 word39_89 gnd C_wl
Rw40_89 word40_89 word39_89 R_wl
Cwl_40_89 word40_89 gnd C_wl
Rw41_89 word41_89 word40_89 R_wl
Cwl_41_89 word41_89 gnd C_wl
Rw42_89 word42_89 word41_89 R_wl
Cwl_42_89 word42_89 gnd C_wl
Rw43_89 word43_89 word42_89 R_wl
Cwl_43_89 word43_89 gnd C_wl
Rw44_89 word44_89 word43_89 R_wl
Cwl_44_89 word44_89 gnd C_wl
Rw45_89 word45_89 word44_89 R_wl
Cwl_45_89 word45_89 gnd C_wl
Rw46_89 word46_89 word45_89 R_wl
Cwl_46_89 word46_89 gnd C_wl
Rw47_89 word47_89 word46_89 R_wl
Cwl_47_89 word47_89 gnd C_wl
Rw48_89 word48_89 word47_89 R_wl
Cwl_48_89 word48_89 gnd C_wl
Rw49_89 word49_89 word48_89 R_wl
Cwl_49_89 word49_89 gnd C_wl
Rw50_89 word50_89 word49_89 R_wl
Cwl_50_89 word50_89 gnd C_wl
Rw51_89 word51_89 word50_89 R_wl
Cwl_51_89 word51_89 gnd C_wl
Rw52_89 word52_89 word51_89 R_wl
Cwl_52_89 word52_89 gnd C_wl
Rw53_89 word53_89 word52_89 R_wl
Cwl_53_89 word53_89 gnd C_wl
Rw54_89 word54_89 word53_89 R_wl
Cwl_54_89 word54_89 gnd C_wl
Rw55_89 word55_89 word54_89 R_wl
Cwl_55_89 word55_89 gnd C_wl
Rw56_89 word56_89 word55_89 R_wl
Cwl_56_89 word56_89 gnd C_wl
Rw57_89 word57_89 word56_89 R_wl
Cwl_57_89 word57_89 gnd C_wl
Rw58_89 word58_89 word57_89 R_wl
Cwl_58_89 word58_89 gnd C_wl
Rw59_89 word59_89 word58_89 R_wl
Cwl_59_89 word59_89 gnd C_wl
Rw60_89 word60_89 word59_89 R_wl
Cwl_60_89 word60_89 gnd C_wl
Rw61_89 word61_89 word60_89 R_wl
Cwl_61_89 word61_89 gnd C_wl
Rw62_89 word62_89 word61_89 R_wl
Cwl_62_89 word62_89 gnd C_wl
Rw63_89 word63_89 word62_89 R_wl
Cwl_63_89 word63_89 gnd C_wl
Rw64_89 word64_89 word63_89 R_wl
Cwl_64_89 word64_89 gnd C_wl
Rw65_89 word65_89 word64_89 R_wl
Cwl_65_89 word65_89 gnd C_wl
Rw66_89 word66_89 word65_89 R_wl
Cwl_66_89 word66_89 gnd C_wl
Rw67_89 word67_89 word66_89 R_wl
Cwl_67_89 word67_89 gnd C_wl
Rw68_89 word68_89 word67_89 R_wl
Cwl_68_89 word68_89 gnd C_wl
Rw69_89 word69_89 word68_89 R_wl
Cwl_69_89 word69_89 gnd C_wl
Rw70_89 word70_89 word69_89 R_wl
Cwl_70_89 word70_89 gnd C_wl
Rw71_89 word71_89 word70_89 R_wl
Cwl_71_89 word71_89 gnd C_wl
Rw72_89 word72_89 word71_89 R_wl
Cwl_72_89 word72_89 gnd C_wl
Rw73_89 word73_89 word72_89 R_wl
Cwl_73_89 word73_89 gnd C_wl
Rw74_89 word74_89 word73_89 R_wl
Cwl_74_89 word74_89 gnd C_wl
Rw75_89 word75_89 word74_89 R_wl
Cwl_75_89 word75_89 gnd C_wl
Rw76_89 word76_89 word75_89 R_wl
Cwl_76_89 word76_89 gnd C_wl
Rw77_89 word77_89 word76_89 R_wl
Cwl_77_89 word77_89 gnd C_wl
Rw78_89 word78_89 word77_89 R_wl
Cwl_78_89 word78_89 gnd C_wl
Rw79_89 word79_89 word78_89 R_wl
Cwl_79_89 word79_89 gnd C_wl
Rw80_89 word80_89 word79_89 R_wl
Cwl_80_89 word80_89 gnd C_wl
Rw81_89 word81_89 word80_89 R_wl
Cwl_81_89 word81_89 gnd C_wl
Rw82_89 word82_89 word81_89 R_wl
Cwl_82_89 word82_89 gnd C_wl
Rw83_89 word83_89 word82_89 R_wl
Cwl_83_89 word83_89 gnd C_wl
Rw84_89 word84_89 word83_89 R_wl
Cwl_84_89 word84_89 gnd C_wl
Rw85_89 word85_89 word84_89 R_wl
Cwl_85_89 word85_89 gnd C_wl
Rw86_89 word86_89 word85_89 R_wl
Cwl_86_89 word86_89 gnd C_wl
Rw87_89 word87_89 word86_89 R_wl
Cwl_87_89 word87_89 gnd C_wl
Rw88_89 word88_89 word87_89 R_wl
Cwl_88_89 word88_89 gnd C_wl
Rw89_89 word89_89 word88_89 R_wl
Cwl_89_89 word89_89 gnd C_wl
Rw90_89 word90_89 word89_89 R_wl
Cwl_90_89 word90_89 gnd C_wl
Rw91_89 word91_89 word90_89 R_wl
Cwl_91_89 word91_89 gnd C_wl
Rw92_89 word92_89 word91_89 R_wl
Cwl_92_89 word92_89 gnd C_wl
Rw93_89 word93_89 word92_89 R_wl
Cwl_93_89 word93_89 gnd C_wl
Rw94_89 word94_89 word93_89 R_wl
Cwl_94_89 word94_89 gnd C_wl
Rw95_89 word95_89 word94_89 R_wl
Cwl_95_89 word95_89 gnd C_wl
Rw96_89 word96_89 word95_89 R_wl
Cwl_96_89 word96_89 gnd C_wl
Rw97_89 word97_89 word96_89 R_wl
Cwl_97_89 word97_89 gnd C_wl
Rw98_89 word98_89 word97_89 R_wl
Cwl_98_89 word98_89 gnd C_wl
Rw99_89 word99_89 word98_89 R_wl
Cwl_99_89 word99_89 gnd C_wl
Vwl_90 word_90 0 0
Rw0_90 word_90 word0_90 R_wl
Cwl_0_90 word0_90 gnd C_wl
Rw1_90 word1_90 word0_90 R_wl
Cwl_1_90 word1_90 gnd C_wl
Rw2_90 word2_90 word1_90 R_wl
Cwl_2_90 word2_90 gnd C_wl
Rw3_90 word3_90 word2_90 R_wl
Cwl_3_90 word3_90 gnd C_wl
Rw4_90 word4_90 word3_90 R_wl
Cwl_4_90 word4_90 gnd C_wl
Rw5_90 word5_90 word4_90 R_wl
Cwl_5_90 word5_90 gnd C_wl
Rw6_90 word6_90 word5_90 R_wl
Cwl_6_90 word6_90 gnd C_wl
Rw7_90 word7_90 word6_90 R_wl
Cwl_7_90 word7_90 gnd C_wl
Rw8_90 word8_90 word7_90 R_wl
Cwl_8_90 word8_90 gnd C_wl
Rw9_90 word9_90 word8_90 R_wl
Cwl_9_90 word9_90 gnd C_wl
Rw10_90 word10_90 word9_90 R_wl
Cwl_10_90 word10_90 gnd C_wl
Rw11_90 word11_90 word10_90 R_wl
Cwl_11_90 word11_90 gnd C_wl
Rw12_90 word12_90 word11_90 R_wl
Cwl_12_90 word12_90 gnd C_wl
Rw13_90 word13_90 word12_90 R_wl
Cwl_13_90 word13_90 gnd C_wl
Rw14_90 word14_90 word13_90 R_wl
Cwl_14_90 word14_90 gnd C_wl
Rw15_90 word15_90 word14_90 R_wl
Cwl_15_90 word15_90 gnd C_wl
Rw16_90 word16_90 word15_90 R_wl
Cwl_16_90 word16_90 gnd C_wl
Rw17_90 word17_90 word16_90 R_wl
Cwl_17_90 word17_90 gnd C_wl
Rw18_90 word18_90 word17_90 R_wl
Cwl_18_90 word18_90 gnd C_wl
Rw19_90 word19_90 word18_90 R_wl
Cwl_19_90 word19_90 gnd C_wl
Rw20_90 word20_90 word19_90 R_wl
Cwl_20_90 word20_90 gnd C_wl
Rw21_90 word21_90 word20_90 R_wl
Cwl_21_90 word21_90 gnd C_wl
Rw22_90 word22_90 word21_90 R_wl
Cwl_22_90 word22_90 gnd C_wl
Rw23_90 word23_90 word22_90 R_wl
Cwl_23_90 word23_90 gnd C_wl
Rw24_90 word24_90 word23_90 R_wl
Cwl_24_90 word24_90 gnd C_wl
Rw25_90 word25_90 word24_90 R_wl
Cwl_25_90 word25_90 gnd C_wl
Rw26_90 word26_90 word25_90 R_wl
Cwl_26_90 word26_90 gnd C_wl
Rw27_90 word27_90 word26_90 R_wl
Cwl_27_90 word27_90 gnd C_wl
Rw28_90 word28_90 word27_90 R_wl
Cwl_28_90 word28_90 gnd C_wl
Rw29_90 word29_90 word28_90 R_wl
Cwl_29_90 word29_90 gnd C_wl
Rw30_90 word30_90 word29_90 R_wl
Cwl_30_90 word30_90 gnd C_wl
Rw31_90 word31_90 word30_90 R_wl
Cwl_31_90 word31_90 gnd C_wl
Rw32_90 word32_90 word31_90 R_wl
Cwl_32_90 word32_90 gnd C_wl
Rw33_90 word33_90 word32_90 R_wl
Cwl_33_90 word33_90 gnd C_wl
Rw34_90 word34_90 word33_90 R_wl
Cwl_34_90 word34_90 gnd C_wl
Rw35_90 word35_90 word34_90 R_wl
Cwl_35_90 word35_90 gnd C_wl
Rw36_90 word36_90 word35_90 R_wl
Cwl_36_90 word36_90 gnd C_wl
Rw37_90 word37_90 word36_90 R_wl
Cwl_37_90 word37_90 gnd C_wl
Rw38_90 word38_90 word37_90 R_wl
Cwl_38_90 word38_90 gnd C_wl
Rw39_90 word39_90 word38_90 R_wl
Cwl_39_90 word39_90 gnd C_wl
Rw40_90 word40_90 word39_90 R_wl
Cwl_40_90 word40_90 gnd C_wl
Rw41_90 word41_90 word40_90 R_wl
Cwl_41_90 word41_90 gnd C_wl
Rw42_90 word42_90 word41_90 R_wl
Cwl_42_90 word42_90 gnd C_wl
Rw43_90 word43_90 word42_90 R_wl
Cwl_43_90 word43_90 gnd C_wl
Rw44_90 word44_90 word43_90 R_wl
Cwl_44_90 word44_90 gnd C_wl
Rw45_90 word45_90 word44_90 R_wl
Cwl_45_90 word45_90 gnd C_wl
Rw46_90 word46_90 word45_90 R_wl
Cwl_46_90 word46_90 gnd C_wl
Rw47_90 word47_90 word46_90 R_wl
Cwl_47_90 word47_90 gnd C_wl
Rw48_90 word48_90 word47_90 R_wl
Cwl_48_90 word48_90 gnd C_wl
Rw49_90 word49_90 word48_90 R_wl
Cwl_49_90 word49_90 gnd C_wl
Rw50_90 word50_90 word49_90 R_wl
Cwl_50_90 word50_90 gnd C_wl
Rw51_90 word51_90 word50_90 R_wl
Cwl_51_90 word51_90 gnd C_wl
Rw52_90 word52_90 word51_90 R_wl
Cwl_52_90 word52_90 gnd C_wl
Rw53_90 word53_90 word52_90 R_wl
Cwl_53_90 word53_90 gnd C_wl
Rw54_90 word54_90 word53_90 R_wl
Cwl_54_90 word54_90 gnd C_wl
Rw55_90 word55_90 word54_90 R_wl
Cwl_55_90 word55_90 gnd C_wl
Rw56_90 word56_90 word55_90 R_wl
Cwl_56_90 word56_90 gnd C_wl
Rw57_90 word57_90 word56_90 R_wl
Cwl_57_90 word57_90 gnd C_wl
Rw58_90 word58_90 word57_90 R_wl
Cwl_58_90 word58_90 gnd C_wl
Rw59_90 word59_90 word58_90 R_wl
Cwl_59_90 word59_90 gnd C_wl
Rw60_90 word60_90 word59_90 R_wl
Cwl_60_90 word60_90 gnd C_wl
Rw61_90 word61_90 word60_90 R_wl
Cwl_61_90 word61_90 gnd C_wl
Rw62_90 word62_90 word61_90 R_wl
Cwl_62_90 word62_90 gnd C_wl
Rw63_90 word63_90 word62_90 R_wl
Cwl_63_90 word63_90 gnd C_wl
Rw64_90 word64_90 word63_90 R_wl
Cwl_64_90 word64_90 gnd C_wl
Rw65_90 word65_90 word64_90 R_wl
Cwl_65_90 word65_90 gnd C_wl
Rw66_90 word66_90 word65_90 R_wl
Cwl_66_90 word66_90 gnd C_wl
Rw67_90 word67_90 word66_90 R_wl
Cwl_67_90 word67_90 gnd C_wl
Rw68_90 word68_90 word67_90 R_wl
Cwl_68_90 word68_90 gnd C_wl
Rw69_90 word69_90 word68_90 R_wl
Cwl_69_90 word69_90 gnd C_wl
Rw70_90 word70_90 word69_90 R_wl
Cwl_70_90 word70_90 gnd C_wl
Rw71_90 word71_90 word70_90 R_wl
Cwl_71_90 word71_90 gnd C_wl
Rw72_90 word72_90 word71_90 R_wl
Cwl_72_90 word72_90 gnd C_wl
Rw73_90 word73_90 word72_90 R_wl
Cwl_73_90 word73_90 gnd C_wl
Rw74_90 word74_90 word73_90 R_wl
Cwl_74_90 word74_90 gnd C_wl
Rw75_90 word75_90 word74_90 R_wl
Cwl_75_90 word75_90 gnd C_wl
Rw76_90 word76_90 word75_90 R_wl
Cwl_76_90 word76_90 gnd C_wl
Rw77_90 word77_90 word76_90 R_wl
Cwl_77_90 word77_90 gnd C_wl
Rw78_90 word78_90 word77_90 R_wl
Cwl_78_90 word78_90 gnd C_wl
Rw79_90 word79_90 word78_90 R_wl
Cwl_79_90 word79_90 gnd C_wl
Rw80_90 word80_90 word79_90 R_wl
Cwl_80_90 word80_90 gnd C_wl
Rw81_90 word81_90 word80_90 R_wl
Cwl_81_90 word81_90 gnd C_wl
Rw82_90 word82_90 word81_90 R_wl
Cwl_82_90 word82_90 gnd C_wl
Rw83_90 word83_90 word82_90 R_wl
Cwl_83_90 word83_90 gnd C_wl
Rw84_90 word84_90 word83_90 R_wl
Cwl_84_90 word84_90 gnd C_wl
Rw85_90 word85_90 word84_90 R_wl
Cwl_85_90 word85_90 gnd C_wl
Rw86_90 word86_90 word85_90 R_wl
Cwl_86_90 word86_90 gnd C_wl
Rw87_90 word87_90 word86_90 R_wl
Cwl_87_90 word87_90 gnd C_wl
Rw88_90 word88_90 word87_90 R_wl
Cwl_88_90 word88_90 gnd C_wl
Rw89_90 word89_90 word88_90 R_wl
Cwl_89_90 word89_90 gnd C_wl
Rw90_90 word90_90 word89_90 R_wl
Cwl_90_90 word90_90 gnd C_wl
Rw91_90 word91_90 word90_90 R_wl
Cwl_91_90 word91_90 gnd C_wl
Rw92_90 word92_90 word91_90 R_wl
Cwl_92_90 word92_90 gnd C_wl
Rw93_90 word93_90 word92_90 R_wl
Cwl_93_90 word93_90 gnd C_wl
Rw94_90 word94_90 word93_90 R_wl
Cwl_94_90 word94_90 gnd C_wl
Rw95_90 word95_90 word94_90 R_wl
Cwl_95_90 word95_90 gnd C_wl
Rw96_90 word96_90 word95_90 R_wl
Cwl_96_90 word96_90 gnd C_wl
Rw97_90 word97_90 word96_90 R_wl
Cwl_97_90 word97_90 gnd C_wl
Rw98_90 word98_90 word97_90 R_wl
Cwl_98_90 word98_90 gnd C_wl
Rw99_90 word99_90 word98_90 R_wl
Cwl_99_90 word99_90 gnd C_wl
Vwl_91 word_91 0 0
Rw0_91 word_91 word0_91 R_wl
Cwl_0_91 word0_91 gnd C_wl
Rw1_91 word1_91 word0_91 R_wl
Cwl_1_91 word1_91 gnd C_wl
Rw2_91 word2_91 word1_91 R_wl
Cwl_2_91 word2_91 gnd C_wl
Rw3_91 word3_91 word2_91 R_wl
Cwl_3_91 word3_91 gnd C_wl
Rw4_91 word4_91 word3_91 R_wl
Cwl_4_91 word4_91 gnd C_wl
Rw5_91 word5_91 word4_91 R_wl
Cwl_5_91 word5_91 gnd C_wl
Rw6_91 word6_91 word5_91 R_wl
Cwl_6_91 word6_91 gnd C_wl
Rw7_91 word7_91 word6_91 R_wl
Cwl_7_91 word7_91 gnd C_wl
Rw8_91 word8_91 word7_91 R_wl
Cwl_8_91 word8_91 gnd C_wl
Rw9_91 word9_91 word8_91 R_wl
Cwl_9_91 word9_91 gnd C_wl
Rw10_91 word10_91 word9_91 R_wl
Cwl_10_91 word10_91 gnd C_wl
Rw11_91 word11_91 word10_91 R_wl
Cwl_11_91 word11_91 gnd C_wl
Rw12_91 word12_91 word11_91 R_wl
Cwl_12_91 word12_91 gnd C_wl
Rw13_91 word13_91 word12_91 R_wl
Cwl_13_91 word13_91 gnd C_wl
Rw14_91 word14_91 word13_91 R_wl
Cwl_14_91 word14_91 gnd C_wl
Rw15_91 word15_91 word14_91 R_wl
Cwl_15_91 word15_91 gnd C_wl
Rw16_91 word16_91 word15_91 R_wl
Cwl_16_91 word16_91 gnd C_wl
Rw17_91 word17_91 word16_91 R_wl
Cwl_17_91 word17_91 gnd C_wl
Rw18_91 word18_91 word17_91 R_wl
Cwl_18_91 word18_91 gnd C_wl
Rw19_91 word19_91 word18_91 R_wl
Cwl_19_91 word19_91 gnd C_wl
Rw20_91 word20_91 word19_91 R_wl
Cwl_20_91 word20_91 gnd C_wl
Rw21_91 word21_91 word20_91 R_wl
Cwl_21_91 word21_91 gnd C_wl
Rw22_91 word22_91 word21_91 R_wl
Cwl_22_91 word22_91 gnd C_wl
Rw23_91 word23_91 word22_91 R_wl
Cwl_23_91 word23_91 gnd C_wl
Rw24_91 word24_91 word23_91 R_wl
Cwl_24_91 word24_91 gnd C_wl
Rw25_91 word25_91 word24_91 R_wl
Cwl_25_91 word25_91 gnd C_wl
Rw26_91 word26_91 word25_91 R_wl
Cwl_26_91 word26_91 gnd C_wl
Rw27_91 word27_91 word26_91 R_wl
Cwl_27_91 word27_91 gnd C_wl
Rw28_91 word28_91 word27_91 R_wl
Cwl_28_91 word28_91 gnd C_wl
Rw29_91 word29_91 word28_91 R_wl
Cwl_29_91 word29_91 gnd C_wl
Rw30_91 word30_91 word29_91 R_wl
Cwl_30_91 word30_91 gnd C_wl
Rw31_91 word31_91 word30_91 R_wl
Cwl_31_91 word31_91 gnd C_wl
Rw32_91 word32_91 word31_91 R_wl
Cwl_32_91 word32_91 gnd C_wl
Rw33_91 word33_91 word32_91 R_wl
Cwl_33_91 word33_91 gnd C_wl
Rw34_91 word34_91 word33_91 R_wl
Cwl_34_91 word34_91 gnd C_wl
Rw35_91 word35_91 word34_91 R_wl
Cwl_35_91 word35_91 gnd C_wl
Rw36_91 word36_91 word35_91 R_wl
Cwl_36_91 word36_91 gnd C_wl
Rw37_91 word37_91 word36_91 R_wl
Cwl_37_91 word37_91 gnd C_wl
Rw38_91 word38_91 word37_91 R_wl
Cwl_38_91 word38_91 gnd C_wl
Rw39_91 word39_91 word38_91 R_wl
Cwl_39_91 word39_91 gnd C_wl
Rw40_91 word40_91 word39_91 R_wl
Cwl_40_91 word40_91 gnd C_wl
Rw41_91 word41_91 word40_91 R_wl
Cwl_41_91 word41_91 gnd C_wl
Rw42_91 word42_91 word41_91 R_wl
Cwl_42_91 word42_91 gnd C_wl
Rw43_91 word43_91 word42_91 R_wl
Cwl_43_91 word43_91 gnd C_wl
Rw44_91 word44_91 word43_91 R_wl
Cwl_44_91 word44_91 gnd C_wl
Rw45_91 word45_91 word44_91 R_wl
Cwl_45_91 word45_91 gnd C_wl
Rw46_91 word46_91 word45_91 R_wl
Cwl_46_91 word46_91 gnd C_wl
Rw47_91 word47_91 word46_91 R_wl
Cwl_47_91 word47_91 gnd C_wl
Rw48_91 word48_91 word47_91 R_wl
Cwl_48_91 word48_91 gnd C_wl
Rw49_91 word49_91 word48_91 R_wl
Cwl_49_91 word49_91 gnd C_wl
Rw50_91 word50_91 word49_91 R_wl
Cwl_50_91 word50_91 gnd C_wl
Rw51_91 word51_91 word50_91 R_wl
Cwl_51_91 word51_91 gnd C_wl
Rw52_91 word52_91 word51_91 R_wl
Cwl_52_91 word52_91 gnd C_wl
Rw53_91 word53_91 word52_91 R_wl
Cwl_53_91 word53_91 gnd C_wl
Rw54_91 word54_91 word53_91 R_wl
Cwl_54_91 word54_91 gnd C_wl
Rw55_91 word55_91 word54_91 R_wl
Cwl_55_91 word55_91 gnd C_wl
Rw56_91 word56_91 word55_91 R_wl
Cwl_56_91 word56_91 gnd C_wl
Rw57_91 word57_91 word56_91 R_wl
Cwl_57_91 word57_91 gnd C_wl
Rw58_91 word58_91 word57_91 R_wl
Cwl_58_91 word58_91 gnd C_wl
Rw59_91 word59_91 word58_91 R_wl
Cwl_59_91 word59_91 gnd C_wl
Rw60_91 word60_91 word59_91 R_wl
Cwl_60_91 word60_91 gnd C_wl
Rw61_91 word61_91 word60_91 R_wl
Cwl_61_91 word61_91 gnd C_wl
Rw62_91 word62_91 word61_91 R_wl
Cwl_62_91 word62_91 gnd C_wl
Rw63_91 word63_91 word62_91 R_wl
Cwl_63_91 word63_91 gnd C_wl
Rw64_91 word64_91 word63_91 R_wl
Cwl_64_91 word64_91 gnd C_wl
Rw65_91 word65_91 word64_91 R_wl
Cwl_65_91 word65_91 gnd C_wl
Rw66_91 word66_91 word65_91 R_wl
Cwl_66_91 word66_91 gnd C_wl
Rw67_91 word67_91 word66_91 R_wl
Cwl_67_91 word67_91 gnd C_wl
Rw68_91 word68_91 word67_91 R_wl
Cwl_68_91 word68_91 gnd C_wl
Rw69_91 word69_91 word68_91 R_wl
Cwl_69_91 word69_91 gnd C_wl
Rw70_91 word70_91 word69_91 R_wl
Cwl_70_91 word70_91 gnd C_wl
Rw71_91 word71_91 word70_91 R_wl
Cwl_71_91 word71_91 gnd C_wl
Rw72_91 word72_91 word71_91 R_wl
Cwl_72_91 word72_91 gnd C_wl
Rw73_91 word73_91 word72_91 R_wl
Cwl_73_91 word73_91 gnd C_wl
Rw74_91 word74_91 word73_91 R_wl
Cwl_74_91 word74_91 gnd C_wl
Rw75_91 word75_91 word74_91 R_wl
Cwl_75_91 word75_91 gnd C_wl
Rw76_91 word76_91 word75_91 R_wl
Cwl_76_91 word76_91 gnd C_wl
Rw77_91 word77_91 word76_91 R_wl
Cwl_77_91 word77_91 gnd C_wl
Rw78_91 word78_91 word77_91 R_wl
Cwl_78_91 word78_91 gnd C_wl
Rw79_91 word79_91 word78_91 R_wl
Cwl_79_91 word79_91 gnd C_wl
Rw80_91 word80_91 word79_91 R_wl
Cwl_80_91 word80_91 gnd C_wl
Rw81_91 word81_91 word80_91 R_wl
Cwl_81_91 word81_91 gnd C_wl
Rw82_91 word82_91 word81_91 R_wl
Cwl_82_91 word82_91 gnd C_wl
Rw83_91 word83_91 word82_91 R_wl
Cwl_83_91 word83_91 gnd C_wl
Rw84_91 word84_91 word83_91 R_wl
Cwl_84_91 word84_91 gnd C_wl
Rw85_91 word85_91 word84_91 R_wl
Cwl_85_91 word85_91 gnd C_wl
Rw86_91 word86_91 word85_91 R_wl
Cwl_86_91 word86_91 gnd C_wl
Rw87_91 word87_91 word86_91 R_wl
Cwl_87_91 word87_91 gnd C_wl
Rw88_91 word88_91 word87_91 R_wl
Cwl_88_91 word88_91 gnd C_wl
Rw89_91 word89_91 word88_91 R_wl
Cwl_89_91 word89_91 gnd C_wl
Rw90_91 word90_91 word89_91 R_wl
Cwl_90_91 word90_91 gnd C_wl
Rw91_91 word91_91 word90_91 R_wl
Cwl_91_91 word91_91 gnd C_wl
Rw92_91 word92_91 word91_91 R_wl
Cwl_92_91 word92_91 gnd C_wl
Rw93_91 word93_91 word92_91 R_wl
Cwl_93_91 word93_91 gnd C_wl
Rw94_91 word94_91 word93_91 R_wl
Cwl_94_91 word94_91 gnd C_wl
Rw95_91 word95_91 word94_91 R_wl
Cwl_95_91 word95_91 gnd C_wl
Rw96_91 word96_91 word95_91 R_wl
Cwl_96_91 word96_91 gnd C_wl
Rw97_91 word97_91 word96_91 R_wl
Cwl_97_91 word97_91 gnd C_wl
Rw98_91 word98_91 word97_91 R_wl
Cwl_98_91 word98_91 gnd C_wl
Rw99_91 word99_91 word98_91 R_wl
Cwl_99_91 word99_91 gnd C_wl
Vwl_92 word_92 0 0
Rw0_92 word_92 word0_92 R_wl
Cwl_0_92 word0_92 gnd C_wl
Rw1_92 word1_92 word0_92 R_wl
Cwl_1_92 word1_92 gnd C_wl
Rw2_92 word2_92 word1_92 R_wl
Cwl_2_92 word2_92 gnd C_wl
Rw3_92 word3_92 word2_92 R_wl
Cwl_3_92 word3_92 gnd C_wl
Rw4_92 word4_92 word3_92 R_wl
Cwl_4_92 word4_92 gnd C_wl
Rw5_92 word5_92 word4_92 R_wl
Cwl_5_92 word5_92 gnd C_wl
Rw6_92 word6_92 word5_92 R_wl
Cwl_6_92 word6_92 gnd C_wl
Rw7_92 word7_92 word6_92 R_wl
Cwl_7_92 word7_92 gnd C_wl
Rw8_92 word8_92 word7_92 R_wl
Cwl_8_92 word8_92 gnd C_wl
Rw9_92 word9_92 word8_92 R_wl
Cwl_9_92 word9_92 gnd C_wl
Rw10_92 word10_92 word9_92 R_wl
Cwl_10_92 word10_92 gnd C_wl
Rw11_92 word11_92 word10_92 R_wl
Cwl_11_92 word11_92 gnd C_wl
Rw12_92 word12_92 word11_92 R_wl
Cwl_12_92 word12_92 gnd C_wl
Rw13_92 word13_92 word12_92 R_wl
Cwl_13_92 word13_92 gnd C_wl
Rw14_92 word14_92 word13_92 R_wl
Cwl_14_92 word14_92 gnd C_wl
Rw15_92 word15_92 word14_92 R_wl
Cwl_15_92 word15_92 gnd C_wl
Rw16_92 word16_92 word15_92 R_wl
Cwl_16_92 word16_92 gnd C_wl
Rw17_92 word17_92 word16_92 R_wl
Cwl_17_92 word17_92 gnd C_wl
Rw18_92 word18_92 word17_92 R_wl
Cwl_18_92 word18_92 gnd C_wl
Rw19_92 word19_92 word18_92 R_wl
Cwl_19_92 word19_92 gnd C_wl
Rw20_92 word20_92 word19_92 R_wl
Cwl_20_92 word20_92 gnd C_wl
Rw21_92 word21_92 word20_92 R_wl
Cwl_21_92 word21_92 gnd C_wl
Rw22_92 word22_92 word21_92 R_wl
Cwl_22_92 word22_92 gnd C_wl
Rw23_92 word23_92 word22_92 R_wl
Cwl_23_92 word23_92 gnd C_wl
Rw24_92 word24_92 word23_92 R_wl
Cwl_24_92 word24_92 gnd C_wl
Rw25_92 word25_92 word24_92 R_wl
Cwl_25_92 word25_92 gnd C_wl
Rw26_92 word26_92 word25_92 R_wl
Cwl_26_92 word26_92 gnd C_wl
Rw27_92 word27_92 word26_92 R_wl
Cwl_27_92 word27_92 gnd C_wl
Rw28_92 word28_92 word27_92 R_wl
Cwl_28_92 word28_92 gnd C_wl
Rw29_92 word29_92 word28_92 R_wl
Cwl_29_92 word29_92 gnd C_wl
Rw30_92 word30_92 word29_92 R_wl
Cwl_30_92 word30_92 gnd C_wl
Rw31_92 word31_92 word30_92 R_wl
Cwl_31_92 word31_92 gnd C_wl
Rw32_92 word32_92 word31_92 R_wl
Cwl_32_92 word32_92 gnd C_wl
Rw33_92 word33_92 word32_92 R_wl
Cwl_33_92 word33_92 gnd C_wl
Rw34_92 word34_92 word33_92 R_wl
Cwl_34_92 word34_92 gnd C_wl
Rw35_92 word35_92 word34_92 R_wl
Cwl_35_92 word35_92 gnd C_wl
Rw36_92 word36_92 word35_92 R_wl
Cwl_36_92 word36_92 gnd C_wl
Rw37_92 word37_92 word36_92 R_wl
Cwl_37_92 word37_92 gnd C_wl
Rw38_92 word38_92 word37_92 R_wl
Cwl_38_92 word38_92 gnd C_wl
Rw39_92 word39_92 word38_92 R_wl
Cwl_39_92 word39_92 gnd C_wl
Rw40_92 word40_92 word39_92 R_wl
Cwl_40_92 word40_92 gnd C_wl
Rw41_92 word41_92 word40_92 R_wl
Cwl_41_92 word41_92 gnd C_wl
Rw42_92 word42_92 word41_92 R_wl
Cwl_42_92 word42_92 gnd C_wl
Rw43_92 word43_92 word42_92 R_wl
Cwl_43_92 word43_92 gnd C_wl
Rw44_92 word44_92 word43_92 R_wl
Cwl_44_92 word44_92 gnd C_wl
Rw45_92 word45_92 word44_92 R_wl
Cwl_45_92 word45_92 gnd C_wl
Rw46_92 word46_92 word45_92 R_wl
Cwl_46_92 word46_92 gnd C_wl
Rw47_92 word47_92 word46_92 R_wl
Cwl_47_92 word47_92 gnd C_wl
Rw48_92 word48_92 word47_92 R_wl
Cwl_48_92 word48_92 gnd C_wl
Rw49_92 word49_92 word48_92 R_wl
Cwl_49_92 word49_92 gnd C_wl
Rw50_92 word50_92 word49_92 R_wl
Cwl_50_92 word50_92 gnd C_wl
Rw51_92 word51_92 word50_92 R_wl
Cwl_51_92 word51_92 gnd C_wl
Rw52_92 word52_92 word51_92 R_wl
Cwl_52_92 word52_92 gnd C_wl
Rw53_92 word53_92 word52_92 R_wl
Cwl_53_92 word53_92 gnd C_wl
Rw54_92 word54_92 word53_92 R_wl
Cwl_54_92 word54_92 gnd C_wl
Rw55_92 word55_92 word54_92 R_wl
Cwl_55_92 word55_92 gnd C_wl
Rw56_92 word56_92 word55_92 R_wl
Cwl_56_92 word56_92 gnd C_wl
Rw57_92 word57_92 word56_92 R_wl
Cwl_57_92 word57_92 gnd C_wl
Rw58_92 word58_92 word57_92 R_wl
Cwl_58_92 word58_92 gnd C_wl
Rw59_92 word59_92 word58_92 R_wl
Cwl_59_92 word59_92 gnd C_wl
Rw60_92 word60_92 word59_92 R_wl
Cwl_60_92 word60_92 gnd C_wl
Rw61_92 word61_92 word60_92 R_wl
Cwl_61_92 word61_92 gnd C_wl
Rw62_92 word62_92 word61_92 R_wl
Cwl_62_92 word62_92 gnd C_wl
Rw63_92 word63_92 word62_92 R_wl
Cwl_63_92 word63_92 gnd C_wl
Rw64_92 word64_92 word63_92 R_wl
Cwl_64_92 word64_92 gnd C_wl
Rw65_92 word65_92 word64_92 R_wl
Cwl_65_92 word65_92 gnd C_wl
Rw66_92 word66_92 word65_92 R_wl
Cwl_66_92 word66_92 gnd C_wl
Rw67_92 word67_92 word66_92 R_wl
Cwl_67_92 word67_92 gnd C_wl
Rw68_92 word68_92 word67_92 R_wl
Cwl_68_92 word68_92 gnd C_wl
Rw69_92 word69_92 word68_92 R_wl
Cwl_69_92 word69_92 gnd C_wl
Rw70_92 word70_92 word69_92 R_wl
Cwl_70_92 word70_92 gnd C_wl
Rw71_92 word71_92 word70_92 R_wl
Cwl_71_92 word71_92 gnd C_wl
Rw72_92 word72_92 word71_92 R_wl
Cwl_72_92 word72_92 gnd C_wl
Rw73_92 word73_92 word72_92 R_wl
Cwl_73_92 word73_92 gnd C_wl
Rw74_92 word74_92 word73_92 R_wl
Cwl_74_92 word74_92 gnd C_wl
Rw75_92 word75_92 word74_92 R_wl
Cwl_75_92 word75_92 gnd C_wl
Rw76_92 word76_92 word75_92 R_wl
Cwl_76_92 word76_92 gnd C_wl
Rw77_92 word77_92 word76_92 R_wl
Cwl_77_92 word77_92 gnd C_wl
Rw78_92 word78_92 word77_92 R_wl
Cwl_78_92 word78_92 gnd C_wl
Rw79_92 word79_92 word78_92 R_wl
Cwl_79_92 word79_92 gnd C_wl
Rw80_92 word80_92 word79_92 R_wl
Cwl_80_92 word80_92 gnd C_wl
Rw81_92 word81_92 word80_92 R_wl
Cwl_81_92 word81_92 gnd C_wl
Rw82_92 word82_92 word81_92 R_wl
Cwl_82_92 word82_92 gnd C_wl
Rw83_92 word83_92 word82_92 R_wl
Cwl_83_92 word83_92 gnd C_wl
Rw84_92 word84_92 word83_92 R_wl
Cwl_84_92 word84_92 gnd C_wl
Rw85_92 word85_92 word84_92 R_wl
Cwl_85_92 word85_92 gnd C_wl
Rw86_92 word86_92 word85_92 R_wl
Cwl_86_92 word86_92 gnd C_wl
Rw87_92 word87_92 word86_92 R_wl
Cwl_87_92 word87_92 gnd C_wl
Rw88_92 word88_92 word87_92 R_wl
Cwl_88_92 word88_92 gnd C_wl
Rw89_92 word89_92 word88_92 R_wl
Cwl_89_92 word89_92 gnd C_wl
Rw90_92 word90_92 word89_92 R_wl
Cwl_90_92 word90_92 gnd C_wl
Rw91_92 word91_92 word90_92 R_wl
Cwl_91_92 word91_92 gnd C_wl
Rw92_92 word92_92 word91_92 R_wl
Cwl_92_92 word92_92 gnd C_wl
Rw93_92 word93_92 word92_92 R_wl
Cwl_93_92 word93_92 gnd C_wl
Rw94_92 word94_92 word93_92 R_wl
Cwl_94_92 word94_92 gnd C_wl
Rw95_92 word95_92 word94_92 R_wl
Cwl_95_92 word95_92 gnd C_wl
Rw96_92 word96_92 word95_92 R_wl
Cwl_96_92 word96_92 gnd C_wl
Rw97_92 word97_92 word96_92 R_wl
Cwl_97_92 word97_92 gnd C_wl
Rw98_92 word98_92 word97_92 R_wl
Cwl_98_92 word98_92 gnd C_wl
Rw99_92 word99_92 word98_92 R_wl
Cwl_99_92 word99_92 gnd C_wl
Vwl_93 word_93 0 0
Rw0_93 word_93 word0_93 R_wl
Cwl_0_93 word0_93 gnd C_wl
Rw1_93 word1_93 word0_93 R_wl
Cwl_1_93 word1_93 gnd C_wl
Rw2_93 word2_93 word1_93 R_wl
Cwl_2_93 word2_93 gnd C_wl
Rw3_93 word3_93 word2_93 R_wl
Cwl_3_93 word3_93 gnd C_wl
Rw4_93 word4_93 word3_93 R_wl
Cwl_4_93 word4_93 gnd C_wl
Rw5_93 word5_93 word4_93 R_wl
Cwl_5_93 word5_93 gnd C_wl
Rw6_93 word6_93 word5_93 R_wl
Cwl_6_93 word6_93 gnd C_wl
Rw7_93 word7_93 word6_93 R_wl
Cwl_7_93 word7_93 gnd C_wl
Rw8_93 word8_93 word7_93 R_wl
Cwl_8_93 word8_93 gnd C_wl
Rw9_93 word9_93 word8_93 R_wl
Cwl_9_93 word9_93 gnd C_wl
Rw10_93 word10_93 word9_93 R_wl
Cwl_10_93 word10_93 gnd C_wl
Rw11_93 word11_93 word10_93 R_wl
Cwl_11_93 word11_93 gnd C_wl
Rw12_93 word12_93 word11_93 R_wl
Cwl_12_93 word12_93 gnd C_wl
Rw13_93 word13_93 word12_93 R_wl
Cwl_13_93 word13_93 gnd C_wl
Rw14_93 word14_93 word13_93 R_wl
Cwl_14_93 word14_93 gnd C_wl
Rw15_93 word15_93 word14_93 R_wl
Cwl_15_93 word15_93 gnd C_wl
Rw16_93 word16_93 word15_93 R_wl
Cwl_16_93 word16_93 gnd C_wl
Rw17_93 word17_93 word16_93 R_wl
Cwl_17_93 word17_93 gnd C_wl
Rw18_93 word18_93 word17_93 R_wl
Cwl_18_93 word18_93 gnd C_wl
Rw19_93 word19_93 word18_93 R_wl
Cwl_19_93 word19_93 gnd C_wl
Rw20_93 word20_93 word19_93 R_wl
Cwl_20_93 word20_93 gnd C_wl
Rw21_93 word21_93 word20_93 R_wl
Cwl_21_93 word21_93 gnd C_wl
Rw22_93 word22_93 word21_93 R_wl
Cwl_22_93 word22_93 gnd C_wl
Rw23_93 word23_93 word22_93 R_wl
Cwl_23_93 word23_93 gnd C_wl
Rw24_93 word24_93 word23_93 R_wl
Cwl_24_93 word24_93 gnd C_wl
Rw25_93 word25_93 word24_93 R_wl
Cwl_25_93 word25_93 gnd C_wl
Rw26_93 word26_93 word25_93 R_wl
Cwl_26_93 word26_93 gnd C_wl
Rw27_93 word27_93 word26_93 R_wl
Cwl_27_93 word27_93 gnd C_wl
Rw28_93 word28_93 word27_93 R_wl
Cwl_28_93 word28_93 gnd C_wl
Rw29_93 word29_93 word28_93 R_wl
Cwl_29_93 word29_93 gnd C_wl
Rw30_93 word30_93 word29_93 R_wl
Cwl_30_93 word30_93 gnd C_wl
Rw31_93 word31_93 word30_93 R_wl
Cwl_31_93 word31_93 gnd C_wl
Rw32_93 word32_93 word31_93 R_wl
Cwl_32_93 word32_93 gnd C_wl
Rw33_93 word33_93 word32_93 R_wl
Cwl_33_93 word33_93 gnd C_wl
Rw34_93 word34_93 word33_93 R_wl
Cwl_34_93 word34_93 gnd C_wl
Rw35_93 word35_93 word34_93 R_wl
Cwl_35_93 word35_93 gnd C_wl
Rw36_93 word36_93 word35_93 R_wl
Cwl_36_93 word36_93 gnd C_wl
Rw37_93 word37_93 word36_93 R_wl
Cwl_37_93 word37_93 gnd C_wl
Rw38_93 word38_93 word37_93 R_wl
Cwl_38_93 word38_93 gnd C_wl
Rw39_93 word39_93 word38_93 R_wl
Cwl_39_93 word39_93 gnd C_wl
Rw40_93 word40_93 word39_93 R_wl
Cwl_40_93 word40_93 gnd C_wl
Rw41_93 word41_93 word40_93 R_wl
Cwl_41_93 word41_93 gnd C_wl
Rw42_93 word42_93 word41_93 R_wl
Cwl_42_93 word42_93 gnd C_wl
Rw43_93 word43_93 word42_93 R_wl
Cwl_43_93 word43_93 gnd C_wl
Rw44_93 word44_93 word43_93 R_wl
Cwl_44_93 word44_93 gnd C_wl
Rw45_93 word45_93 word44_93 R_wl
Cwl_45_93 word45_93 gnd C_wl
Rw46_93 word46_93 word45_93 R_wl
Cwl_46_93 word46_93 gnd C_wl
Rw47_93 word47_93 word46_93 R_wl
Cwl_47_93 word47_93 gnd C_wl
Rw48_93 word48_93 word47_93 R_wl
Cwl_48_93 word48_93 gnd C_wl
Rw49_93 word49_93 word48_93 R_wl
Cwl_49_93 word49_93 gnd C_wl
Rw50_93 word50_93 word49_93 R_wl
Cwl_50_93 word50_93 gnd C_wl
Rw51_93 word51_93 word50_93 R_wl
Cwl_51_93 word51_93 gnd C_wl
Rw52_93 word52_93 word51_93 R_wl
Cwl_52_93 word52_93 gnd C_wl
Rw53_93 word53_93 word52_93 R_wl
Cwl_53_93 word53_93 gnd C_wl
Rw54_93 word54_93 word53_93 R_wl
Cwl_54_93 word54_93 gnd C_wl
Rw55_93 word55_93 word54_93 R_wl
Cwl_55_93 word55_93 gnd C_wl
Rw56_93 word56_93 word55_93 R_wl
Cwl_56_93 word56_93 gnd C_wl
Rw57_93 word57_93 word56_93 R_wl
Cwl_57_93 word57_93 gnd C_wl
Rw58_93 word58_93 word57_93 R_wl
Cwl_58_93 word58_93 gnd C_wl
Rw59_93 word59_93 word58_93 R_wl
Cwl_59_93 word59_93 gnd C_wl
Rw60_93 word60_93 word59_93 R_wl
Cwl_60_93 word60_93 gnd C_wl
Rw61_93 word61_93 word60_93 R_wl
Cwl_61_93 word61_93 gnd C_wl
Rw62_93 word62_93 word61_93 R_wl
Cwl_62_93 word62_93 gnd C_wl
Rw63_93 word63_93 word62_93 R_wl
Cwl_63_93 word63_93 gnd C_wl
Rw64_93 word64_93 word63_93 R_wl
Cwl_64_93 word64_93 gnd C_wl
Rw65_93 word65_93 word64_93 R_wl
Cwl_65_93 word65_93 gnd C_wl
Rw66_93 word66_93 word65_93 R_wl
Cwl_66_93 word66_93 gnd C_wl
Rw67_93 word67_93 word66_93 R_wl
Cwl_67_93 word67_93 gnd C_wl
Rw68_93 word68_93 word67_93 R_wl
Cwl_68_93 word68_93 gnd C_wl
Rw69_93 word69_93 word68_93 R_wl
Cwl_69_93 word69_93 gnd C_wl
Rw70_93 word70_93 word69_93 R_wl
Cwl_70_93 word70_93 gnd C_wl
Rw71_93 word71_93 word70_93 R_wl
Cwl_71_93 word71_93 gnd C_wl
Rw72_93 word72_93 word71_93 R_wl
Cwl_72_93 word72_93 gnd C_wl
Rw73_93 word73_93 word72_93 R_wl
Cwl_73_93 word73_93 gnd C_wl
Rw74_93 word74_93 word73_93 R_wl
Cwl_74_93 word74_93 gnd C_wl
Rw75_93 word75_93 word74_93 R_wl
Cwl_75_93 word75_93 gnd C_wl
Rw76_93 word76_93 word75_93 R_wl
Cwl_76_93 word76_93 gnd C_wl
Rw77_93 word77_93 word76_93 R_wl
Cwl_77_93 word77_93 gnd C_wl
Rw78_93 word78_93 word77_93 R_wl
Cwl_78_93 word78_93 gnd C_wl
Rw79_93 word79_93 word78_93 R_wl
Cwl_79_93 word79_93 gnd C_wl
Rw80_93 word80_93 word79_93 R_wl
Cwl_80_93 word80_93 gnd C_wl
Rw81_93 word81_93 word80_93 R_wl
Cwl_81_93 word81_93 gnd C_wl
Rw82_93 word82_93 word81_93 R_wl
Cwl_82_93 word82_93 gnd C_wl
Rw83_93 word83_93 word82_93 R_wl
Cwl_83_93 word83_93 gnd C_wl
Rw84_93 word84_93 word83_93 R_wl
Cwl_84_93 word84_93 gnd C_wl
Rw85_93 word85_93 word84_93 R_wl
Cwl_85_93 word85_93 gnd C_wl
Rw86_93 word86_93 word85_93 R_wl
Cwl_86_93 word86_93 gnd C_wl
Rw87_93 word87_93 word86_93 R_wl
Cwl_87_93 word87_93 gnd C_wl
Rw88_93 word88_93 word87_93 R_wl
Cwl_88_93 word88_93 gnd C_wl
Rw89_93 word89_93 word88_93 R_wl
Cwl_89_93 word89_93 gnd C_wl
Rw90_93 word90_93 word89_93 R_wl
Cwl_90_93 word90_93 gnd C_wl
Rw91_93 word91_93 word90_93 R_wl
Cwl_91_93 word91_93 gnd C_wl
Rw92_93 word92_93 word91_93 R_wl
Cwl_92_93 word92_93 gnd C_wl
Rw93_93 word93_93 word92_93 R_wl
Cwl_93_93 word93_93 gnd C_wl
Rw94_93 word94_93 word93_93 R_wl
Cwl_94_93 word94_93 gnd C_wl
Rw95_93 word95_93 word94_93 R_wl
Cwl_95_93 word95_93 gnd C_wl
Rw96_93 word96_93 word95_93 R_wl
Cwl_96_93 word96_93 gnd C_wl
Rw97_93 word97_93 word96_93 R_wl
Cwl_97_93 word97_93 gnd C_wl
Rw98_93 word98_93 word97_93 R_wl
Cwl_98_93 word98_93 gnd C_wl
Rw99_93 word99_93 word98_93 R_wl
Cwl_99_93 word99_93 gnd C_wl
Vwl_94 word_94 0 0
Rw0_94 word_94 word0_94 R_wl
Cwl_0_94 word0_94 gnd C_wl
Rw1_94 word1_94 word0_94 R_wl
Cwl_1_94 word1_94 gnd C_wl
Rw2_94 word2_94 word1_94 R_wl
Cwl_2_94 word2_94 gnd C_wl
Rw3_94 word3_94 word2_94 R_wl
Cwl_3_94 word3_94 gnd C_wl
Rw4_94 word4_94 word3_94 R_wl
Cwl_4_94 word4_94 gnd C_wl
Rw5_94 word5_94 word4_94 R_wl
Cwl_5_94 word5_94 gnd C_wl
Rw6_94 word6_94 word5_94 R_wl
Cwl_6_94 word6_94 gnd C_wl
Rw7_94 word7_94 word6_94 R_wl
Cwl_7_94 word7_94 gnd C_wl
Rw8_94 word8_94 word7_94 R_wl
Cwl_8_94 word8_94 gnd C_wl
Rw9_94 word9_94 word8_94 R_wl
Cwl_9_94 word9_94 gnd C_wl
Rw10_94 word10_94 word9_94 R_wl
Cwl_10_94 word10_94 gnd C_wl
Rw11_94 word11_94 word10_94 R_wl
Cwl_11_94 word11_94 gnd C_wl
Rw12_94 word12_94 word11_94 R_wl
Cwl_12_94 word12_94 gnd C_wl
Rw13_94 word13_94 word12_94 R_wl
Cwl_13_94 word13_94 gnd C_wl
Rw14_94 word14_94 word13_94 R_wl
Cwl_14_94 word14_94 gnd C_wl
Rw15_94 word15_94 word14_94 R_wl
Cwl_15_94 word15_94 gnd C_wl
Rw16_94 word16_94 word15_94 R_wl
Cwl_16_94 word16_94 gnd C_wl
Rw17_94 word17_94 word16_94 R_wl
Cwl_17_94 word17_94 gnd C_wl
Rw18_94 word18_94 word17_94 R_wl
Cwl_18_94 word18_94 gnd C_wl
Rw19_94 word19_94 word18_94 R_wl
Cwl_19_94 word19_94 gnd C_wl
Rw20_94 word20_94 word19_94 R_wl
Cwl_20_94 word20_94 gnd C_wl
Rw21_94 word21_94 word20_94 R_wl
Cwl_21_94 word21_94 gnd C_wl
Rw22_94 word22_94 word21_94 R_wl
Cwl_22_94 word22_94 gnd C_wl
Rw23_94 word23_94 word22_94 R_wl
Cwl_23_94 word23_94 gnd C_wl
Rw24_94 word24_94 word23_94 R_wl
Cwl_24_94 word24_94 gnd C_wl
Rw25_94 word25_94 word24_94 R_wl
Cwl_25_94 word25_94 gnd C_wl
Rw26_94 word26_94 word25_94 R_wl
Cwl_26_94 word26_94 gnd C_wl
Rw27_94 word27_94 word26_94 R_wl
Cwl_27_94 word27_94 gnd C_wl
Rw28_94 word28_94 word27_94 R_wl
Cwl_28_94 word28_94 gnd C_wl
Rw29_94 word29_94 word28_94 R_wl
Cwl_29_94 word29_94 gnd C_wl
Rw30_94 word30_94 word29_94 R_wl
Cwl_30_94 word30_94 gnd C_wl
Rw31_94 word31_94 word30_94 R_wl
Cwl_31_94 word31_94 gnd C_wl
Rw32_94 word32_94 word31_94 R_wl
Cwl_32_94 word32_94 gnd C_wl
Rw33_94 word33_94 word32_94 R_wl
Cwl_33_94 word33_94 gnd C_wl
Rw34_94 word34_94 word33_94 R_wl
Cwl_34_94 word34_94 gnd C_wl
Rw35_94 word35_94 word34_94 R_wl
Cwl_35_94 word35_94 gnd C_wl
Rw36_94 word36_94 word35_94 R_wl
Cwl_36_94 word36_94 gnd C_wl
Rw37_94 word37_94 word36_94 R_wl
Cwl_37_94 word37_94 gnd C_wl
Rw38_94 word38_94 word37_94 R_wl
Cwl_38_94 word38_94 gnd C_wl
Rw39_94 word39_94 word38_94 R_wl
Cwl_39_94 word39_94 gnd C_wl
Rw40_94 word40_94 word39_94 R_wl
Cwl_40_94 word40_94 gnd C_wl
Rw41_94 word41_94 word40_94 R_wl
Cwl_41_94 word41_94 gnd C_wl
Rw42_94 word42_94 word41_94 R_wl
Cwl_42_94 word42_94 gnd C_wl
Rw43_94 word43_94 word42_94 R_wl
Cwl_43_94 word43_94 gnd C_wl
Rw44_94 word44_94 word43_94 R_wl
Cwl_44_94 word44_94 gnd C_wl
Rw45_94 word45_94 word44_94 R_wl
Cwl_45_94 word45_94 gnd C_wl
Rw46_94 word46_94 word45_94 R_wl
Cwl_46_94 word46_94 gnd C_wl
Rw47_94 word47_94 word46_94 R_wl
Cwl_47_94 word47_94 gnd C_wl
Rw48_94 word48_94 word47_94 R_wl
Cwl_48_94 word48_94 gnd C_wl
Rw49_94 word49_94 word48_94 R_wl
Cwl_49_94 word49_94 gnd C_wl
Rw50_94 word50_94 word49_94 R_wl
Cwl_50_94 word50_94 gnd C_wl
Rw51_94 word51_94 word50_94 R_wl
Cwl_51_94 word51_94 gnd C_wl
Rw52_94 word52_94 word51_94 R_wl
Cwl_52_94 word52_94 gnd C_wl
Rw53_94 word53_94 word52_94 R_wl
Cwl_53_94 word53_94 gnd C_wl
Rw54_94 word54_94 word53_94 R_wl
Cwl_54_94 word54_94 gnd C_wl
Rw55_94 word55_94 word54_94 R_wl
Cwl_55_94 word55_94 gnd C_wl
Rw56_94 word56_94 word55_94 R_wl
Cwl_56_94 word56_94 gnd C_wl
Rw57_94 word57_94 word56_94 R_wl
Cwl_57_94 word57_94 gnd C_wl
Rw58_94 word58_94 word57_94 R_wl
Cwl_58_94 word58_94 gnd C_wl
Rw59_94 word59_94 word58_94 R_wl
Cwl_59_94 word59_94 gnd C_wl
Rw60_94 word60_94 word59_94 R_wl
Cwl_60_94 word60_94 gnd C_wl
Rw61_94 word61_94 word60_94 R_wl
Cwl_61_94 word61_94 gnd C_wl
Rw62_94 word62_94 word61_94 R_wl
Cwl_62_94 word62_94 gnd C_wl
Rw63_94 word63_94 word62_94 R_wl
Cwl_63_94 word63_94 gnd C_wl
Rw64_94 word64_94 word63_94 R_wl
Cwl_64_94 word64_94 gnd C_wl
Rw65_94 word65_94 word64_94 R_wl
Cwl_65_94 word65_94 gnd C_wl
Rw66_94 word66_94 word65_94 R_wl
Cwl_66_94 word66_94 gnd C_wl
Rw67_94 word67_94 word66_94 R_wl
Cwl_67_94 word67_94 gnd C_wl
Rw68_94 word68_94 word67_94 R_wl
Cwl_68_94 word68_94 gnd C_wl
Rw69_94 word69_94 word68_94 R_wl
Cwl_69_94 word69_94 gnd C_wl
Rw70_94 word70_94 word69_94 R_wl
Cwl_70_94 word70_94 gnd C_wl
Rw71_94 word71_94 word70_94 R_wl
Cwl_71_94 word71_94 gnd C_wl
Rw72_94 word72_94 word71_94 R_wl
Cwl_72_94 word72_94 gnd C_wl
Rw73_94 word73_94 word72_94 R_wl
Cwl_73_94 word73_94 gnd C_wl
Rw74_94 word74_94 word73_94 R_wl
Cwl_74_94 word74_94 gnd C_wl
Rw75_94 word75_94 word74_94 R_wl
Cwl_75_94 word75_94 gnd C_wl
Rw76_94 word76_94 word75_94 R_wl
Cwl_76_94 word76_94 gnd C_wl
Rw77_94 word77_94 word76_94 R_wl
Cwl_77_94 word77_94 gnd C_wl
Rw78_94 word78_94 word77_94 R_wl
Cwl_78_94 word78_94 gnd C_wl
Rw79_94 word79_94 word78_94 R_wl
Cwl_79_94 word79_94 gnd C_wl
Rw80_94 word80_94 word79_94 R_wl
Cwl_80_94 word80_94 gnd C_wl
Rw81_94 word81_94 word80_94 R_wl
Cwl_81_94 word81_94 gnd C_wl
Rw82_94 word82_94 word81_94 R_wl
Cwl_82_94 word82_94 gnd C_wl
Rw83_94 word83_94 word82_94 R_wl
Cwl_83_94 word83_94 gnd C_wl
Rw84_94 word84_94 word83_94 R_wl
Cwl_84_94 word84_94 gnd C_wl
Rw85_94 word85_94 word84_94 R_wl
Cwl_85_94 word85_94 gnd C_wl
Rw86_94 word86_94 word85_94 R_wl
Cwl_86_94 word86_94 gnd C_wl
Rw87_94 word87_94 word86_94 R_wl
Cwl_87_94 word87_94 gnd C_wl
Rw88_94 word88_94 word87_94 R_wl
Cwl_88_94 word88_94 gnd C_wl
Rw89_94 word89_94 word88_94 R_wl
Cwl_89_94 word89_94 gnd C_wl
Rw90_94 word90_94 word89_94 R_wl
Cwl_90_94 word90_94 gnd C_wl
Rw91_94 word91_94 word90_94 R_wl
Cwl_91_94 word91_94 gnd C_wl
Rw92_94 word92_94 word91_94 R_wl
Cwl_92_94 word92_94 gnd C_wl
Rw93_94 word93_94 word92_94 R_wl
Cwl_93_94 word93_94 gnd C_wl
Rw94_94 word94_94 word93_94 R_wl
Cwl_94_94 word94_94 gnd C_wl
Rw95_94 word95_94 word94_94 R_wl
Cwl_95_94 word95_94 gnd C_wl
Rw96_94 word96_94 word95_94 R_wl
Cwl_96_94 word96_94 gnd C_wl
Rw97_94 word97_94 word96_94 R_wl
Cwl_97_94 word97_94 gnd C_wl
Rw98_94 word98_94 word97_94 R_wl
Cwl_98_94 word98_94 gnd C_wl
Rw99_94 word99_94 word98_94 R_wl
Cwl_99_94 word99_94 gnd C_wl
Vwl_95 word_95 0 0
Rw0_95 word_95 word0_95 R_wl
Cwl_0_95 word0_95 gnd C_wl
Rw1_95 word1_95 word0_95 R_wl
Cwl_1_95 word1_95 gnd C_wl
Rw2_95 word2_95 word1_95 R_wl
Cwl_2_95 word2_95 gnd C_wl
Rw3_95 word3_95 word2_95 R_wl
Cwl_3_95 word3_95 gnd C_wl
Rw4_95 word4_95 word3_95 R_wl
Cwl_4_95 word4_95 gnd C_wl
Rw5_95 word5_95 word4_95 R_wl
Cwl_5_95 word5_95 gnd C_wl
Rw6_95 word6_95 word5_95 R_wl
Cwl_6_95 word6_95 gnd C_wl
Rw7_95 word7_95 word6_95 R_wl
Cwl_7_95 word7_95 gnd C_wl
Rw8_95 word8_95 word7_95 R_wl
Cwl_8_95 word8_95 gnd C_wl
Rw9_95 word9_95 word8_95 R_wl
Cwl_9_95 word9_95 gnd C_wl
Rw10_95 word10_95 word9_95 R_wl
Cwl_10_95 word10_95 gnd C_wl
Rw11_95 word11_95 word10_95 R_wl
Cwl_11_95 word11_95 gnd C_wl
Rw12_95 word12_95 word11_95 R_wl
Cwl_12_95 word12_95 gnd C_wl
Rw13_95 word13_95 word12_95 R_wl
Cwl_13_95 word13_95 gnd C_wl
Rw14_95 word14_95 word13_95 R_wl
Cwl_14_95 word14_95 gnd C_wl
Rw15_95 word15_95 word14_95 R_wl
Cwl_15_95 word15_95 gnd C_wl
Rw16_95 word16_95 word15_95 R_wl
Cwl_16_95 word16_95 gnd C_wl
Rw17_95 word17_95 word16_95 R_wl
Cwl_17_95 word17_95 gnd C_wl
Rw18_95 word18_95 word17_95 R_wl
Cwl_18_95 word18_95 gnd C_wl
Rw19_95 word19_95 word18_95 R_wl
Cwl_19_95 word19_95 gnd C_wl
Rw20_95 word20_95 word19_95 R_wl
Cwl_20_95 word20_95 gnd C_wl
Rw21_95 word21_95 word20_95 R_wl
Cwl_21_95 word21_95 gnd C_wl
Rw22_95 word22_95 word21_95 R_wl
Cwl_22_95 word22_95 gnd C_wl
Rw23_95 word23_95 word22_95 R_wl
Cwl_23_95 word23_95 gnd C_wl
Rw24_95 word24_95 word23_95 R_wl
Cwl_24_95 word24_95 gnd C_wl
Rw25_95 word25_95 word24_95 R_wl
Cwl_25_95 word25_95 gnd C_wl
Rw26_95 word26_95 word25_95 R_wl
Cwl_26_95 word26_95 gnd C_wl
Rw27_95 word27_95 word26_95 R_wl
Cwl_27_95 word27_95 gnd C_wl
Rw28_95 word28_95 word27_95 R_wl
Cwl_28_95 word28_95 gnd C_wl
Rw29_95 word29_95 word28_95 R_wl
Cwl_29_95 word29_95 gnd C_wl
Rw30_95 word30_95 word29_95 R_wl
Cwl_30_95 word30_95 gnd C_wl
Rw31_95 word31_95 word30_95 R_wl
Cwl_31_95 word31_95 gnd C_wl
Rw32_95 word32_95 word31_95 R_wl
Cwl_32_95 word32_95 gnd C_wl
Rw33_95 word33_95 word32_95 R_wl
Cwl_33_95 word33_95 gnd C_wl
Rw34_95 word34_95 word33_95 R_wl
Cwl_34_95 word34_95 gnd C_wl
Rw35_95 word35_95 word34_95 R_wl
Cwl_35_95 word35_95 gnd C_wl
Rw36_95 word36_95 word35_95 R_wl
Cwl_36_95 word36_95 gnd C_wl
Rw37_95 word37_95 word36_95 R_wl
Cwl_37_95 word37_95 gnd C_wl
Rw38_95 word38_95 word37_95 R_wl
Cwl_38_95 word38_95 gnd C_wl
Rw39_95 word39_95 word38_95 R_wl
Cwl_39_95 word39_95 gnd C_wl
Rw40_95 word40_95 word39_95 R_wl
Cwl_40_95 word40_95 gnd C_wl
Rw41_95 word41_95 word40_95 R_wl
Cwl_41_95 word41_95 gnd C_wl
Rw42_95 word42_95 word41_95 R_wl
Cwl_42_95 word42_95 gnd C_wl
Rw43_95 word43_95 word42_95 R_wl
Cwl_43_95 word43_95 gnd C_wl
Rw44_95 word44_95 word43_95 R_wl
Cwl_44_95 word44_95 gnd C_wl
Rw45_95 word45_95 word44_95 R_wl
Cwl_45_95 word45_95 gnd C_wl
Rw46_95 word46_95 word45_95 R_wl
Cwl_46_95 word46_95 gnd C_wl
Rw47_95 word47_95 word46_95 R_wl
Cwl_47_95 word47_95 gnd C_wl
Rw48_95 word48_95 word47_95 R_wl
Cwl_48_95 word48_95 gnd C_wl
Rw49_95 word49_95 word48_95 R_wl
Cwl_49_95 word49_95 gnd C_wl
Rw50_95 word50_95 word49_95 R_wl
Cwl_50_95 word50_95 gnd C_wl
Rw51_95 word51_95 word50_95 R_wl
Cwl_51_95 word51_95 gnd C_wl
Rw52_95 word52_95 word51_95 R_wl
Cwl_52_95 word52_95 gnd C_wl
Rw53_95 word53_95 word52_95 R_wl
Cwl_53_95 word53_95 gnd C_wl
Rw54_95 word54_95 word53_95 R_wl
Cwl_54_95 word54_95 gnd C_wl
Rw55_95 word55_95 word54_95 R_wl
Cwl_55_95 word55_95 gnd C_wl
Rw56_95 word56_95 word55_95 R_wl
Cwl_56_95 word56_95 gnd C_wl
Rw57_95 word57_95 word56_95 R_wl
Cwl_57_95 word57_95 gnd C_wl
Rw58_95 word58_95 word57_95 R_wl
Cwl_58_95 word58_95 gnd C_wl
Rw59_95 word59_95 word58_95 R_wl
Cwl_59_95 word59_95 gnd C_wl
Rw60_95 word60_95 word59_95 R_wl
Cwl_60_95 word60_95 gnd C_wl
Rw61_95 word61_95 word60_95 R_wl
Cwl_61_95 word61_95 gnd C_wl
Rw62_95 word62_95 word61_95 R_wl
Cwl_62_95 word62_95 gnd C_wl
Rw63_95 word63_95 word62_95 R_wl
Cwl_63_95 word63_95 gnd C_wl
Rw64_95 word64_95 word63_95 R_wl
Cwl_64_95 word64_95 gnd C_wl
Rw65_95 word65_95 word64_95 R_wl
Cwl_65_95 word65_95 gnd C_wl
Rw66_95 word66_95 word65_95 R_wl
Cwl_66_95 word66_95 gnd C_wl
Rw67_95 word67_95 word66_95 R_wl
Cwl_67_95 word67_95 gnd C_wl
Rw68_95 word68_95 word67_95 R_wl
Cwl_68_95 word68_95 gnd C_wl
Rw69_95 word69_95 word68_95 R_wl
Cwl_69_95 word69_95 gnd C_wl
Rw70_95 word70_95 word69_95 R_wl
Cwl_70_95 word70_95 gnd C_wl
Rw71_95 word71_95 word70_95 R_wl
Cwl_71_95 word71_95 gnd C_wl
Rw72_95 word72_95 word71_95 R_wl
Cwl_72_95 word72_95 gnd C_wl
Rw73_95 word73_95 word72_95 R_wl
Cwl_73_95 word73_95 gnd C_wl
Rw74_95 word74_95 word73_95 R_wl
Cwl_74_95 word74_95 gnd C_wl
Rw75_95 word75_95 word74_95 R_wl
Cwl_75_95 word75_95 gnd C_wl
Rw76_95 word76_95 word75_95 R_wl
Cwl_76_95 word76_95 gnd C_wl
Rw77_95 word77_95 word76_95 R_wl
Cwl_77_95 word77_95 gnd C_wl
Rw78_95 word78_95 word77_95 R_wl
Cwl_78_95 word78_95 gnd C_wl
Rw79_95 word79_95 word78_95 R_wl
Cwl_79_95 word79_95 gnd C_wl
Rw80_95 word80_95 word79_95 R_wl
Cwl_80_95 word80_95 gnd C_wl
Rw81_95 word81_95 word80_95 R_wl
Cwl_81_95 word81_95 gnd C_wl
Rw82_95 word82_95 word81_95 R_wl
Cwl_82_95 word82_95 gnd C_wl
Rw83_95 word83_95 word82_95 R_wl
Cwl_83_95 word83_95 gnd C_wl
Rw84_95 word84_95 word83_95 R_wl
Cwl_84_95 word84_95 gnd C_wl
Rw85_95 word85_95 word84_95 R_wl
Cwl_85_95 word85_95 gnd C_wl
Rw86_95 word86_95 word85_95 R_wl
Cwl_86_95 word86_95 gnd C_wl
Rw87_95 word87_95 word86_95 R_wl
Cwl_87_95 word87_95 gnd C_wl
Rw88_95 word88_95 word87_95 R_wl
Cwl_88_95 word88_95 gnd C_wl
Rw89_95 word89_95 word88_95 R_wl
Cwl_89_95 word89_95 gnd C_wl
Rw90_95 word90_95 word89_95 R_wl
Cwl_90_95 word90_95 gnd C_wl
Rw91_95 word91_95 word90_95 R_wl
Cwl_91_95 word91_95 gnd C_wl
Rw92_95 word92_95 word91_95 R_wl
Cwl_92_95 word92_95 gnd C_wl
Rw93_95 word93_95 word92_95 R_wl
Cwl_93_95 word93_95 gnd C_wl
Rw94_95 word94_95 word93_95 R_wl
Cwl_94_95 word94_95 gnd C_wl
Rw95_95 word95_95 word94_95 R_wl
Cwl_95_95 word95_95 gnd C_wl
Rw96_95 word96_95 word95_95 R_wl
Cwl_96_95 word96_95 gnd C_wl
Rw97_95 word97_95 word96_95 R_wl
Cwl_97_95 word97_95 gnd C_wl
Rw98_95 word98_95 word97_95 R_wl
Cwl_98_95 word98_95 gnd C_wl
Rw99_95 word99_95 word98_95 R_wl
Cwl_99_95 word99_95 gnd C_wl
Vwl_96 word_96 0 0
Rw0_96 word_96 word0_96 R_wl
Cwl_0_96 word0_96 gnd C_wl
Rw1_96 word1_96 word0_96 R_wl
Cwl_1_96 word1_96 gnd C_wl
Rw2_96 word2_96 word1_96 R_wl
Cwl_2_96 word2_96 gnd C_wl
Rw3_96 word3_96 word2_96 R_wl
Cwl_3_96 word3_96 gnd C_wl
Rw4_96 word4_96 word3_96 R_wl
Cwl_4_96 word4_96 gnd C_wl
Rw5_96 word5_96 word4_96 R_wl
Cwl_5_96 word5_96 gnd C_wl
Rw6_96 word6_96 word5_96 R_wl
Cwl_6_96 word6_96 gnd C_wl
Rw7_96 word7_96 word6_96 R_wl
Cwl_7_96 word7_96 gnd C_wl
Rw8_96 word8_96 word7_96 R_wl
Cwl_8_96 word8_96 gnd C_wl
Rw9_96 word9_96 word8_96 R_wl
Cwl_9_96 word9_96 gnd C_wl
Rw10_96 word10_96 word9_96 R_wl
Cwl_10_96 word10_96 gnd C_wl
Rw11_96 word11_96 word10_96 R_wl
Cwl_11_96 word11_96 gnd C_wl
Rw12_96 word12_96 word11_96 R_wl
Cwl_12_96 word12_96 gnd C_wl
Rw13_96 word13_96 word12_96 R_wl
Cwl_13_96 word13_96 gnd C_wl
Rw14_96 word14_96 word13_96 R_wl
Cwl_14_96 word14_96 gnd C_wl
Rw15_96 word15_96 word14_96 R_wl
Cwl_15_96 word15_96 gnd C_wl
Rw16_96 word16_96 word15_96 R_wl
Cwl_16_96 word16_96 gnd C_wl
Rw17_96 word17_96 word16_96 R_wl
Cwl_17_96 word17_96 gnd C_wl
Rw18_96 word18_96 word17_96 R_wl
Cwl_18_96 word18_96 gnd C_wl
Rw19_96 word19_96 word18_96 R_wl
Cwl_19_96 word19_96 gnd C_wl
Rw20_96 word20_96 word19_96 R_wl
Cwl_20_96 word20_96 gnd C_wl
Rw21_96 word21_96 word20_96 R_wl
Cwl_21_96 word21_96 gnd C_wl
Rw22_96 word22_96 word21_96 R_wl
Cwl_22_96 word22_96 gnd C_wl
Rw23_96 word23_96 word22_96 R_wl
Cwl_23_96 word23_96 gnd C_wl
Rw24_96 word24_96 word23_96 R_wl
Cwl_24_96 word24_96 gnd C_wl
Rw25_96 word25_96 word24_96 R_wl
Cwl_25_96 word25_96 gnd C_wl
Rw26_96 word26_96 word25_96 R_wl
Cwl_26_96 word26_96 gnd C_wl
Rw27_96 word27_96 word26_96 R_wl
Cwl_27_96 word27_96 gnd C_wl
Rw28_96 word28_96 word27_96 R_wl
Cwl_28_96 word28_96 gnd C_wl
Rw29_96 word29_96 word28_96 R_wl
Cwl_29_96 word29_96 gnd C_wl
Rw30_96 word30_96 word29_96 R_wl
Cwl_30_96 word30_96 gnd C_wl
Rw31_96 word31_96 word30_96 R_wl
Cwl_31_96 word31_96 gnd C_wl
Rw32_96 word32_96 word31_96 R_wl
Cwl_32_96 word32_96 gnd C_wl
Rw33_96 word33_96 word32_96 R_wl
Cwl_33_96 word33_96 gnd C_wl
Rw34_96 word34_96 word33_96 R_wl
Cwl_34_96 word34_96 gnd C_wl
Rw35_96 word35_96 word34_96 R_wl
Cwl_35_96 word35_96 gnd C_wl
Rw36_96 word36_96 word35_96 R_wl
Cwl_36_96 word36_96 gnd C_wl
Rw37_96 word37_96 word36_96 R_wl
Cwl_37_96 word37_96 gnd C_wl
Rw38_96 word38_96 word37_96 R_wl
Cwl_38_96 word38_96 gnd C_wl
Rw39_96 word39_96 word38_96 R_wl
Cwl_39_96 word39_96 gnd C_wl
Rw40_96 word40_96 word39_96 R_wl
Cwl_40_96 word40_96 gnd C_wl
Rw41_96 word41_96 word40_96 R_wl
Cwl_41_96 word41_96 gnd C_wl
Rw42_96 word42_96 word41_96 R_wl
Cwl_42_96 word42_96 gnd C_wl
Rw43_96 word43_96 word42_96 R_wl
Cwl_43_96 word43_96 gnd C_wl
Rw44_96 word44_96 word43_96 R_wl
Cwl_44_96 word44_96 gnd C_wl
Rw45_96 word45_96 word44_96 R_wl
Cwl_45_96 word45_96 gnd C_wl
Rw46_96 word46_96 word45_96 R_wl
Cwl_46_96 word46_96 gnd C_wl
Rw47_96 word47_96 word46_96 R_wl
Cwl_47_96 word47_96 gnd C_wl
Rw48_96 word48_96 word47_96 R_wl
Cwl_48_96 word48_96 gnd C_wl
Rw49_96 word49_96 word48_96 R_wl
Cwl_49_96 word49_96 gnd C_wl
Rw50_96 word50_96 word49_96 R_wl
Cwl_50_96 word50_96 gnd C_wl
Rw51_96 word51_96 word50_96 R_wl
Cwl_51_96 word51_96 gnd C_wl
Rw52_96 word52_96 word51_96 R_wl
Cwl_52_96 word52_96 gnd C_wl
Rw53_96 word53_96 word52_96 R_wl
Cwl_53_96 word53_96 gnd C_wl
Rw54_96 word54_96 word53_96 R_wl
Cwl_54_96 word54_96 gnd C_wl
Rw55_96 word55_96 word54_96 R_wl
Cwl_55_96 word55_96 gnd C_wl
Rw56_96 word56_96 word55_96 R_wl
Cwl_56_96 word56_96 gnd C_wl
Rw57_96 word57_96 word56_96 R_wl
Cwl_57_96 word57_96 gnd C_wl
Rw58_96 word58_96 word57_96 R_wl
Cwl_58_96 word58_96 gnd C_wl
Rw59_96 word59_96 word58_96 R_wl
Cwl_59_96 word59_96 gnd C_wl
Rw60_96 word60_96 word59_96 R_wl
Cwl_60_96 word60_96 gnd C_wl
Rw61_96 word61_96 word60_96 R_wl
Cwl_61_96 word61_96 gnd C_wl
Rw62_96 word62_96 word61_96 R_wl
Cwl_62_96 word62_96 gnd C_wl
Rw63_96 word63_96 word62_96 R_wl
Cwl_63_96 word63_96 gnd C_wl
Rw64_96 word64_96 word63_96 R_wl
Cwl_64_96 word64_96 gnd C_wl
Rw65_96 word65_96 word64_96 R_wl
Cwl_65_96 word65_96 gnd C_wl
Rw66_96 word66_96 word65_96 R_wl
Cwl_66_96 word66_96 gnd C_wl
Rw67_96 word67_96 word66_96 R_wl
Cwl_67_96 word67_96 gnd C_wl
Rw68_96 word68_96 word67_96 R_wl
Cwl_68_96 word68_96 gnd C_wl
Rw69_96 word69_96 word68_96 R_wl
Cwl_69_96 word69_96 gnd C_wl
Rw70_96 word70_96 word69_96 R_wl
Cwl_70_96 word70_96 gnd C_wl
Rw71_96 word71_96 word70_96 R_wl
Cwl_71_96 word71_96 gnd C_wl
Rw72_96 word72_96 word71_96 R_wl
Cwl_72_96 word72_96 gnd C_wl
Rw73_96 word73_96 word72_96 R_wl
Cwl_73_96 word73_96 gnd C_wl
Rw74_96 word74_96 word73_96 R_wl
Cwl_74_96 word74_96 gnd C_wl
Rw75_96 word75_96 word74_96 R_wl
Cwl_75_96 word75_96 gnd C_wl
Rw76_96 word76_96 word75_96 R_wl
Cwl_76_96 word76_96 gnd C_wl
Rw77_96 word77_96 word76_96 R_wl
Cwl_77_96 word77_96 gnd C_wl
Rw78_96 word78_96 word77_96 R_wl
Cwl_78_96 word78_96 gnd C_wl
Rw79_96 word79_96 word78_96 R_wl
Cwl_79_96 word79_96 gnd C_wl
Rw80_96 word80_96 word79_96 R_wl
Cwl_80_96 word80_96 gnd C_wl
Rw81_96 word81_96 word80_96 R_wl
Cwl_81_96 word81_96 gnd C_wl
Rw82_96 word82_96 word81_96 R_wl
Cwl_82_96 word82_96 gnd C_wl
Rw83_96 word83_96 word82_96 R_wl
Cwl_83_96 word83_96 gnd C_wl
Rw84_96 word84_96 word83_96 R_wl
Cwl_84_96 word84_96 gnd C_wl
Rw85_96 word85_96 word84_96 R_wl
Cwl_85_96 word85_96 gnd C_wl
Rw86_96 word86_96 word85_96 R_wl
Cwl_86_96 word86_96 gnd C_wl
Rw87_96 word87_96 word86_96 R_wl
Cwl_87_96 word87_96 gnd C_wl
Rw88_96 word88_96 word87_96 R_wl
Cwl_88_96 word88_96 gnd C_wl
Rw89_96 word89_96 word88_96 R_wl
Cwl_89_96 word89_96 gnd C_wl
Rw90_96 word90_96 word89_96 R_wl
Cwl_90_96 word90_96 gnd C_wl
Rw91_96 word91_96 word90_96 R_wl
Cwl_91_96 word91_96 gnd C_wl
Rw92_96 word92_96 word91_96 R_wl
Cwl_92_96 word92_96 gnd C_wl
Rw93_96 word93_96 word92_96 R_wl
Cwl_93_96 word93_96 gnd C_wl
Rw94_96 word94_96 word93_96 R_wl
Cwl_94_96 word94_96 gnd C_wl
Rw95_96 word95_96 word94_96 R_wl
Cwl_95_96 word95_96 gnd C_wl
Rw96_96 word96_96 word95_96 R_wl
Cwl_96_96 word96_96 gnd C_wl
Rw97_96 word97_96 word96_96 R_wl
Cwl_97_96 word97_96 gnd C_wl
Rw98_96 word98_96 word97_96 R_wl
Cwl_98_96 word98_96 gnd C_wl
Rw99_96 word99_96 word98_96 R_wl
Cwl_99_96 word99_96 gnd C_wl
Vwl_97 word_97 0 0
Rw0_97 word_97 word0_97 R_wl
Cwl_0_97 word0_97 gnd C_wl
Rw1_97 word1_97 word0_97 R_wl
Cwl_1_97 word1_97 gnd C_wl
Rw2_97 word2_97 word1_97 R_wl
Cwl_2_97 word2_97 gnd C_wl
Rw3_97 word3_97 word2_97 R_wl
Cwl_3_97 word3_97 gnd C_wl
Rw4_97 word4_97 word3_97 R_wl
Cwl_4_97 word4_97 gnd C_wl
Rw5_97 word5_97 word4_97 R_wl
Cwl_5_97 word5_97 gnd C_wl
Rw6_97 word6_97 word5_97 R_wl
Cwl_6_97 word6_97 gnd C_wl
Rw7_97 word7_97 word6_97 R_wl
Cwl_7_97 word7_97 gnd C_wl
Rw8_97 word8_97 word7_97 R_wl
Cwl_8_97 word8_97 gnd C_wl
Rw9_97 word9_97 word8_97 R_wl
Cwl_9_97 word9_97 gnd C_wl
Rw10_97 word10_97 word9_97 R_wl
Cwl_10_97 word10_97 gnd C_wl
Rw11_97 word11_97 word10_97 R_wl
Cwl_11_97 word11_97 gnd C_wl
Rw12_97 word12_97 word11_97 R_wl
Cwl_12_97 word12_97 gnd C_wl
Rw13_97 word13_97 word12_97 R_wl
Cwl_13_97 word13_97 gnd C_wl
Rw14_97 word14_97 word13_97 R_wl
Cwl_14_97 word14_97 gnd C_wl
Rw15_97 word15_97 word14_97 R_wl
Cwl_15_97 word15_97 gnd C_wl
Rw16_97 word16_97 word15_97 R_wl
Cwl_16_97 word16_97 gnd C_wl
Rw17_97 word17_97 word16_97 R_wl
Cwl_17_97 word17_97 gnd C_wl
Rw18_97 word18_97 word17_97 R_wl
Cwl_18_97 word18_97 gnd C_wl
Rw19_97 word19_97 word18_97 R_wl
Cwl_19_97 word19_97 gnd C_wl
Rw20_97 word20_97 word19_97 R_wl
Cwl_20_97 word20_97 gnd C_wl
Rw21_97 word21_97 word20_97 R_wl
Cwl_21_97 word21_97 gnd C_wl
Rw22_97 word22_97 word21_97 R_wl
Cwl_22_97 word22_97 gnd C_wl
Rw23_97 word23_97 word22_97 R_wl
Cwl_23_97 word23_97 gnd C_wl
Rw24_97 word24_97 word23_97 R_wl
Cwl_24_97 word24_97 gnd C_wl
Rw25_97 word25_97 word24_97 R_wl
Cwl_25_97 word25_97 gnd C_wl
Rw26_97 word26_97 word25_97 R_wl
Cwl_26_97 word26_97 gnd C_wl
Rw27_97 word27_97 word26_97 R_wl
Cwl_27_97 word27_97 gnd C_wl
Rw28_97 word28_97 word27_97 R_wl
Cwl_28_97 word28_97 gnd C_wl
Rw29_97 word29_97 word28_97 R_wl
Cwl_29_97 word29_97 gnd C_wl
Rw30_97 word30_97 word29_97 R_wl
Cwl_30_97 word30_97 gnd C_wl
Rw31_97 word31_97 word30_97 R_wl
Cwl_31_97 word31_97 gnd C_wl
Rw32_97 word32_97 word31_97 R_wl
Cwl_32_97 word32_97 gnd C_wl
Rw33_97 word33_97 word32_97 R_wl
Cwl_33_97 word33_97 gnd C_wl
Rw34_97 word34_97 word33_97 R_wl
Cwl_34_97 word34_97 gnd C_wl
Rw35_97 word35_97 word34_97 R_wl
Cwl_35_97 word35_97 gnd C_wl
Rw36_97 word36_97 word35_97 R_wl
Cwl_36_97 word36_97 gnd C_wl
Rw37_97 word37_97 word36_97 R_wl
Cwl_37_97 word37_97 gnd C_wl
Rw38_97 word38_97 word37_97 R_wl
Cwl_38_97 word38_97 gnd C_wl
Rw39_97 word39_97 word38_97 R_wl
Cwl_39_97 word39_97 gnd C_wl
Rw40_97 word40_97 word39_97 R_wl
Cwl_40_97 word40_97 gnd C_wl
Rw41_97 word41_97 word40_97 R_wl
Cwl_41_97 word41_97 gnd C_wl
Rw42_97 word42_97 word41_97 R_wl
Cwl_42_97 word42_97 gnd C_wl
Rw43_97 word43_97 word42_97 R_wl
Cwl_43_97 word43_97 gnd C_wl
Rw44_97 word44_97 word43_97 R_wl
Cwl_44_97 word44_97 gnd C_wl
Rw45_97 word45_97 word44_97 R_wl
Cwl_45_97 word45_97 gnd C_wl
Rw46_97 word46_97 word45_97 R_wl
Cwl_46_97 word46_97 gnd C_wl
Rw47_97 word47_97 word46_97 R_wl
Cwl_47_97 word47_97 gnd C_wl
Rw48_97 word48_97 word47_97 R_wl
Cwl_48_97 word48_97 gnd C_wl
Rw49_97 word49_97 word48_97 R_wl
Cwl_49_97 word49_97 gnd C_wl
Rw50_97 word50_97 word49_97 R_wl
Cwl_50_97 word50_97 gnd C_wl
Rw51_97 word51_97 word50_97 R_wl
Cwl_51_97 word51_97 gnd C_wl
Rw52_97 word52_97 word51_97 R_wl
Cwl_52_97 word52_97 gnd C_wl
Rw53_97 word53_97 word52_97 R_wl
Cwl_53_97 word53_97 gnd C_wl
Rw54_97 word54_97 word53_97 R_wl
Cwl_54_97 word54_97 gnd C_wl
Rw55_97 word55_97 word54_97 R_wl
Cwl_55_97 word55_97 gnd C_wl
Rw56_97 word56_97 word55_97 R_wl
Cwl_56_97 word56_97 gnd C_wl
Rw57_97 word57_97 word56_97 R_wl
Cwl_57_97 word57_97 gnd C_wl
Rw58_97 word58_97 word57_97 R_wl
Cwl_58_97 word58_97 gnd C_wl
Rw59_97 word59_97 word58_97 R_wl
Cwl_59_97 word59_97 gnd C_wl
Rw60_97 word60_97 word59_97 R_wl
Cwl_60_97 word60_97 gnd C_wl
Rw61_97 word61_97 word60_97 R_wl
Cwl_61_97 word61_97 gnd C_wl
Rw62_97 word62_97 word61_97 R_wl
Cwl_62_97 word62_97 gnd C_wl
Rw63_97 word63_97 word62_97 R_wl
Cwl_63_97 word63_97 gnd C_wl
Rw64_97 word64_97 word63_97 R_wl
Cwl_64_97 word64_97 gnd C_wl
Rw65_97 word65_97 word64_97 R_wl
Cwl_65_97 word65_97 gnd C_wl
Rw66_97 word66_97 word65_97 R_wl
Cwl_66_97 word66_97 gnd C_wl
Rw67_97 word67_97 word66_97 R_wl
Cwl_67_97 word67_97 gnd C_wl
Rw68_97 word68_97 word67_97 R_wl
Cwl_68_97 word68_97 gnd C_wl
Rw69_97 word69_97 word68_97 R_wl
Cwl_69_97 word69_97 gnd C_wl
Rw70_97 word70_97 word69_97 R_wl
Cwl_70_97 word70_97 gnd C_wl
Rw71_97 word71_97 word70_97 R_wl
Cwl_71_97 word71_97 gnd C_wl
Rw72_97 word72_97 word71_97 R_wl
Cwl_72_97 word72_97 gnd C_wl
Rw73_97 word73_97 word72_97 R_wl
Cwl_73_97 word73_97 gnd C_wl
Rw74_97 word74_97 word73_97 R_wl
Cwl_74_97 word74_97 gnd C_wl
Rw75_97 word75_97 word74_97 R_wl
Cwl_75_97 word75_97 gnd C_wl
Rw76_97 word76_97 word75_97 R_wl
Cwl_76_97 word76_97 gnd C_wl
Rw77_97 word77_97 word76_97 R_wl
Cwl_77_97 word77_97 gnd C_wl
Rw78_97 word78_97 word77_97 R_wl
Cwl_78_97 word78_97 gnd C_wl
Rw79_97 word79_97 word78_97 R_wl
Cwl_79_97 word79_97 gnd C_wl
Rw80_97 word80_97 word79_97 R_wl
Cwl_80_97 word80_97 gnd C_wl
Rw81_97 word81_97 word80_97 R_wl
Cwl_81_97 word81_97 gnd C_wl
Rw82_97 word82_97 word81_97 R_wl
Cwl_82_97 word82_97 gnd C_wl
Rw83_97 word83_97 word82_97 R_wl
Cwl_83_97 word83_97 gnd C_wl
Rw84_97 word84_97 word83_97 R_wl
Cwl_84_97 word84_97 gnd C_wl
Rw85_97 word85_97 word84_97 R_wl
Cwl_85_97 word85_97 gnd C_wl
Rw86_97 word86_97 word85_97 R_wl
Cwl_86_97 word86_97 gnd C_wl
Rw87_97 word87_97 word86_97 R_wl
Cwl_87_97 word87_97 gnd C_wl
Rw88_97 word88_97 word87_97 R_wl
Cwl_88_97 word88_97 gnd C_wl
Rw89_97 word89_97 word88_97 R_wl
Cwl_89_97 word89_97 gnd C_wl
Rw90_97 word90_97 word89_97 R_wl
Cwl_90_97 word90_97 gnd C_wl
Rw91_97 word91_97 word90_97 R_wl
Cwl_91_97 word91_97 gnd C_wl
Rw92_97 word92_97 word91_97 R_wl
Cwl_92_97 word92_97 gnd C_wl
Rw93_97 word93_97 word92_97 R_wl
Cwl_93_97 word93_97 gnd C_wl
Rw94_97 word94_97 word93_97 R_wl
Cwl_94_97 word94_97 gnd C_wl
Rw95_97 word95_97 word94_97 R_wl
Cwl_95_97 word95_97 gnd C_wl
Rw96_97 word96_97 word95_97 R_wl
Cwl_96_97 word96_97 gnd C_wl
Rw97_97 word97_97 word96_97 R_wl
Cwl_97_97 word97_97 gnd C_wl
Rw98_97 word98_97 word97_97 R_wl
Cwl_98_97 word98_97 gnd C_wl
Rw99_97 word99_97 word98_97 R_wl
Cwl_99_97 word99_97 gnd C_wl
Vwl_98 word_98 0 0
Rw0_98 word_98 word0_98 R_wl
Cwl_0_98 word0_98 gnd C_wl
Rw1_98 word1_98 word0_98 R_wl
Cwl_1_98 word1_98 gnd C_wl
Rw2_98 word2_98 word1_98 R_wl
Cwl_2_98 word2_98 gnd C_wl
Rw3_98 word3_98 word2_98 R_wl
Cwl_3_98 word3_98 gnd C_wl
Rw4_98 word4_98 word3_98 R_wl
Cwl_4_98 word4_98 gnd C_wl
Rw5_98 word5_98 word4_98 R_wl
Cwl_5_98 word5_98 gnd C_wl
Rw6_98 word6_98 word5_98 R_wl
Cwl_6_98 word6_98 gnd C_wl
Rw7_98 word7_98 word6_98 R_wl
Cwl_7_98 word7_98 gnd C_wl
Rw8_98 word8_98 word7_98 R_wl
Cwl_8_98 word8_98 gnd C_wl
Rw9_98 word9_98 word8_98 R_wl
Cwl_9_98 word9_98 gnd C_wl
Rw10_98 word10_98 word9_98 R_wl
Cwl_10_98 word10_98 gnd C_wl
Rw11_98 word11_98 word10_98 R_wl
Cwl_11_98 word11_98 gnd C_wl
Rw12_98 word12_98 word11_98 R_wl
Cwl_12_98 word12_98 gnd C_wl
Rw13_98 word13_98 word12_98 R_wl
Cwl_13_98 word13_98 gnd C_wl
Rw14_98 word14_98 word13_98 R_wl
Cwl_14_98 word14_98 gnd C_wl
Rw15_98 word15_98 word14_98 R_wl
Cwl_15_98 word15_98 gnd C_wl
Rw16_98 word16_98 word15_98 R_wl
Cwl_16_98 word16_98 gnd C_wl
Rw17_98 word17_98 word16_98 R_wl
Cwl_17_98 word17_98 gnd C_wl
Rw18_98 word18_98 word17_98 R_wl
Cwl_18_98 word18_98 gnd C_wl
Rw19_98 word19_98 word18_98 R_wl
Cwl_19_98 word19_98 gnd C_wl
Rw20_98 word20_98 word19_98 R_wl
Cwl_20_98 word20_98 gnd C_wl
Rw21_98 word21_98 word20_98 R_wl
Cwl_21_98 word21_98 gnd C_wl
Rw22_98 word22_98 word21_98 R_wl
Cwl_22_98 word22_98 gnd C_wl
Rw23_98 word23_98 word22_98 R_wl
Cwl_23_98 word23_98 gnd C_wl
Rw24_98 word24_98 word23_98 R_wl
Cwl_24_98 word24_98 gnd C_wl
Rw25_98 word25_98 word24_98 R_wl
Cwl_25_98 word25_98 gnd C_wl
Rw26_98 word26_98 word25_98 R_wl
Cwl_26_98 word26_98 gnd C_wl
Rw27_98 word27_98 word26_98 R_wl
Cwl_27_98 word27_98 gnd C_wl
Rw28_98 word28_98 word27_98 R_wl
Cwl_28_98 word28_98 gnd C_wl
Rw29_98 word29_98 word28_98 R_wl
Cwl_29_98 word29_98 gnd C_wl
Rw30_98 word30_98 word29_98 R_wl
Cwl_30_98 word30_98 gnd C_wl
Rw31_98 word31_98 word30_98 R_wl
Cwl_31_98 word31_98 gnd C_wl
Rw32_98 word32_98 word31_98 R_wl
Cwl_32_98 word32_98 gnd C_wl
Rw33_98 word33_98 word32_98 R_wl
Cwl_33_98 word33_98 gnd C_wl
Rw34_98 word34_98 word33_98 R_wl
Cwl_34_98 word34_98 gnd C_wl
Rw35_98 word35_98 word34_98 R_wl
Cwl_35_98 word35_98 gnd C_wl
Rw36_98 word36_98 word35_98 R_wl
Cwl_36_98 word36_98 gnd C_wl
Rw37_98 word37_98 word36_98 R_wl
Cwl_37_98 word37_98 gnd C_wl
Rw38_98 word38_98 word37_98 R_wl
Cwl_38_98 word38_98 gnd C_wl
Rw39_98 word39_98 word38_98 R_wl
Cwl_39_98 word39_98 gnd C_wl
Rw40_98 word40_98 word39_98 R_wl
Cwl_40_98 word40_98 gnd C_wl
Rw41_98 word41_98 word40_98 R_wl
Cwl_41_98 word41_98 gnd C_wl
Rw42_98 word42_98 word41_98 R_wl
Cwl_42_98 word42_98 gnd C_wl
Rw43_98 word43_98 word42_98 R_wl
Cwl_43_98 word43_98 gnd C_wl
Rw44_98 word44_98 word43_98 R_wl
Cwl_44_98 word44_98 gnd C_wl
Rw45_98 word45_98 word44_98 R_wl
Cwl_45_98 word45_98 gnd C_wl
Rw46_98 word46_98 word45_98 R_wl
Cwl_46_98 word46_98 gnd C_wl
Rw47_98 word47_98 word46_98 R_wl
Cwl_47_98 word47_98 gnd C_wl
Rw48_98 word48_98 word47_98 R_wl
Cwl_48_98 word48_98 gnd C_wl
Rw49_98 word49_98 word48_98 R_wl
Cwl_49_98 word49_98 gnd C_wl
Rw50_98 word50_98 word49_98 R_wl
Cwl_50_98 word50_98 gnd C_wl
Rw51_98 word51_98 word50_98 R_wl
Cwl_51_98 word51_98 gnd C_wl
Rw52_98 word52_98 word51_98 R_wl
Cwl_52_98 word52_98 gnd C_wl
Rw53_98 word53_98 word52_98 R_wl
Cwl_53_98 word53_98 gnd C_wl
Rw54_98 word54_98 word53_98 R_wl
Cwl_54_98 word54_98 gnd C_wl
Rw55_98 word55_98 word54_98 R_wl
Cwl_55_98 word55_98 gnd C_wl
Rw56_98 word56_98 word55_98 R_wl
Cwl_56_98 word56_98 gnd C_wl
Rw57_98 word57_98 word56_98 R_wl
Cwl_57_98 word57_98 gnd C_wl
Rw58_98 word58_98 word57_98 R_wl
Cwl_58_98 word58_98 gnd C_wl
Rw59_98 word59_98 word58_98 R_wl
Cwl_59_98 word59_98 gnd C_wl
Rw60_98 word60_98 word59_98 R_wl
Cwl_60_98 word60_98 gnd C_wl
Rw61_98 word61_98 word60_98 R_wl
Cwl_61_98 word61_98 gnd C_wl
Rw62_98 word62_98 word61_98 R_wl
Cwl_62_98 word62_98 gnd C_wl
Rw63_98 word63_98 word62_98 R_wl
Cwl_63_98 word63_98 gnd C_wl
Rw64_98 word64_98 word63_98 R_wl
Cwl_64_98 word64_98 gnd C_wl
Rw65_98 word65_98 word64_98 R_wl
Cwl_65_98 word65_98 gnd C_wl
Rw66_98 word66_98 word65_98 R_wl
Cwl_66_98 word66_98 gnd C_wl
Rw67_98 word67_98 word66_98 R_wl
Cwl_67_98 word67_98 gnd C_wl
Rw68_98 word68_98 word67_98 R_wl
Cwl_68_98 word68_98 gnd C_wl
Rw69_98 word69_98 word68_98 R_wl
Cwl_69_98 word69_98 gnd C_wl
Rw70_98 word70_98 word69_98 R_wl
Cwl_70_98 word70_98 gnd C_wl
Rw71_98 word71_98 word70_98 R_wl
Cwl_71_98 word71_98 gnd C_wl
Rw72_98 word72_98 word71_98 R_wl
Cwl_72_98 word72_98 gnd C_wl
Rw73_98 word73_98 word72_98 R_wl
Cwl_73_98 word73_98 gnd C_wl
Rw74_98 word74_98 word73_98 R_wl
Cwl_74_98 word74_98 gnd C_wl
Rw75_98 word75_98 word74_98 R_wl
Cwl_75_98 word75_98 gnd C_wl
Rw76_98 word76_98 word75_98 R_wl
Cwl_76_98 word76_98 gnd C_wl
Rw77_98 word77_98 word76_98 R_wl
Cwl_77_98 word77_98 gnd C_wl
Rw78_98 word78_98 word77_98 R_wl
Cwl_78_98 word78_98 gnd C_wl
Rw79_98 word79_98 word78_98 R_wl
Cwl_79_98 word79_98 gnd C_wl
Rw80_98 word80_98 word79_98 R_wl
Cwl_80_98 word80_98 gnd C_wl
Rw81_98 word81_98 word80_98 R_wl
Cwl_81_98 word81_98 gnd C_wl
Rw82_98 word82_98 word81_98 R_wl
Cwl_82_98 word82_98 gnd C_wl
Rw83_98 word83_98 word82_98 R_wl
Cwl_83_98 word83_98 gnd C_wl
Rw84_98 word84_98 word83_98 R_wl
Cwl_84_98 word84_98 gnd C_wl
Rw85_98 word85_98 word84_98 R_wl
Cwl_85_98 word85_98 gnd C_wl
Rw86_98 word86_98 word85_98 R_wl
Cwl_86_98 word86_98 gnd C_wl
Rw87_98 word87_98 word86_98 R_wl
Cwl_87_98 word87_98 gnd C_wl
Rw88_98 word88_98 word87_98 R_wl
Cwl_88_98 word88_98 gnd C_wl
Rw89_98 word89_98 word88_98 R_wl
Cwl_89_98 word89_98 gnd C_wl
Rw90_98 word90_98 word89_98 R_wl
Cwl_90_98 word90_98 gnd C_wl
Rw91_98 word91_98 word90_98 R_wl
Cwl_91_98 word91_98 gnd C_wl
Rw92_98 word92_98 word91_98 R_wl
Cwl_92_98 word92_98 gnd C_wl
Rw93_98 word93_98 word92_98 R_wl
Cwl_93_98 word93_98 gnd C_wl
Rw94_98 word94_98 word93_98 R_wl
Cwl_94_98 word94_98 gnd C_wl
Rw95_98 word95_98 word94_98 R_wl
Cwl_95_98 word95_98 gnd C_wl
Rw96_98 word96_98 word95_98 R_wl
Cwl_96_98 word96_98 gnd C_wl
Rw97_98 word97_98 word96_98 R_wl
Cwl_97_98 word97_98 gnd C_wl
Rw98_98 word98_98 word97_98 R_wl
Cwl_98_98 word98_98 gnd C_wl
Rw99_98 word99_98 word98_98 R_wl
Cwl_99_98 word99_98 gnd C_wl
Vwl_99 word_99 gnd pwl 0 0 (16n) 0 (17n) 1.8 50n 1.8 (51n) 0 
Rw0_99 word_99 word0_99 R_wl
Cwl_0_99 word0_99 gnd C_wl
Rw1_99 word1_99 word0_99 R_wl
Cwl_1_99 word1_99 gnd C_wl
Rw2_99 word2_99 word1_99 R_wl
Cwl_2_99 word2_99 gnd C_wl
Rw3_99 word3_99 word2_99 R_wl
Cwl_3_99 word3_99 gnd C_wl
Rw4_99 word4_99 word3_99 R_wl
Cwl_4_99 word4_99 gnd C_wl
Rw5_99 word5_99 word4_99 R_wl
Cwl_5_99 word5_99 gnd C_wl
Rw6_99 word6_99 word5_99 R_wl
Cwl_6_99 word6_99 gnd C_wl
Rw7_99 word7_99 word6_99 R_wl
Cwl_7_99 word7_99 gnd C_wl
Rw8_99 word8_99 word7_99 R_wl
Cwl_8_99 word8_99 gnd C_wl
Rw9_99 word9_99 word8_99 R_wl
Cwl_9_99 word9_99 gnd C_wl
Rw10_99 word10_99 word9_99 R_wl
Cwl_10_99 word10_99 gnd C_wl
Rw11_99 word11_99 word10_99 R_wl
Cwl_11_99 word11_99 gnd C_wl
Rw12_99 word12_99 word11_99 R_wl
Cwl_12_99 word12_99 gnd C_wl
Rw13_99 word13_99 word12_99 R_wl
Cwl_13_99 word13_99 gnd C_wl
Rw14_99 word14_99 word13_99 R_wl
Cwl_14_99 word14_99 gnd C_wl
Rw15_99 word15_99 word14_99 R_wl
Cwl_15_99 word15_99 gnd C_wl
Rw16_99 word16_99 word15_99 R_wl
Cwl_16_99 word16_99 gnd C_wl
Rw17_99 word17_99 word16_99 R_wl
Cwl_17_99 word17_99 gnd C_wl
Rw18_99 word18_99 word17_99 R_wl
Cwl_18_99 word18_99 gnd C_wl
Rw19_99 word19_99 word18_99 R_wl
Cwl_19_99 word19_99 gnd C_wl
Rw20_99 word20_99 word19_99 R_wl
Cwl_20_99 word20_99 gnd C_wl
Rw21_99 word21_99 word20_99 R_wl
Cwl_21_99 word21_99 gnd C_wl
Rw22_99 word22_99 word21_99 R_wl
Cwl_22_99 word22_99 gnd C_wl
Rw23_99 word23_99 word22_99 R_wl
Cwl_23_99 word23_99 gnd C_wl
Rw24_99 word24_99 word23_99 R_wl
Cwl_24_99 word24_99 gnd C_wl
Rw25_99 word25_99 word24_99 R_wl
Cwl_25_99 word25_99 gnd C_wl
Rw26_99 word26_99 word25_99 R_wl
Cwl_26_99 word26_99 gnd C_wl
Rw27_99 word27_99 word26_99 R_wl
Cwl_27_99 word27_99 gnd C_wl
Rw28_99 word28_99 word27_99 R_wl
Cwl_28_99 word28_99 gnd C_wl
Rw29_99 word29_99 word28_99 R_wl
Cwl_29_99 word29_99 gnd C_wl
Rw30_99 word30_99 word29_99 R_wl
Cwl_30_99 word30_99 gnd C_wl
Rw31_99 word31_99 word30_99 R_wl
Cwl_31_99 word31_99 gnd C_wl
Rw32_99 word32_99 word31_99 R_wl
Cwl_32_99 word32_99 gnd C_wl
Rw33_99 word33_99 word32_99 R_wl
Cwl_33_99 word33_99 gnd C_wl
Rw34_99 word34_99 word33_99 R_wl
Cwl_34_99 word34_99 gnd C_wl
Rw35_99 word35_99 word34_99 R_wl
Cwl_35_99 word35_99 gnd C_wl
Rw36_99 word36_99 word35_99 R_wl
Cwl_36_99 word36_99 gnd C_wl
Rw37_99 word37_99 word36_99 R_wl
Cwl_37_99 word37_99 gnd C_wl
Rw38_99 word38_99 word37_99 R_wl
Cwl_38_99 word38_99 gnd C_wl
Rw39_99 word39_99 word38_99 R_wl
Cwl_39_99 word39_99 gnd C_wl
Rw40_99 word40_99 word39_99 R_wl
Cwl_40_99 word40_99 gnd C_wl
Rw41_99 word41_99 word40_99 R_wl
Cwl_41_99 word41_99 gnd C_wl
Rw42_99 word42_99 word41_99 R_wl
Cwl_42_99 word42_99 gnd C_wl
Rw43_99 word43_99 word42_99 R_wl
Cwl_43_99 word43_99 gnd C_wl
Rw44_99 word44_99 word43_99 R_wl
Cwl_44_99 word44_99 gnd C_wl
Rw45_99 word45_99 word44_99 R_wl
Cwl_45_99 word45_99 gnd C_wl
Rw46_99 word46_99 word45_99 R_wl
Cwl_46_99 word46_99 gnd C_wl
Rw47_99 word47_99 word46_99 R_wl
Cwl_47_99 word47_99 gnd C_wl
Rw48_99 word48_99 word47_99 R_wl
Cwl_48_99 word48_99 gnd C_wl
Rw49_99 word49_99 word48_99 R_wl
Cwl_49_99 word49_99 gnd C_wl
Rw50_99 word50_99 word49_99 R_wl
Cwl_50_99 word50_99 gnd C_wl
Rw51_99 word51_99 word50_99 R_wl
Cwl_51_99 word51_99 gnd C_wl
Rw52_99 word52_99 word51_99 R_wl
Cwl_52_99 word52_99 gnd C_wl
Rw53_99 word53_99 word52_99 R_wl
Cwl_53_99 word53_99 gnd C_wl
Rw54_99 word54_99 word53_99 R_wl
Cwl_54_99 word54_99 gnd C_wl
Rw55_99 word55_99 word54_99 R_wl
Cwl_55_99 word55_99 gnd C_wl
Rw56_99 word56_99 word55_99 R_wl
Cwl_56_99 word56_99 gnd C_wl
Rw57_99 word57_99 word56_99 R_wl
Cwl_57_99 word57_99 gnd C_wl
Rw58_99 word58_99 word57_99 R_wl
Cwl_58_99 word58_99 gnd C_wl
Rw59_99 word59_99 word58_99 R_wl
Cwl_59_99 word59_99 gnd C_wl
Rw60_99 word60_99 word59_99 R_wl
Cwl_60_99 word60_99 gnd C_wl
Rw61_99 word61_99 word60_99 R_wl
Cwl_61_99 word61_99 gnd C_wl
Rw62_99 word62_99 word61_99 R_wl
Cwl_62_99 word62_99 gnd C_wl
Rw63_99 word63_99 word62_99 R_wl
Cwl_63_99 word63_99 gnd C_wl
Rw64_99 word64_99 word63_99 R_wl
Cwl_64_99 word64_99 gnd C_wl
Rw65_99 word65_99 word64_99 R_wl
Cwl_65_99 word65_99 gnd C_wl
Rw66_99 word66_99 word65_99 R_wl
Cwl_66_99 word66_99 gnd C_wl
Rw67_99 word67_99 word66_99 R_wl
Cwl_67_99 word67_99 gnd C_wl
Rw68_99 word68_99 word67_99 R_wl
Cwl_68_99 word68_99 gnd C_wl
Rw69_99 word69_99 word68_99 R_wl
Cwl_69_99 word69_99 gnd C_wl
Rw70_99 word70_99 word69_99 R_wl
Cwl_70_99 word70_99 gnd C_wl
Rw71_99 word71_99 word70_99 R_wl
Cwl_71_99 word71_99 gnd C_wl
Rw72_99 word72_99 word71_99 R_wl
Cwl_72_99 word72_99 gnd C_wl
Rw73_99 word73_99 word72_99 R_wl
Cwl_73_99 word73_99 gnd C_wl
Rw74_99 word74_99 word73_99 R_wl
Cwl_74_99 word74_99 gnd C_wl
Rw75_99 word75_99 word74_99 R_wl
Cwl_75_99 word75_99 gnd C_wl
Rw76_99 word76_99 word75_99 R_wl
Cwl_76_99 word76_99 gnd C_wl
Rw77_99 word77_99 word76_99 R_wl
Cwl_77_99 word77_99 gnd C_wl
Rw78_99 word78_99 word77_99 R_wl
Cwl_78_99 word78_99 gnd C_wl
Rw79_99 word79_99 word78_99 R_wl
Cwl_79_99 word79_99 gnd C_wl
Rw80_99 word80_99 word79_99 R_wl
Cwl_80_99 word80_99 gnd C_wl
Rw81_99 word81_99 word80_99 R_wl
Cwl_81_99 word81_99 gnd C_wl
Rw82_99 word82_99 word81_99 R_wl
Cwl_82_99 word82_99 gnd C_wl
Rw83_99 word83_99 word82_99 R_wl
Cwl_83_99 word83_99 gnd C_wl
Rw84_99 word84_99 word83_99 R_wl
Cwl_84_99 word84_99 gnd C_wl
Rw85_99 word85_99 word84_99 R_wl
Cwl_85_99 word85_99 gnd C_wl
Rw86_99 word86_99 word85_99 R_wl
Cwl_86_99 word86_99 gnd C_wl
Rw87_99 word87_99 word86_99 R_wl
Cwl_87_99 word87_99 gnd C_wl
Rw88_99 word88_99 word87_99 R_wl
Cwl_88_99 word88_99 gnd C_wl
Rw89_99 word89_99 word88_99 R_wl
Cwl_89_99 word89_99 gnd C_wl
Rw90_99 word90_99 word89_99 R_wl
Cwl_90_99 word90_99 gnd C_wl
Rw91_99 word91_99 word90_99 R_wl
Cwl_91_99 word91_99 gnd C_wl
Rw92_99 word92_99 word91_99 R_wl
Cwl_92_99 word92_99 gnd C_wl
Rw93_99 word93_99 word92_99 R_wl
Cwl_93_99 word93_99 gnd C_wl
Rw94_99 word94_99 word93_99 R_wl
Cwl_94_99 word94_99 gnd C_wl
Rw95_99 word95_99 word94_99 R_wl
Cwl_95_99 word95_99 gnd C_wl
Rw96_99 word96_99 word95_99 R_wl
Cwl_96_99 word96_99 gnd C_wl
Rw97_99 word97_99 word96_99 R_wl
Cwl_97_99 word97_99 gnd C_wl
Rw98_99 word98_99 word97_99 R_wl
Cwl_98_99 word98_99 gnd C_wl
Rw99_99 word99_99 word98_99 R_wl
Cwl_99_99 word99_99 gnd C_wl
*Column access, activates at 110n
Vcol_write_0 col_write_0 gnd dc 0
Vcol_read_0 col_read_0 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_1 col_write_1 gnd dc 0
Vcol_read_1 col_read_1 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_2 col_write_2 gnd dc 0
Vcol_read_2 col_read_2 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_3 col_write_3 gnd dc 0
Vcol_read_3 col_read_3 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_4 col_write_4 gnd dc 0
Vcol_read_4 col_read_4 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_5 col_write_5 gnd dc 0
Vcol_read_5 col_read_5 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_6 col_write_6 gnd dc 0
Vcol_read_6 col_read_6 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_7 col_write_7 gnd dc 0
Vcol_read_7 col_read_7 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_8 col_write_8 gnd dc 0
Vcol_read_8 col_read_8 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_9 col_write_9 gnd dc 0
Vcol_read_9 col_read_9 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_10 col_write_10 gnd dc 0
Vcol_read_10 col_read_10 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_11 col_write_11 gnd dc 0
Vcol_read_11 col_read_11 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_12 col_write_12 gnd dc 0
Vcol_read_12 col_read_12 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_13 col_write_13 gnd dc 0
Vcol_read_13 col_read_13 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_14 col_write_14 gnd dc 0
Vcol_read_14 col_read_14 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_15 col_write_15 gnd dc 0
Vcol_read_15 col_read_15 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_16 col_write_16 gnd dc 0
Vcol_read_16 col_read_16 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_17 col_write_17 gnd dc 0
Vcol_read_17 col_read_17 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_18 col_write_18 gnd dc 0
Vcol_read_18 col_read_18 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_19 col_write_19 gnd dc 0
Vcol_read_19 col_read_19 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_20 col_write_20 gnd dc 0
Vcol_read_20 col_read_20 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_21 col_write_21 gnd dc 0
Vcol_read_21 col_read_21 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_22 col_write_22 gnd dc 0
Vcol_read_22 col_read_22 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_23 col_write_23 gnd dc 0
Vcol_read_23 col_read_23 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_24 col_write_24 gnd dc 0
Vcol_read_24 col_read_24 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_25 col_write_25 gnd dc 0
Vcol_read_25 col_read_25 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_26 col_write_26 gnd dc 0
Vcol_read_26 col_read_26 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_27 col_write_27 gnd dc 0
Vcol_read_27 col_read_27 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_28 col_write_28 gnd dc 0
Vcol_read_28 col_read_28 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_29 col_write_29 gnd dc 0
Vcol_read_29 col_read_29 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_30 col_write_30 gnd dc 0
Vcol_read_30 col_read_30 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_31 col_write_31 gnd dc 0
Vcol_read_31 col_read_31 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_32 col_write_32 gnd dc 0
Vcol_read_32 col_read_32 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_33 col_write_33 gnd dc 0
Vcol_read_33 col_read_33 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_34 col_write_34 gnd dc 0
Vcol_read_34 col_read_34 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_35 col_write_35 gnd dc 0
Vcol_read_35 col_read_35 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_36 col_write_36 gnd dc 0
Vcol_read_36 col_read_36 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_37 col_write_37 gnd dc 0
Vcol_read_37 col_read_37 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_38 col_write_38 gnd dc 0
Vcol_read_38 col_read_38 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_39 col_write_39 gnd dc 0
Vcol_read_39 col_read_39 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_40 col_write_40 gnd dc 0
Vcol_read_40 col_read_40 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_41 col_write_41 gnd dc 0
Vcol_read_41 col_read_41 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_42 col_write_42 gnd dc 0
Vcol_read_42 col_read_42 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_43 col_write_43 gnd dc 0
Vcol_read_43 col_read_43 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_44 col_write_44 gnd dc 0
Vcol_read_44 col_read_44 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_45 col_write_45 gnd dc 0
Vcol_read_45 col_read_45 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_46 col_write_46 gnd dc 0
Vcol_read_46 col_read_46 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_47 col_write_47 gnd dc 0
Vcol_read_47 col_read_47 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_48 col_write_48 gnd dc 0
Vcol_read_48 col_read_48 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_49 col_write_49 gnd dc 0
Vcol_read_49 col_read_49 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_50 col_write_50 gnd dc 0
Vcol_read_50 col_read_50 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_51 col_write_51 gnd dc 0
Vcol_read_51 col_read_51 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_52 col_write_52 gnd dc 0
Vcol_read_52 col_read_52 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_53 col_write_53 gnd dc 0
Vcol_read_53 col_read_53 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_54 col_write_54 gnd dc 0
Vcol_read_54 col_read_54 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_55 col_write_55 gnd dc 0
Vcol_read_55 col_read_55 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_56 col_write_56 gnd dc 0
Vcol_read_56 col_read_56 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_57 col_write_57 gnd dc 0
Vcol_read_57 col_read_57 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_58 col_write_58 gnd dc 0
Vcol_read_58 col_read_58 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_59 col_write_59 gnd dc 0
Vcol_read_59 col_read_59 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_60 col_write_60 gnd dc 0
Vcol_read_60 col_read_60 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_61 col_write_61 gnd dc 0
Vcol_read_61 col_read_61 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_62 col_write_62 gnd dc 0
Vcol_read_62 col_read_62 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_63 col_write_63 gnd dc 0
Vcol_read_63 col_read_63 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_64 col_write_64 gnd dc 0
Vcol_read_64 col_read_64 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_65 col_write_65 gnd dc 0
Vcol_read_65 col_read_65 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_66 col_write_66 gnd dc 0
Vcol_read_66 col_read_66 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_67 col_write_67 gnd dc 0
Vcol_read_67 col_read_67 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_68 col_write_68 gnd dc 0
Vcol_read_68 col_read_68 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_69 col_write_69 gnd dc 0
Vcol_read_69 col_read_69 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_70 col_write_70 gnd dc 0
Vcol_read_70 col_read_70 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_71 col_write_71 gnd dc 0
Vcol_read_71 col_read_71 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_72 col_write_72 gnd dc 0
Vcol_read_72 col_read_72 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_73 col_write_73 gnd dc 0
Vcol_read_73 col_read_73 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_74 col_write_74 gnd dc 0
Vcol_read_74 col_read_74 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_75 col_write_75 gnd dc 0
Vcol_read_75 col_read_75 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_76 col_write_76 gnd dc 0
Vcol_read_76 col_read_76 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_77 col_write_77 gnd dc 0
Vcol_read_77 col_read_77 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_78 col_write_78 gnd dc 0
Vcol_read_78 col_read_78 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_79 col_write_79 gnd dc 0
Vcol_read_79 col_read_79 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_80 col_write_80 gnd dc 0
Vcol_read_80 col_read_80 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_81 col_write_81 gnd dc 0
Vcol_read_81 col_read_81 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_82 col_write_82 gnd dc 0
Vcol_read_82 col_read_82 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_83 col_write_83 gnd dc 0
Vcol_read_83 col_read_83 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_84 col_write_84 gnd dc 0
Vcol_read_84 col_read_84 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_85 col_write_85 gnd dc 0
Vcol_read_85 col_read_85 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_86 col_write_86 gnd dc 0
Vcol_read_86 col_read_86 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_87 col_write_87 gnd dc 0
Vcol_read_87 col_read_87 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_88 col_write_88 gnd dc 0
Vcol_read_88 col_read_88 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_89 col_write_89 gnd dc 0
Vcol_read_89 col_read_89 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_90 col_write_90 gnd dc 0
Vcol_read_90 col_read_90 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_91 col_write_91 gnd dc 0
Vcol_read_91 col_read_91 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_92 col_write_92 gnd dc 0
Vcol_read_92 col_read_92 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_93 col_write_93 gnd dc 0
Vcol_read_93 col_read_93 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_94 col_write_94 gnd dc 0
Vcol_read_94 col_read_94 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_95 col_write_95 gnd dc 0
Vcol_read_95 col_read_95 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_96 col_write_96 gnd dc 0
Vcol_read_96 col_read_96 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_97 col_write_97 gnd dc 0
Vcol_read_97 col_read_97 gnd dc 1.8
*Column access, activates at 110n
Vcol_write_98 col_write_98 gnd dc 0
Vcol_read_98 col_read_98 gnd dc 1.8
*Column access, activates at 110n
Vcol_read_99 col_read_99 gnd pwl 0 1.8 (17n) 1.8 (18n) 0 50n 0 (51n) 1.8
Vcol_write_99 col_write_99 gnd pwl 0 0 (17n) 0 (18n) 1.8 50n 1.8 (51n) 0
*Precharge, activates at 10n
Vpc_0 pc_0 gnd dc 1.8
*Precharge, activates at 10n
Vpc_1 pc_1 gnd dc 1.8
*Precharge, activates at 10n
Vpc_2 pc_2 gnd dc 1.8
*Precharge, activates at 10n
Vpc_3 pc_3 gnd dc 1.8
*Precharge, activates at 10n
Vpc_4 pc_4 gnd dc 1.8
*Precharge, activates at 10n
Vpc_5 pc_5 gnd dc 1.8
*Precharge, activates at 10n
Vpc_6 pc_6 gnd dc 1.8
*Precharge, activates at 10n
Vpc_7 pc_7 gnd dc 1.8
*Precharge, activates at 10n
Vpc_8 pc_8 gnd dc 1.8
*Precharge, activates at 10n
Vpc_9 pc_9 gnd dc 1.8
*Precharge, activates at 10n
Vpc_10 pc_10 gnd dc 1.8
*Precharge, activates at 10n
Vpc_11 pc_11 gnd dc 1.8
*Precharge, activates at 10n
Vpc_12 pc_12 gnd dc 1.8
*Precharge, activates at 10n
Vpc_13 pc_13 gnd dc 1.8
*Precharge, activates at 10n
Vpc_14 pc_14 gnd dc 1.8
*Precharge, activates at 10n
Vpc_15 pc_15 gnd dc 1.8
*Precharge, activates at 10n
Vpc_16 pc_16 gnd dc 1.8
*Precharge, activates at 10n
Vpc_17 pc_17 gnd dc 1.8
*Precharge, activates at 10n
Vpc_18 pc_18 gnd dc 1.8
*Precharge, activates at 10n
Vpc_19 pc_19 gnd dc 1.8
*Precharge, activates at 10n
Vpc_20 pc_20 gnd dc 1.8
*Precharge, activates at 10n
Vpc_21 pc_21 gnd dc 1.8
*Precharge, activates at 10n
Vpc_22 pc_22 gnd dc 1.8
*Precharge, activates at 10n
Vpc_23 pc_23 gnd dc 1.8
*Precharge, activates at 10n
Vpc_24 pc_24 gnd dc 1.8
*Precharge, activates at 10n
Vpc_25 pc_25 gnd dc 1.8
*Precharge, activates at 10n
Vpc_26 pc_26 gnd dc 1.8
*Precharge, activates at 10n
Vpc_27 pc_27 gnd dc 1.8
*Precharge, activates at 10n
Vpc_28 pc_28 gnd dc 1.8
*Precharge, activates at 10n
Vpc_29 pc_29 gnd dc 1.8
*Precharge, activates at 10n
Vpc_30 pc_30 gnd dc 1.8
*Precharge, activates at 10n
Vpc_31 pc_31 gnd dc 1.8
*Precharge, activates at 10n
Vpc_32 pc_32 gnd dc 1.8
*Precharge, activates at 10n
Vpc_33 pc_33 gnd dc 1.8
*Precharge, activates at 10n
Vpc_34 pc_34 gnd dc 1.8
*Precharge, activates at 10n
Vpc_35 pc_35 gnd dc 1.8
*Precharge, activates at 10n
Vpc_36 pc_36 gnd dc 1.8
*Precharge, activates at 10n
Vpc_37 pc_37 gnd dc 1.8
*Precharge, activates at 10n
Vpc_38 pc_38 gnd dc 1.8
*Precharge, activates at 10n
Vpc_39 pc_39 gnd dc 1.8
*Precharge, activates at 10n
Vpc_40 pc_40 gnd dc 1.8
*Precharge, activates at 10n
Vpc_41 pc_41 gnd dc 1.8
*Precharge, activates at 10n
Vpc_42 pc_42 gnd dc 1.8
*Precharge, activates at 10n
Vpc_43 pc_43 gnd dc 1.8
*Precharge, activates at 10n
Vpc_44 pc_44 gnd dc 1.8
*Precharge, activates at 10n
Vpc_45 pc_45 gnd dc 1.8
*Precharge, activates at 10n
Vpc_46 pc_46 gnd dc 1.8
*Precharge, activates at 10n
Vpc_47 pc_47 gnd dc 1.8
*Precharge, activates at 10n
Vpc_48 pc_48 gnd dc 1.8
*Precharge, activates at 10n
Vpc_49 pc_49 gnd dc 1.8
*Precharge, activates at 10n
Vpc_50 pc_50 gnd dc 1.8
*Precharge, activates at 10n
Vpc_51 pc_51 gnd dc 1.8
*Precharge, activates at 10n
Vpc_52 pc_52 gnd dc 1.8
*Precharge, activates at 10n
Vpc_53 pc_53 gnd dc 1.8
*Precharge, activates at 10n
Vpc_54 pc_54 gnd dc 1.8
*Precharge, activates at 10n
Vpc_55 pc_55 gnd dc 1.8
*Precharge, activates at 10n
Vpc_56 pc_56 gnd dc 1.8
*Precharge, activates at 10n
Vpc_57 pc_57 gnd dc 1.8
*Precharge, activates at 10n
Vpc_58 pc_58 gnd dc 1.8
*Precharge, activates at 10n
Vpc_59 pc_59 gnd dc 1.8
*Precharge, activates at 10n
Vpc_60 pc_60 gnd dc 1.8
*Precharge, activates at 10n
Vpc_61 pc_61 gnd dc 1.8
*Precharge, activates at 10n
Vpc_62 pc_62 gnd dc 1.8
*Precharge, activates at 10n
Vpc_63 pc_63 gnd dc 1.8
*Precharge, activates at 10n
Vpc_64 pc_64 gnd dc 1.8
*Precharge, activates at 10n
Vpc_65 pc_65 gnd dc 1.8
*Precharge, activates at 10n
Vpc_66 pc_66 gnd dc 1.8
*Precharge, activates at 10n
Vpc_67 pc_67 gnd dc 1.8
*Precharge, activates at 10n
Vpc_68 pc_68 gnd dc 1.8
*Precharge, activates at 10n
Vpc_69 pc_69 gnd dc 1.8
*Precharge, activates at 10n
Vpc_70 pc_70 gnd dc 1.8
*Precharge, activates at 10n
Vpc_71 pc_71 gnd dc 1.8
*Precharge, activates at 10n
Vpc_72 pc_72 gnd dc 1.8
*Precharge, activates at 10n
Vpc_73 pc_73 gnd dc 1.8
*Precharge, activates at 10n
Vpc_74 pc_74 gnd dc 1.8
*Precharge, activates at 10n
Vpc_75 pc_75 gnd dc 1.8
*Precharge, activates at 10n
Vpc_76 pc_76 gnd dc 1.8
*Precharge, activates at 10n
Vpc_77 pc_77 gnd dc 1.8
*Precharge, activates at 10n
Vpc_78 pc_78 gnd dc 1.8
*Precharge, activates at 10n
Vpc_79 pc_79 gnd dc 1.8
*Precharge, activates at 10n
Vpc_80 pc_80 gnd dc 1.8
*Precharge, activates at 10n
Vpc_81 pc_81 gnd dc 1.8
*Precharge, activates at 10n
Vpc_82 pc_82 gnd dc 1.8
*Precharge, activates at 10n
Vpc_83 pc_83 gnd dc 1.8
*Precharge, activates at 10n
Vpc_84 pc_84 gnd dc 1.8
*Precharge, activates at 10n
Vpc_85 pc_85 gnd dc 1.8
*Precharge, activates at 10n
Vpc_86 pc_86 gnd dc 1.8
*Precharge, activates at 10n
Vpc_87 pc_87 gnd dc 1.8
*Precharge, activates at 10n
Vpc_88 pc_88 gnd dc 1.8
*Precharge, activates at 10n
Vpc_89 pc_89 gnd dc 1.8
*Precharge, activates at 10n
Vpc_90 pc_90 gnd dc 1.8
*Precharge, activates at 10n
Vpc_91 pc_91 gnd dc 1.8
*Precharge, activates at 10n
Vpc_92 pc_92 gnd dc 1.8
*Precharge, activates at 10n
Vpc_93 pc_93 gnd dc 1.8
*Precharge, activates at 10n
Vpc_94 pc_94 gnd dc 1.8
*Precharge, activates at 10n
Vpc_95 pc_95 gnd dc 1.8
*Precharge, activates at 10n
Vpc_96 pc_96 gnd dc 1.8
*Precharge, activates at 10n
Vpc_97 pc_97 gnd dc 1.8
*Precharge, activates at 10n
Vpc_98 pc_98 gnd dc 1.8
*Precharge, activates at 10n
Vpc_99 pc_99 gnd pwl 0 1.8 10n 1.8 11n 0 14n 0 15n 1.8
*Sense amp bias supply
Vsa sa_vcs gnd dc 0.7
.param R_bl=0.5
.param C_bl=3.789f
Rb_0_0 bit_0_0 bit_0_1 R_bl
Rbb_0_0 bitb_0_0 bitb_0_1 R_bl
Cb_0_0 bit_0_0 gnd C_bl
Cbb_0_0 bitb_0_0 gnd C_bl
Rb_0_1 bit_0_1 bit_0_2 R_bl
Rbb_0_1 bitb_0_1 bitb_0_2 R_bl
Cb_0_1 bit_0_1 gnd C_bl
Cbb_0_1 bitb_0_1 gnd C_bl
Rb_0_2 bit_0_2 bit_0_3 R_bl
Rbb_0_2 bitb_0_2 bitb_0_3 R_bl
Cb_0_2 bit_0_2 gnd C_bl
Cbb_0_2 bitb_0_2 gnd C_bl
Rb_0_3 bit_0_3 bit_0_4 R_bl
Rbb_0_3 bitb_0_3 bitb_0_4 R_bl
Cb_0_3 bit_0_3 gnd C_bl
Cbb_0_3 bitb_0_3 gnd C_bl
Rb_0_4 bit_0_4 bit_0_5 R_bl
Rbb_0_4 bitb_0_4 bitb_0_5 R_bl
Cb_0_4 bit_0_4 gnd C_bl
Cbb_0_4 bitb_0_4 gnd C_bl
Rb_0_5 bit_0_5 bit_0_6 R_bl
Rbb_0_5 bitb_0_5 bitb_0_6 R_bl
Cb_0_5 bit_0_5 gnd C_bl
Cbb_0_5 bitb_0_5 gnd C_bl
Rb_0_6 bit_0_6 bit_0_7 R_bl
Rbb_0_6 bitb_0_6 bitb_0_7 R_bl
Cb_0_6 bit_0_6 gnd C_bl
Cbb_0_6 bitb_0_6 gnd C_bl
Rb_0_7 bit_0_7 bit_0_8 R_bl
Rbb_0_7 bitb_0_7 bitb_0_8 R_bl
Cb_0_7 bit_0_7 gnd C_bl
Cbb_0_7 bitb_0_7 gnd C_bl
Rb_0_8 bit_0_8 bit_0_9 R_bl
Rbb_0_8 bitb_0_8 bitb_0_9 R_bl
Cb_0_8 bit_0_8 gnd C_bl
Cbb_0_8 bitb_0_8 gnd C_bl
Rb_0_9 bit_0_9 bit_0_10 R_bl
Rbb_0_9 bitb_0_9 bitb_0_10 R_bl
Cb_0_9 bit_0_9 gnd C_bl
Cbb_0_9 bitb_0_9 gnd C_bl
Rb_0_10 bit_0_10 bit_0_11 R_bl
Rbb_0_10 bitb_0_10 bitb_0_11 R_bl
Cb_0_10 bit_0_10 gnd C_bl
Cbb_0_10 bitb_0_10 gnd C_bl
Rb_0_11 bit_0_11 bit_0_12 R_bl
Rbb_0_11 bitb_0_11 bitb_0_12 R_bl
Cb_0_11 bit_0_11 gnd C_bl
Cbb_0_11 bitb_0_11 gnd C_bl
Rb_0_12 bit_0_12 bit_0_13 R_bl
Rbb_0_12 bitb_0_12 bitb_0_13 R_bl
Cb_0_12 bit_0_12 gnd C_bl
Cbb_0_12 bitb_0_12 gnd C_bl
Rb_0_13 bit_0_13 bit_0_14 R_bl
Rbb_0_13 bitb_0_13 bitb_0_14 R_bl
Cb_0_13 bit_0_13 gnd C_bl
Cbb_0_13 bitb_0_13 gnd C_bl
Rb_0_14 bit_0_14 bit_0_15 R_bl
Rbb_0_14 bitb_0_14 bitb_0_15 R_bl
Cb_0_14 bit_0_14 gnd C_bl
Cbb_0_14 bitb_0_14 gnd C_bl
Rb_0_15 bit_0_15 bit_0_16 R_bl
Rbb_0_15 bitb_0_15 bitb_0_16 R_bl
Cb_0_15 bit_0_15 gnd C_bl
Cbb_0_15 bitb_0_15 gnd C_bl
Rb_0_16 bit_0_16 bit_0_17 R_bl
Rbb_0_16 bitb_0_16 bitb_0_17 R_bl
Cb_0_16 bit_0_16 gnd C_bl
Cbb_0_16 bitb_0_16 gnd C_bl
Rb_0_17 bit_0_17 bit_0_18 R_bl
Rbb_0_17 bitb_0_17 bitb_0_18 R_bl
Cb_0_17 bit_0_17 gnd C_bl
Cbb_0_17 bitb_0_17 gnd C_bl
Rb_0_18 bit_0_18 bit_0_19 R_bl
Rbb_0_18 bitb_0_18 bitb_0_19 R_bl
Cb_0_18 bit_0_18 gnd C_bl
Cbb_0_18 bitb_0_18 gnd C_bl
Rb_0_19 bit_0_19 bit_0_20 R_bl
Rbb_0_19 bitb_0_19 bitb_0_20 R_bl
Cb_0_19 bit_0_19 gnd C_bl
Cbb_0_19 bitb_0_19 gnd C_bl
Rb_0_20 bit_0_20 bit_0_21 R_bl
Rbb_0_20 bitb_0_20 bitb_0_21 R_bl
Cb_0_20 bit_0_20 gnd C_bl
Cbb_0_20 bitb_0_20 gnd C_bl
Rb_0_21 bit_0_21 bit_0_22 R_bl
Rbb_0_21 bitb_0_21 bitb_0_22 R_bl
Cb_0_21 bit_0_21 gnd C_bl
Cbb_0_21 bitb_0_21 gnd C_bl
Rb_0_22 bit_0_22 bit_0_23 R_bl
Rbb_0_22 bitb_0_22 bitb_0_23 R_bl
Cb_0_22 bit_0_22 gnd C_bl
Cbb_0_22 bitb_0_22 gnd C_bl
Rb_0_23 bit_0_23 bit_0_24 R_bl
Rbb_0_23 bitb_0_23 bitb_0_24 R_bl
Cb_0_23 bit_0_23 gnd C_bl
Cbb_0_23 bitb_0_23 gnd C_bl
Rb_0_24 bit_0_24 bit_0_25 R_bl
Rbb_0_24 bitb_0_24 bitb_0_25 R_bl
Cb_0_24 bit_0_24 gnd C_bl
Cbb_0_24 bitb_0_24 gnd C_bl
Rb_0_25 bit_0_25 bit_0_26 R_bl
Rbb_0_25 bitb_0_25 bitb_0_26 R_bl
Cb_0_25 bit_0_25 gnd C_bl
Cbb_0_25 bitb_0_25 gnd C_bl
Rb_0_26 bit_0_26 bit_0_27 R_bl
Rbb_0_26 bitb_0_26 bitb_0_27 R_bl
Cb_0_26 bit_0_26 gnd C_bl
Cbb_0_26 bitb_0_26 gnd C_bl
Rb_0_27 bit_0_27 bit_0_28 R_bl
Rbb_0_27 bitb_0_27 bitb_0_28 R_bl
Cb_0_27 bit_0_27 gnd C_bl
Cbb_0_27 bitb_0_27 gnd C_bl
Rb_0_28 bit_0_28 bit_0_29 R_bl
Rbb_0_28 bitb_0_28 bitb_0_29 R_bl
Cb_0_28 bit_0_28 gnd C_bl
Cbb_0_28 bitb_0_28 gnd C_bl
Rb_0_29 bit_0_29 bit_0_30 R_bl
Rbb_0_29 bitb_0_29 bitb_0_30 R_bl
Cb_0_29 bit_0_29 gnd C_bl
Cbb_0_29 bitb_0_29 gnd C_bl
Rb_0_30 bit_0_30 bit_0_31 R_bl
Rbb_0_30 bitb_0_30 bitb_0_31 R_bl
Cb_0_30 bit_0_30 gnd C_bl
Cbb_0_30 bitb_0_30 gnd C_bl
Rb_0_31 bit_0_31 bit_0_32 R_bl
Rbb_0_31 bitb_0_31 bitb_0_32 R_bl
Cb_0_31 bit_0_31 gnd C_bl
Cbb_0_31 bitb_0_31 gnd C_bl
Rb_0_32 bit_0_32 bit_0_33 R_bl
Rbb_0_32 bitb_0_32 bitb_0_33 R_bl
Cb_0_32 bit_0_32 gnd C_bl
Cbb_0_32 bitb_0_32 gnd C_bl
Rb_0_33 bit_0_33 bit_0_34 R_bl
Rbb_0_33 bitb_0_33 bitb_0_34 R_bl
Cb_0_33 bit_0_33 gnd C_bl
Cbb_0_33 bitb_0_33 gnd C_bl
Rb_0_34 bit_0_34 bit_0_35 R_bl
Rbb_0_34 bitb_0_34 bitb_0_35 R_bl
Cb_0_34 bit_0_34 gnd C_bl
Cbb_0_34 bitb_0_34 gnd C_bl
Rb_0_35 bit_0_35 bit_0_36 R_bl
Rbb_0_35 bitb_0_35 bitb_0_36 R_bl
Cb_0_35 bit_0_35 gnd C_bl
Cbb_0_35 bitb_0_35 gnd C_bl
Rb_0_36 bit_0_36 bit_0_37 R_bl
Rbb_0_36 bitb_0_36 bitb_0_37 R_bl
Cb_0_36 bit_0_36 gnd C_bl
Cbb_0_36 bitb_0_36 gnd C_bl
Rb_0_37 bit_0_37 bit_0_38 R_bl
Rbb_0_37 bitb_0_37 bitb_0_38 R_bl
Cb_0_37 bit_0_37 gnd C_bl
Cbb_0_37 bitb_0_37 gnd C_bl
Rb_0_38 bit_0_38 bit_0_39 R_bl
Rbb_0_38 bitb_0_38 bitb_0_39 R_bl
Cb_0_38 bit_0_38 gnd C_bl
Cbb_0_38 bitb_0_38 gnd C_bl
Rb_0_39 bit_0_39 bit_0_40 R_bl
Rbb_0_39 bitb_0_39 bitb_0_40 R_bl
Cb_0_39 bit_0_39 gnd C_bl
Cbb_0_39 bitb_0_39 gnd C_bl
Rb_0_40 bit_0_40 bit_0_41 R_bl
Rbb_0_40 bitb_0_40 bitb_0_41 R_bl
Cb_0_40 bit_0_40 gnd C_bl
Cbb_0_40 bitb_0_40 gnd C_bl
Rb_0_41 bit_0_41 bit_0_42 R_bl
Rbb_0_41 bitb_0_41 bitb_0_42 R_bl
Cb_0_41 bit_0_41 gnd C_bl
Cbb_0_41 bitb_0_41 gnd C_bl
Rb_0_42 bit_0_42 bit_0_43 R_bl
Rbb_0_42 bitb_0_42 bitb_0_43 R_bl
Cb_0_42 bit_0_42 gnd C_bl
Cbb_0_42 bitb_0_42 gnd C_bl
Rb_0_43 bit_0_43 bit_0_44 R_bl
Rbb_0_43 bitb_0_43 bitb_0_44 R_bl
Cb_0_43 bit_0_43 gnd C_bl
Cbb_0_43 bitb_0_43 gnd C_bl
Rb_0_44 bit_0_44 bit_0_45 R_bl
Rbb_0_44 bitb_0_44 bitb_0_45 R_bl
Cb_0_44 bit_0_44 gnd C_bl
Cbb_0_44 bitb_0_44 gnd C_bl
Rb_0_45 bit_0_45 bit_0_46 R_bl
Rbb_0_45 bitb_0_45 bitb_0_46 R_bl
Cb_0_45 bit_0_45 gnd C_bl
Cbb_0_45 bitb_0_45 gnd C_bl
Rb_0_46 bit_0_46 bit_0_47 R_bl
Rbb_0_46 bitb_0_46 bitb_0_47 R_bl
Cb_0_46 bit_0_46 gnd C_bl
Cbb_0_46 bitb_0_46 gnd C_bl
Rb_0_47 bit_0_47 bit_0_48 R_bl
Rbb_0_47 bitb_0_47 bitb_0_48 R_bl
Cb_0_47 bit_0_47 gnd C_bl
Cbb_0_47 bitb_0_47 gnd C_bl
Rb_0_48 bit_0_48 bit_0_49 R_bl
Rbb_0_48 bitb_0_48 bitb_0_49 R_bl
Cb_0_48 bit_0_48 gnd C_bl
Cbb_0_48 bitb_0_48 gnd C_bl
Rb_0_49 bit_0_49 bit_0_50 R_bl
Rbb_0_49 bitb_0_49 bitb_0_50 R_bl
Cb_0_49 bit_0_49 gnd C_bl
Cbb_0_49 bitb_0_49 gnd C_bl
Rb_0_50 bit_0_50 bit_0_51 R_bl
Rbb_0_50 bitb_0_50 bitb_0_51 R_bl
Cb_0_50 bit_0_50 gnd C_bl
Cbb_0_50 bitb_0_50 gnd C_bl
Rb_0_51 bit_0_51 bit_0_52 R_bl
Rbb_0_51 bitb_0_51 bitb_0_52 R_bl
Cb_0_51 bit_0_51 gnd C_bl
Cbb_0_51 bitb_0_51 gnd C_bl
Rb_0_52 bit_0_52 bit_0_53 R_bl
Rbb_0_52 bitb_0_52 bitb_0_53 R_bl
Cb_0_52 bit_0_52 gnd C_bl
Cbb_0_52 bitb_0_52 gnd C_bl
Rb_0_53 bit_0_53 bit_0_54 R_bl
Rbb_0_53 bitb_0_53 bitb_0_54 R_bl
Cb_0_53 bit_0_53 gnd C_bl
Cbb_0_53 bitb_0_53 gnd C_bl
Rb_0_54 bit_0_54 bit_0_55 R_bl
Rbb_0_54 bitb_0_54 bitb_0_55 R_bl
Cb_0_54 bit_0_54 gnd C_bl
Cbb_0_54 bitb_0_54 gnd C_bl
Rb_0_55 bit_0_55 bit_0_56 R_bl
Rbb_0_55 bitb_0_55 bitb_0_56 R_bl
Cb_0_55 bit_0_55 gnd C_bl
Cbb_0_55 bitb_0_55 gnd C_bl
Rb_0_56 bit_0_56 bit_0_57 R_bl
Rbb_0_56 bitb_0_56 bitb_0_57 R_bl
Cb_0_56 bit_0_56 gnd C_bl
Cbb_0_56 bitb_0_56 gnd C_bl
Rb_0_57 bit_0_57 bit_0_58 R_bl
Rbb_0_57 bitb_0_57 bitb_0_58 R_bl
Cb_0_57 bit_0_57 gnd C_bl
Cbb_0_57 bitb_0_57 gnd C_bl
Rb_0_58 bit_0_58 bit_0_59 R_bl
Rbb_0_58 bitb_0_58 bitb_0_59 R_bl
Cb_0_58 bit_0_58 gnd C_bl
Cbb_0_58 bitb_0_58 gnd C_bl
Rb_0_59 bit_0_59 bit_0_60 R_bl
Rbb_0_59 bitb_0_59 bitb_0_60 R_bl
Cb_0_59 bit_0_59 gnd C_bl
Cbb_0_59 bitb_0_59 gnd C_bl
Rb_0_60 bit_0_60 bit_0_61 R_bl
Rbb_0_60 bitb_0_60 bitb_0_61 R_bl
Cb_0_60 bit_0_60 gnd C_bl
Cbb_0_60 bitb_0_60 gnd C_bl
Rb_0_61 bit_0_61 bit_0_62 R_bl
Rbb_0_61 bitb_0_61 bitb_0_62 R_bl
Cb_0_61 bit_0_61 gnd C_bl
Cbb_0_61 bitb_0_61 gnd C_bl
Rb_0_62 bit_0_62 bit_0_63 R_bl
Rbb_0_62 bitb_0_62 bitb_0_63 R_bl
Cb_0_62 bit_0_62 gnd C_bl
Cbb_0_62 bitb_0_62 gnd C_bl
Rb_0_63 bit_0_63 bit_0_64 R_bl
Rbb_0_63 bitb_0_63 bitb_0_64 R_bl
Cb_0_63 bit_0_63 gnd C_bl
Cbb_0_63 bitb_0_63 gnd C_bl
Rb_0_64 bit_0_64 bit_0_65 R_bl
Rbb_0_64 bitb_0_64 bitb_0_65 R_bl
Cb_0_64 bit_0_64 gnd C_bl
Cbb_0_64 bitb_0_64 gnd C_bl
Rb_0_65 bit_0_65 bit_0_66 R_bl
Rbb_0_65 bitb_0_65 bitb_0_66 R_bl
Cb_0_65 bit_0_65 gnd C_bl
Cbb_0_65 bitb_0_65 gnd C_bl
Rb_0_66 bit_0_66 bit_0_67 R_bl
Rbb_0_66 bitb_0_66 bitb_0_67 R_bl
Cb_0_66 bit_0_66 gnd C_bl
Cbb_0_66 bitb_0_66 gnd C_bl
Rb_0_67 bit_0_67 bit_0_68 R_bl
Rbb_0_67 bitb_0_67 bitb_0_68 R_bl
Cb_0_67 bit_0_67 gnd C_bl
Cbb_0_67 bitb_0_67 gnd C_bl
Rb_0_68 bit_0_68 bit_0_69 R_bl
Rbb_0_68 bitb_0_68 bitb_0_69 R_bl
Cb_0_68 bit_0_68 gnd C_bl
Cbb_0_68 bitb_0_68 gnd C_bl
Rb_0_69 bit_0_69 bit_0_70 R_bl
Rbb_0_69 bitb_0_69 bitb_0_70 R_bl
Cb_0_69 bit_0_69 gnd C_bl
Cbb_0_69 bitb_0_69 gnd C_bl
Rb_0_70 bit_0_70 bit_0_71 R_bl
Rbb_0_70 bitb_0_70 bitb_0_71 R_bl
Cb_0_70 bit_0_70 gnd C_bl
Cbb_0_70 bitb_0_70 gnd C_bl
Rb_0_71 bit_0_71 bit_0_72 R_bl
Rbb_0_71 bitb_0_71 bitb_0_72 R_bl
Cb_0_71 bit_0_71 gnd C_bl
Cbb_0_71 bitb_0_71 gnd C_bl
Rb_0_72 bit_0_72 bit_0_73 R_bl
Rbb_0_72 bitb_0_72 bitb_0_73 R_bl
Cb_0_72 bit_0_72 gnd C_bl
Cbb_0_72 bitb_0_72 gnd C_bl
Rb_0_73 bit_0_73 bit_0_74 R_bl
Rbb_0_73 bitb_0_73 bitb_0_74 R_bl
Cb_0_73 bit_0_73 gnd C_bl
Cbb_0_73 bitb_0_73 gnd C_bl
Rb_0_74 bit_0_74 bit_0_75 R_bl
Rbb_0_74 bitb_0_74 bitb_0_75 R_bl
Cb_0_74 bit_0_74 gnd C_bl
Cbb_0_74 bitb_0_74 gnd C_bl
Rb_0_75 bit_0_75 bit_0_76 R_bl
Rbb_0_75 bitb_0_75 bitb_0_76 R_bl
Cb_0_75 bit_0_75 gnd C_bl
Cbb_0_75 bitb_0_75 gnd C_bl
Rb_0_76 bit_0_76 bit_0_77 R_bl
Rbb_0_76 bitb_0_76 bitb_0_77 R_bl
Cb_0_76 bit_0_76 gnd C_bl
Cbb_0_76 bitb_0_76 gnd C_bl
Rb_0_77 bit_0_77 bit_0_78 R_bl
Rbb_0_77 bitb_0_77 bitb_0_78 R_bl
Cb_0_77 bit_0_77 gnd C_bl
Cbb_0_77 bitb_0_77 gnd C_bl
Rb_0_78 bit_0_78 bit_0_79 R_bl
Rbb_0_78 bitb_0_78 bitb_0_79 R_bl
Cb_0_78 bit_0_78 gnd C_bl
Cbb_0_78 bitb_0_78 gnd C_bl
Rb_0_79 bit_0_79 bit_0_80 R_bl
Rbb_0_79 bitb_0_79 bitb_0_80 R_bl
Cb_0_79 bit_0_79 gnd C_bl
Cbb_0_79 bitb_0_79 gnd C_bl
Rb_0_80 bit_0_80 bit_0_81 R_bl
Rbb_0_80 bitb_0_80 bitb_0_81 R_bl
Cb_0_80 bit_0_80 gnd C_bl
Cbb_0_80 bitb_0_80 gnd C_bl
Rb_0_81 bit_0_81 bit_0_82 R_bl
Rbb_0_81 bitb_0_81 bitb_0_82 R_bl
Cb_0_81 bit_0_81 gnd C_bl
Cbb_0_81 bitb_0_81 gnd C_bl
Rb_0_82 bit_0_82 bit_0_83 R_bl
Rbb_0_82 bitb_0_82 bitb_0_83 R_bl
Cb_0_82 bit_0_82 gnd C_bl
Cbb_0_82 bitb_0_82 gnd C_bl
Rb_0_83 bit_0_83 bit_0_84 R_bl
Rbb_0_83 bitb_0_83 bitb_0_84 R_bl
Cb_0_83 bit_0_83 gnd C_bl
Cbb_0_83 bitb_0_83 gnd C_bl
Rb_0_84 bit_0_84 bit_0_85 R_bl
Rbb_0_84 bitb_0_84 bitb_0_85 R_bl
Cb_0_84 bit_0_84 gnd C_bl
Cbb_0_84 bitb_0_84 gnd C_bl
Rb_0_85 bit_0_85 bit_0_86 R_bl
Rbb_0_85 bitb_0_85 bitb_0_86 R_bl
Cb_0_85 bit_0_85 gnd C_bl
Cbb_0_85 bitb_0_85 gnd C_bl
Rb_0_86 bit_0_86 bit_0_87 R_bl
Rbb_0_86 bitb_0_86 bitb_0_87 R_bl
Cb_0_86 bit_0_86 gnd C_bl
Cbb_0_86 bitb_0_86 gnd C_bl
Rb_0_87 bit_0_87 bit_0_88 R_bl
Rbb_0_87 bitb_0_87 bitb_0_88 R_bl
Cb_0_87 bit_0_87 gnd C_bl
Cbb_0_87 bitb_0_87 gnd C_bl
Rb_0_88 bit_0_88 bit_0_89 R_bl
Rbb_0_88 bitb_0_88 bitb_0_89 R_bl
Cb_0_88 bit_0_88 gnd C_bl
Cbb_0_88 bitb_0_88 gnd C_bl
Rb_0_89 bit_0_89 bit_0_90 R_bl
Rbb_0_89 bitb_0_89 bitb_0_90 R_bl
Cb_0_89 bit_0_89 gnd C_bl
Cbb_0_89 bitb_0_89 gnd C_bl
Rb_0_90 bit_0_90 bit_0_91 R_bl
Rbb_0_90 bitb_0_90 bitb_0_91 R_bl
Cb_0_90 bit_0_90 gnd C_bl
Cbb_0_90 bitb_0_90 gnd C_bl
Rb_0_91 bit_0_91 bit_0_92 R_bl
Rbb_0_91 bitb_0_91 bitb_0_92 R_bl
Cb_0_91 bit_0_91 gnd C_bl
Cbb_0_91 bitb_0_91 gnd C_bl
Rb_0_92 bit_0_92 bit_0_93 R_bl
Rbb_0_92 bitb_0_92 bitb_0_93 R_bl
Cb_0_92 bit_0_92 gnd C_bl
Cbb_0_92 bitb_0_92 gnd C_bl
Rb_0_93 bit_0_93 bit_0_94 R_bl
Rbb_0_93 bitb_0_93 bitb_0_94 R_bl
Cb_0_93 bit_0_93 gnd C_bl
Cbb_0_93 bitb_0_93 gnd C_bl
Rb_0_94 bit_0_94 bit_0_95 R_bl
Rbb_0_94 bitb_0_94 bitb_0_95 R_bl
Cb_0_94 bit_0_94 gnd C_bl
Cbb_0_94 bitb_0_94 gnd C_bl
Rb_0_95 bit_0_95 bit_0_96 R_bl
Rbb_0_95 bitb_0_95 bitb_0_96 R_bl
Cb_0_95 bit_0_95 gnd C_bl
Cbb_0_95 bitb_0_95 gnd C_bl
Rb_0_96 bit_0_96 bit_0_97 R_bl
Rbb_0_96 bitb_0_96 bitb_0_97 R_bl
Cb_0_96 bit_0_96 gnd C_bl
Cbb_0_96 bitb_0_96 gnd C_bl
Rb_0_97 bit_0_97 bit_0_98 R_bl
Rbb_0_97 bitb_0_97 bitb_0_98 R_bl
Cb_0_97 bit_0_97 gnd C_bl
Cbb_0_97 bitb_0_97 gnd C_bl
Rb_0_98 bit_0_98 bit_0_99 R_bl
Rbb_0_98 bitb_0_98 bitb_0_99 R_bl
Cb_0_98 bit_0_98 gnd C_bl
Cbb_0_98 bitb_0_98 gnd C_bl
Rb_0_99 bit_0_99 bit_0_100 R_bl
Rbb_0_99 bitb_0_99 bitb_0_100 R_bl
Cb_0_99 bit_0_99 gnd C_bl
Cbb_0_99 bitb_0_99 gnd C_bl
Rb_1_0 bit_1_0 bit_1_1 R_bl
Rbb_1_0 bitb_1_0 bitb_1_1 R_bl
Cb_1_0 bit_1_0 gnd C_bl
Cbb_1_0 bitb_1_0 gnd C_bl
Rb_1_1 bit_1_1 bit_1_2 R_bl
Rbb_1_1 bitb_1_1 bitb_1_2 R_bl
Cb_1_1 bit_1_1 gnd C_bl
Cbb_1_1 bitb_1_1 gnd C_bl
Rb_1_2 bit_1_2 bit_1_3 R_bl
Rbb_1_2 bitb_1_2 bitb_1_3 R_bl
Cb_1_2 bit_1_2 gnd C_bl
Cbb_1_2 bitb_1_2 gnd C_bl
Rb_1_3 bit_1_3 bit_1_4 R_bl
Rbb_1_3 bitb_1_3 bitb_1_4 R_bl
Cb_1_3 bit_1_3 gnd C_bl
Cbb_1_3 bitb_1_3 gnd C_bl
Rb_1_4 bit_1_4 bit_1_5 R_bl
Rbb_1_4 bitb_1_4 bitb_1_5 R_bl
Cb_1_4 bit_1_4 gnd C_bl
Cbb_1_4 bitb_1_4 gnd C_bl
Rb_1_5 bit_1_5 bit_1_6 R_bl
Rbb_1_5 bitb_1_5 bitb_1_6 R_bl
Cb_1_5 bit_1_5 gnd C_bl
Cbb_1_5 bitb_1_5 gnd C_bl
Rb_1_6 bit_1_6 bit_1_7 R_bl
Rbb_1_6 bitb_1_6 bitb_1_7 R_bl
Cb_1_6 bit_1_6 gnd C_bl
Cbb_1_6 bitb_1_6 gnd C_bl
Rb_1_7 bit_1_7 bit_1_8 R_bl
Rbb_1_7 bitb_1_7 bitb_1_8 R_bl
Cb_1_7 bit_1_7 gnd C_bl
Cbb_1_7 bitb_1_7 gnd C_bl
Rb_1_8 bit_1_8 bit_1_9 R_bl
Rbb_1_8 bitb_1_8 bitb_1_9 R_bl
Cb_1_8 bit_1_8 gnd C_bl
Cbb_1_8 bitb_1_8 gnd C_bl
Rb_1_9 bit_1_9 bit_1_10 R_bl
Rbb_1_9 bitb_1_9 bitb_1_10 R_bl
Cb_1_9 bit_1_9 gnd C_bl
Cbb_1_9 bitb_1_9 gnd C_bl
Rb_1_10 bit_1_10 bit_1_11 R_bl
Rbb_1_10 bitb_1_10 bitb_1_11 R_bl
Cb_1_10 bit_1_10 gnd C_bl
Cbb_1_10 bitb_1_10 gnd C_bl
Rb_1_11 bit_1_11 bit_1_12 R_bl
Rbb_1_11 bitb_1_11 bitb_1_12 R_bl
Cb_1_11 bit_1_11 gnd C_bl
Cbb_1_11 bitb_1_11 gnd C_bl
Rb_1_12 bit_1_12 bit_1_13 R_bl
Rbb_1_12 bitb_1_12 bitb_1_13 R_bl
Cb_1_12 bit_1_12 gnd C_bl
Cbb_1_12 bitb_1_12 gnd C_bl
Rb_1_13 bit_1_13 bit_1_14 R_bl
Rbb_1_13 bitb_1_13 bitb_1_14 R_bl
Cb_1_13 bit_1_13 gnd C_bl
Cbb_1_13 bitb_1_13 gnd C_bl
Rb_1_14 bit_1_14 bit_1_15 R_bl
Rbb_1_14 bitb_1_14 bitb_1_15 R_bl
Cb_1_14 bit_1_14 gnd C_bl
Cbb_1_14 bitb_1_14 gnd C_bl
Rb_1_15 bit_1_15 bit_1_16 R_bl
Rbb_1_15 bitb_1_15 bitb_1_16 R_bl
Cb_1_15 bit_1_15 gnd C_bl
Cbb_1_15 bitb_1_15 gnd C_bl
Rb_1_16 bit_1_16 bit_1_17 R_bl
Rbb_1_16 bitb_1_16 bitb_1_17 R_bl
Cb_1_16 bit_1_16 gnd C_bl
Cbb_1_16 bitb_1_16 gnd C_bl
Rb_1_17 bit_1_17 bit_1_18 R_bl
Rbb_1_17 bitb_1_17 bitb_1_18 R_bl
Cb_1_17 bit_1_17 gnd C_bl
Cbb_1_17 bitb_1_17 gnd C_bl
Rb_1_18 bit_1_18 bit_1_19 R_bl
Rbb_1_18 bitb_1_18 bitb_1_19 R_bl
Cb_1_18 bit_1_18 gnd C_bl
Cbb_1_18 bitb_1_18 gnd C_bl
Rb_1_19 bit_1_19 bit_1_20 R_bl
Rbb_1_19 bitb_1_19 bitb_1_20 R_bl
Cb_1_19 bit_1_19 gnd C_bl
Cbb_1_19 bitb_1_19 gnd C_bl
Rb_1_20 bit_1_20 bit_1_21 R_bl
Rbb_1_20 bitb_1_20 bitb_1_21 R_bl
Cb_1_20 bit_1_20 gnd C_bl
Cbb_1_20 bitb_1_20 gnd C_bl
Rb_1_21 bit_1_21 bit_1_22 R_bl
Rbb_1_21 bitb_1_21 bitb_1_22 R_bl
Cb_1_21 bit_1_21 gnd C_bl
Cbb_1_21 bitb_1_21 gnd C_bl
Rb_1_22 bit_1_22 bit_1_23 R_bl
Rbb_1_22 bitb_1_22 bitb_1_23 R_bl
Cb_1_22 bit_1_22 gnd C_bl
Cbb_1_22 bitb_1_22 gnd C_bl
Rb_1_23 bit_1_23 bit_1_24 R_bl
Rbb_1_23 bitb_1_23 bitb_1_24 R_bl
Cb_1_23 bit_1_23 gnd C_bl
Cbb_1_23 bitb_1_23 gnd C_bl
Rb_1_24 bit_1_24 bit_1_25 R_bl
Rbb_1_24 bitb_1_24 bitb_1_25 R_bl
Cb_1_24 bit_1_24 gnd C_bl
Cbb_1_24 bitb_1_24 gnd C_bl
Rb_1_25 bit_1_25 bit_1_26 R_bl
Rbb_1_25 bitb_1_25 bitb_1_26 R_bl
Cb_1_25 bit_1_25 gnd C_bl
Cbb_1_25 bitb_1_25 gnd C_bl
Rb_1_26 bit_1_26 bit_1_27 R_bl
Rbb_1_26 bitb_1_26 bitb_1_27 R_bl
Cb_1_26 bit_1_26 gnd C_bl
Cbb_1_26 bitb_1_26 gnd C_bl
Rb_1_27 bit_1_27 bit_1_28 R_bl
Rbb_1_27 bitb_1_27 bitb_1_28 R_bl
Cb_1_27 bit_1_27 gnd C_bl
Cbb_1_27 bitb_1_27 gnd C_bl
Rb_1_28 bit_1_28 bit_1_29 R_bl
Rbb_1_28 bitb_1_28 bitb_1_29 R_bl
Cb_1_28 bit_1_28 gnd C_bl
Cbb_1_28 bitb_1_28 gnd C_bl
Rb_1_29 bit_1_29 bit_1_30 R_bl
Rbb_1_29 bitb_1_29 bitb_1_30 R_bl
Cb_1_29 bit_1_29 gnd C_bl
Cbb_1_29 bitb_1_29 gnd C_bl
Rb_1_30 bit_1_30 bit_1_31 R_bl
Rbb_1_30 bitb_1_30 bitb_1_31 R_bl
Cb_1_30 bit_1_30 gnd C_bl
Cbb_1_30 bitb_1_30 gnd C_bl
Rb_1_31 bit_1_31 bit_1_32 R_bl
Rbb_1_31 bitb_1_31 bitb_1_32 R_bl
Cb_1_31 bit_1_31 gnd C_bl
Cbb_1_31 bitb_1_31 gnd C_bl
Rb_1_32 bit_1_32 bit_1_33 R_bl
Rbb_1_32 bitb_1_32 bitb_1_33 R_bl
Cb_1_32 bit_1_32 gnd C_bl
Cbb_1_32 bitb_1_32 gnd C_bl
Rb_1_33 bit_1_33 bit_1_34 R_bl
Rbb_1_33 bitb_1_33 bitb_1_34 R_bl
Cb_1_33 bit_1_33 gnd C_bl
Cbb_1_33 bitb_1_33 gnd C_bl
Rb_1_34 bit_1_34 bit_1_35 R_bl
Rbb_1_34 bitb_1_34 bitb_1_35 R_bl
Cb_1_34 bit_1_34 gnd C_bl
Cbb_1_34 bitb_1_34 gnd C_bl
Rb_1_35 bit_1_35 bit_1_36 R_bl
Rbb_1_35 bitb_1_35 bitb_1_36 R_bl
Cb_1_35 bit_1_35 gnd C_bl
Cbb_1_35 bitb_1_35 gnd C_bl
Rb_1_36 bit_1_36 bit_1_37 R_bl
Rbb_1_36 bitb_1_36 bitb_1_37 R_bl
Cb_1_36 bit_1_36 gnd C_bl
Cbb_1_36 bitb_1_36 gnd C_bl
Rb_1_37 bit_1_37 bit_1_38 R_bl
Rbb_1_37 bitb_1_37 bitb_1_38 R_bl
Cb_1_37 bit_1_37 gnd C_bl
Cbb_1_37 bitb_1_37 gnd C_bl
Rb_1_38 bit_1_38 bit_1_39 R_bl
Rbb_1_38 bitb_1_38 bitb_1_39 R_bl
Cb_1_38 bit_1_38 gnd C_bl
Cbb_1_38 bitb_1_38 gnd C_bl
Rb_1_39 bit_1_39 bit_1_40 R_bl
Rbb_1_39 bitb_1_39 bitb_1_40 R_bl
Cb_1_39 bit_1_39 gnd C_bl
Cbb_1_39 bitb_1_39 gnd C_bl
Rb_1_40 bit_1_40 bit_1_41 R_bl
Rbb_1_40 bitb_1_40 bitb_1_41 R_bl
Cb_1_40 bit_1_40 gnd C_bl
Cbb_1_40 bitb_1_40 gnd C_bl
Rb_1_41 bit_1_41 bit_1_42 R_bl
Rbb_1_41 bitb_1_41 bitb_1_42 R_bl
Cb_1_41 bit_1_41 gnd C_bl
Cbb_1_41 bitb_1_41 gnd C_bl
Rb_1_42 bit_1_42 bit_1_43 R_bl
Rbb_1_42 bitb_1_42 bitb_1_43 R_bl
Cb_1_42 bit_1_42 gnd C_bl
Cbb_1_42 bitb_1_42 gnd C_bl
Rb_1_43 bit_1_43 bit_1_44 R_bl
Rbb_1_43 bitb_1_43 bitb_1_44 R_bl
Cb_1_43 bit_1_43 gnd C_bl
Cbb_1_43 bitb_1_43 gnd C_bl
Rb_1_44 bit_1_44 bit_1_45 R_bl
Rbb_1_44 bitb_1_44 bitb_1_45 R_bl
Cb_1_44 bit_1_44 gnd C_bl
Cbb_1_44 bitb_1_44 gnd C_bl
Rb_1_45 bit_1_45 bit_1_46 R_bl
Rbb_1_45 bitb_1_45 bitb_1_46 R_bl
Cb_1_45 bit_1_45 gnd C_bl
Cbb_1_45 bitb_1_45 gnd C_bl
Rb_1_46 bit_1_46 bit_1_47 R_bl
Rbb_1_46 bitb_1_46 bitb_1_47 R_bl
Cb_1_46 bit_1_46 gnd C_bl
Cbb_1_46 bitb_1_46 gnd C_bl
Rb_1_47 bit_1_47 bit_1_48 R_bl
Rbb_1_47 bitb_1_47 bitb_1_48 R_bl
Cb_1_47 bit_1_47 gnd C_bl
Cbb_1_47 bitb_1_47 gnd C_bl
Rb_1_48 bit_1_48 bit_1_49 R_bl
Rbb_1_48 bitb_1_48 bitb_1_49 R_bl
Cb_1_48 bit_1_48 gnd C_bl
Cbb_1_48 bitb_1_48 gnd C_bl
Rb_1_49 bit_1_49 bit_1_50 R_bl
Rbb_1_49 bitb_1_49 bitb_1_50 R_bl
Cb_1_49 bit_1_49 gnd C_bl
Cbb_1_49 bitb_1_49 gnd C_bl
Rb_1_50 bit_1_50 bit_1_51 R_bl
Rbb_1_50 bitb_1_50 bitb_1_51 R_bl
Cb_1_50 bit_1_50 gnd C_bl
Cbb_1_50 bitb_1_50 gnd C_bl
Rb_1_51 bit_1_51 bit_1_52 R_bl
Rbb_1_51 bitb_1_51 bitb_1_52 R_bl
Cb_1_51 bit_1_51 gnd C_bl
Cbb_1_51 bitb_1_51 gnd C_bl
Rb_1_52 bit_1_52 bit_1_53 R_bl
Rbb_1_52 bitb_1_52 bitb_1_53 R_bl
Cb_1_52 bit_1_52 gnd C_bl
Cbb_1_52 bitb_1_52 gnd C_bl
Rb_1_53 bit_1_53 bit_1_54 R_bl
Rbb_1_53 bitb_1_53 bitb_1_54 R_bl
Cb_1_53 bit_1_53 gnd C_bl
Cbb_1_53 bitb_1_53 gnd C_bl
Rb_1_54 bit_1_54 bit_1_55 R_bl
Rbb_1_54 bitb_1_54 bitb_1_55 R_bl
Cb_1_54 bit_1_54 gnd C_bl
Cbb_1_54 bitb_1_54 gnd C_bl
Rb_1_55 bit_1_55 bit_1_56 R_bl
Rbb_1_55 bitb_1_55 bitb_1_56 R_bl
Cb_1_55 bit_1_55 gnd C_bl
Cbb_1_55 bitb_1_55 gnd C_bl
Rb_1_56 bit_1_56 bit_1_57 R_bl
Rbb_1_56 bitb_1_56 bitb_1_57 R_bl
Cb_1_56 bit_1_56 gnd C_bl
Cbb_1_56 bitb_1_56 gnd C_bl
Rb_1_57 bit_1_57 bit_1_58 R_bl
Rbb_1_57 bitb_1_57 bitb_1_58 R_bl
Cb_1_57 bit_1_57 gnd C_bl
Cbb_1_57 bitb_1_57 gnd C_bl
Rb_1_58 bit_1_58 bit_1_59 R_bl
Rbb_1_58 bitb_1_58 bitb_1_59 R_bl
Cb_1_58 bit_1_58 gnd C_bl
Cbb_1_58 bitb_1_58 gnd C_bl
Rb_1_59 bit_1_59 bit_1_60 R_bl
Rbb_1_59 bitb_1_59 bitb_1_60 R_bl
Cb_1_59 bit_1_59 gnd C_bl
Cbb_1_59 bitb_1_59 gnd C_bl
Rb_1_60 bit_1_60 bit_1_61 R_bl
Rbb_1_60 bitb_1_60 bitb_1_61 R_bl
Cb_1_60 bit_1_60 gnd C_bl
Cbb_1_60 bitb_1_60 gnd C_bl
Rb_1_61 bit_1_61 bit_1_62 R_bl
Rbb_1_61 bitb_1_61 bitb_1_62 R_bl
Cb_1_61 bit_1_61 gnd C_bl
Cbb_1_61 bitb_1_61 gnd C_bl
Rb_1_62 bit_1_62 bit_1_63 R_bl
Rbb_1_62 bitb_1_62 bitb_1_63 R_bl
Cb_1_62 bit_1_62 gnd C_bl
Cbb_1_62 bitb_1_62 gnd C_bl
Rb_1_63 bit_1_63 bit_1_64 R_bl
Rbb_1_63 bitb_1_63 bitb_1_64 R_bl
Cb_1_63 bit_1_63 gnd C_bl
Cbb_1_63 bitb_1_63 gnd C_bl
Rb_1_64 bit_1_64 bit_1_65 R_bl
Rbb_1_64 bitb_1_64 bitb_1_65 R_bl
Cb_1_64 bit_1_64 gnd C_bl
Cbb_1_64 bitb_1_64 gnd C_bl
Rb_1_65 bit_1_65 bit_1_66 R_bl
Rbb_1_65 bitb_1_65 bitb_1_66 R_bl
Cb_1_65 bit_1_65 gnd C_bl
Cbb_1_65 bitb_1_65 gnd C_bl
Rb_1_66 bit_1_66 bit_1_67 R_bl
Rbb_1_66 bitb_1_66 bitb_1_67 R_bl
Cb_1_66 bit_1_66 gnd C_bl
Cbb_1_66 bitb_1_66 gnd C_bl
Rb_1_67 bit_1_67 bit_1_68 R_bl
Rbb_1_67 bitb_1_67 bitb_1_68 R_bl
Cb_1_67 bit_1_67 gnd C_bl
Cbb_1_67 bitb_1_67 gnd C_bl
Rb_1_68 bit_1_68 bit_1_69 R_bl
Rbb_1_68 bitb_1_68 bitb_1_69 R_bl
Cb_1_68 bit_1_68 gnd C_bl
Cbb_1_68 bitb_1_68 gnd C_bl
Rb_1_69 bit_1_69 bit_1_70 R_bl
Rbb_1_69 bitb_1_69 bitb_1_70 R_bl
Cb_1_69 bit_1_69 gnd C_bl
Cbb_1_69 bitb_1_69 gnd C_bl
Rb_1_70 bit_1_70 bit_1_71 R_bl
Rbb_1_70 bitb_1_70 bitb_1_71 R_bl
Cb_1_70 bit_1_70 gnd C_bl
Cbb_1_70 bitb_1_70 gnd C_bl
Rb_1_71 bit_1_71 bit_1_72 R_bl
Rbb_1_71 bitb_1_71 bitb_1_72 R_bl
Cb_1_71 bit_1_71 gnd C_bl
Cbb_1_71 bitb_1_71 gnd C_bl
Rb_1_72 bit_1_72 bit_1_73 R_bl
Rbb_1_72 bitb_1_72 bitb_1_73 R_bl
Cb_1_72 bit_1_72 gnd C_bl
Cbb_1_72 bitb_1_72 gnd C_bl
Rb_1_73 bit_1_73 bit_1_74 R_bl
Rbb_1_73 bitb_1_73 bitb_1_74 R_bl
Cb_1_73 bit_1_73 gnd C_bl
Cbb_1_73 bitb_1_73 gnd C_bl
Rb_1_74 bit_1_74 bit_1_75 R_bl
Rbb_1_74 bitb_1_74 bitb_1_75 R_bl
Cb_1_74 bit_1_74 gnd C_bl
Cbb_1_74 bitb_1_74 gnd C_bl
Rb_1_75 bit_1_75 bit_1_76 R_bl
Rbb_1_75 bitb_1_75 bitb_1_76 R_bl
Cb_1_75 bit_1_75 gnd C_bl
Cbb_1_75 bitb_1_75 gnd C_bl
Rb_1_76 bit_1_76 bit_1_77 R_bl
Rbb_1_76 bitb_1_76 bitb_1_77 R_bl
Cb_1_76 bit_1_76 gnd C_bl
Cbb_1_76 bitb_1_76 gnd C_bl
Rb_1_77 bit_1_77 bit_1_78 R_bl
Rbb_1_77 bitb_1_77 bitb_1_78 R_bl
Cb_1_77 bit_1_77 gnd C_bl
Cbb_1_77 bitb_1_77 gnd C_bl
Rb_1_78 bit_1_78 bit_1_79 R_bl
Rbb_1_78 bitb_1_78 bitb_1_79 R_bl
Cb_1_78 bit_1_78 gnd C_bl
Cbb_1_78 bitb_1_78 gnd C_bl
Rb_1_79 bit_1_79 bit_1_80 R_bl
Rbb_1_79 bitb_1_79 bitb_1_80 R_bl
Cb_1_79 bit_1_79 gnd C_bl
Cbb_1_79 bitb_1_79 gnd C_bl
Rb_1_80 bit_1_80 bit_1_81 R_bl
Rbb_1_80 bitb_1_80 bitb_1_81 R_bl
Cb_1_80 bit_1_80 gnd C_bl
Cbb_1_80 bitb_1_80 gnd C_bl
Rb_1_81 bit_1_81 bit_1_82 R_bl
Rbb_1_81 bitb_1_81 bitb_1_82 R_bl
Cb_1_81 bit_1_81 gnd C_bl
Cbb_1_81 bitb_1_81 gnd C_bl
Rb_1_82 bit_1_82 bit_1_83 R_bl
Rbb_1_82 bitb_1_82 bitb_1_83 R_bl
Cb_1_82 bit_1_82 gnd C_bl
Cbb_1_82 bitb_1_82 gnd C_bl
Rb_1_83 bit_1_83 bit_1_84 R_bl
Rbb_1_83 bitb_1_83 bitb_1_84 R_bl
Cb_1_83 bit_1_83 gnd C_bl
Cbb_1_83 bitb_1_83 gnd C_bl
Rb_1_84 bit_1_84 bit_1_85 R_bl
Rbb_1_84 bitb_1_84 bitb_1_85 R_bl
Cb_1_84 bit_1_84 gnd C_bl
Cbb_1_84 bitb_1_84 gnd C_bl
Rb_1_85 bit_1_85 bit_1_86 R_bl
Rbb_1_85 bitb_1_85 bitb_1_86 R_bl
Cb_1_85 bit_1_85 gnd C_bl
Cbb_1_85 bitb_1_85 gnd C_bl
Rb_1_86 bit_1_86 bit_1_87 R_bl
Rbb_1_86 bitb_1_86 bitb_1_87 R_bl
Cb_1_86 bit_1_86 gnd C_bl
Cbb_1_86 bitb_1_86 gnd C_bl
Rb_1_87 bit_1_87 bit_1_88 R_bl
Rbb_1_87 bitb_1_87 bitb_1_88 R_bl
Cb_1_87 bit_1_87 gnd C_bl
Cbb_1_87 bitb_1_87 gnd C_bl
Rb_1_88 bit_1_88 bit_1_89 R_bl
Rbb_1_88 bitb_1_88 bitb_1_89 R_bl
Cb_1_88 bit_1_88 gnd C_bl
Cbb_1_88 bitb_1_88 gnd C_bl
Rb_1_89 bit_1_89 bit_1_90 R_bl
Rbb_1_89 bitb_1_89 bitb_1_90 R_bl
Cb_1_89 bit_1_89 gnd C_bl
Cbb_1_89 bitb_1_89 gnd C_bl
Rb_1_90 bit_1_90 bit_1_91 R_bl
Rbb_1_90 bitb_1_90 bitb_1_91 R_bl
Cb_1_90 bit_1_90 gnd C_bl
Cbb_1_90 bitb_1_90 gnd C_bl
Rb_1_91 bit_1_91 bit_1_92 R_bl
Rbb_1_91 bitb_1_91 bitb_1_92 R_bl
Cb_1_91 bit_1_91 gnd C_bl
Cbb_1_91 bitb_1_91 gnd C_bl
Rb_1_92 bit_1_92 bit_1_93 R_bl
Rbb_1_92 bitb_1_92 bitb_1_93 R_bl
Cb_1_92 bit_1_92 gnd C_bl
Cbb_1_92 bitb_1_92 gnd C_bl
Rb_1_93 bit_1_93 bit_1_94 R_bl
Rbb_1_93 bitb_1_93 bitb_1_94 R_bl
Cb_1_93 bit_1_93 gnd C_bl
Cbb_1_93 bitb_1_93 gnd C_bl
Rb_1_94 bit_1_94 bit_1_95 R_bl
Rbb_1_94 bitb_1_94 bitb_1_95 R_bl
Cb_1_94 bit_1_94 gnd C_bl
Cbb_1_94 bitb_1_94 gnd C_bl
Rb_1_95 bit_1_95 bit_1_96 R_bl
Rbb_1_95 bitb_1_95 bitb_1_96 R_bl
Cb_1_95 bit_1_95 gnd C_bl
Cbb_1_95 bitb_1_95 gnd C_bl
Rb_1_96 bit_1_96 bit_1_97 R_bl
Rbb_1_96 bitb_1_96 bitb_1_97 R_bl
Cb_1_96 bit_1_96 gnd C_bl
Cbb_1_96 bitb_1_96 gnd C_bl
Rb_1_97 bit_1_97 bit_1_98 R_bl
Rbb_1_97 bitb_1_97 bitb_1_98 R_bl
Cb_1_97 bit_1_97 gnd C_bl
Cbb_1_97 bitb_1_97 gnd C_bl
Rb_1_98 bit_1_98 bit_1_99 R_bl
Rbb_1_98 bitb_1_98 bitb_1_99 R_bl
Cb_1_98 bit_1_98 gnd C_bl
Cbb_1_98 bitb_1_98 gnd C_bl
Rb_1_99 bit_1_99 bit_1_100 R_bl
Rbb_1_99 bitb_1_99 bitb_1_100 R_bl
Cb_1_99 bit_1_99 gnd C_bl
Cbb_1_99 bitb_1_99 gnd C_bl
Rb_2_0 bit_2_0 bit_2_1 R_bl
Rbb_2_0 bitb_2_0 bitb_2_1 R_bl
Cb_2_0 bit_2_0 gnd C_bl
Cbb_2_0 bitb_2_0 gnd C_bl
Rb_2_1 bit_2_1 bit_2_2 R_bl
Rbb_2_1 bitb_2_1 bitb_2_2 R_bl
Cb_2_1 bit_2_1 gnd C_bl
Cbb_2_1 bitb_2_1 gnd C_bl
Rb_2_2 bit_2_2 bit_2_3 R_bl
Rbb_2_2 bitb_2_2 bitb_2_3 R_bl
Cb_2_2 bit_2_2 gnd C_bl
Cbb_2_2 bitb_2_2 gnd C_bl
Rb_2_3 bit_2_3 bit_2_4 R_bl
Rbb_2_3 bitb_2_3 bitb_2_4 R_bl
Cb_2_3 bit_2_3 gnd C_bl
Cbb_2_3 bitb_2_3 gnd C_bl
Rb_2_4 bit_2_4 bit_2_5 R_bl
Rbb_2_4 bitb_2_4 bitb_2_5 R_bl
Cb_2_4 bit_2_4 gnd C_bl
Cbb_2_4 bitb_2_4 gnd C_bl
Rb_2_5 bit_2_5 bit_2_6 R_bl
Rbb_2_5 bitb_2_5 bitb_2_6 R_bl
Cb_2_5 bit_2_5 gnd C_bl
Cbb_2_5 bitb_2_5 gnd C_bl
Rb_2_6 bit_2_6 bit_2_7 R_bl
Rbb_2_6 bitb_2_6 bitb_2_7 R_bl
Cb_2_6 bit_2_6 gnd C_bl
Cbb_2_6 bitb_2_6 gnd C_bl
Rb_2_7 bit_2_7 bit_2_8 R_bl
Rbb_2_7 bitb_2_7 bitb_2_8 R_bl
Cb_2_7 bit_2_7 gnd C_bl
Cbb_2_7 bitb_2_7 gnd C_bl
Rb_2_8 bit_2_8 bit_2_9 R_bl
Rbb_2_8 bitb_2_8 bitb_2_9 R_bl
Cb_2_8 bit_2_8 gnd C_bl
Cbb_2_8 bitb_2_8 gnd C_bl
Rb_2_9 bit_2_9 bit_2_10 R_bl
Rbb_2_9 bitb_2_9 bitb_2_10 R_bl
Cb_2_9 bit_2_9 gnd C_bl
Cbb_2_9 bitb_2_9 gnd C_bl
Rb_2_10 bit_2_10 bit_2_11 R_bl
Rbb_2_10 bitb_2_10 bitb_2_11 R_bl
Cb_2_10 bit_2_10 gnd C_bl
Cbb_2_10 bitb_2_10 gnd C_bl
Rb_2_11 bit_2_11 bit_2_12 R_bl
Rbb_2_11 bitb_2_11 bitb_2_12 R_bl
Cb_2_11 bit_2_11 gnd C_bl
Cbb_2_11 bitb_2_11 gnd C_bl
Rb_2_12 bit_2_12 bit_2_13 R_bl
Rbb_2_12 bitb_2_12 bitb_2_13 R_bl
Cb_2_12 bit_2_12 gnd C_bl
Cbb_2_12 bitb_2_12 gnd C_bl
Rb_2_13 bit_2_13 bit_2_14 R_bl
Rbb_2_13 bitb_2_13 bitb_2_14 R_bl
Cb_2_13 bit_2_13 gnd C_bl
Cbb_2_13 bitb_2_13 gnd C_bl
Rb_2_14 bit_2_14 bit_2_15 R_bl
Rbb_2_14 bitb_2_14 bitb_2_15 R_bl
Cb_2_14 bit_2_14 gnd C_bl
Cbb_2_14 bitb_2_14 gnd C_bl
Rb_2_15 bit_2_15 bit_2_16 R_bl
Rbb_2_15 bitb_2_15 bitb_2_16 R_bl
Cb_2_15 bit_2_15 gnd C_bl
Cbb_2_15 bitb_2_15 gnd C_bl
Rb_2_16 bit_2_16 bit_2_17 R_bl
Rbb_2_16 bitb_2_16 bitb_2_17 R_bl
Cb_2_16 bit_2_16 gnd C_bl
Cbb_2_16 bitb_2_16 gnd C_bl
Rb_2_17 bit_2_17 bit_2_18 R_bl
Rbb_2_17 bitb_2_17 bitb_2_18 R_bl
Cb_2_17 bit_2_17 gnd C_bl
Cbb_2_17 bitb_2_17 gnd C_bl
Rb_2_18 bit_2_18 bit_2_19 R_bl
Rbb_2_18 bitb_2_18 bitb_2_19 R_bl
Cb_2_18 bit_2_18 gnd C_bl
Cbb_2_18 bitb_2_18 gnd C_bl
Rb_2_19 bit_2_19 bit_2_20 R_bl
Rbb_2_19 bitb_2_19 bitb_2_20 R_bl
Cb_2_19 bit_2_19 gnd C_bl
Cbb_2_19 bitb_2_19 gnd C_bl
Rb_2_20 bit_2_20 bit_2_21 R_bl
Rbb_2_20 bitb_2_20 bitb_2_21 R_bl
Cb_2_20 bit_2_20 gnd C_bl
Cbb_2_20 bitb_2_20 gnd C_bl
Rb_2_21 bit_2_21 bit_2_22 R_bl
Rbb_2_21 bitb_2_21 bitb_2_22 R_bl
Cb_2_21 bit_2_21 gnd C_bl
Cbb_2_21 bitb_2_21 gnd C_bl
Rb_2_22 bit_2_22 bit_2_23 R_bl
Rbb_2_22 bitb_2_22 bitb_2_23 R_bl
Cb_2_22 bit_2_22 gnd C_bl
Cbb_2_22 bitb_2_22 gnd C_bl
Rb_2_23 bit_2_23 bit_2_24 R_bl
Rbb_2_23 bitb_2_23 bitb_2_24 R_bl
Cb_2_23 bit_2_23 gnd C_bl
Cbb_2_23 bitb_2_23 gnd C_bl
Rb_2_24 bit_2_24 bit_2_25 R_bl
Rbb_2_24 bitb_2_24 bitb_2_25 R_bl
Cb_2_24 bit_2_24 gnd C_bl
Cbb_2_24 bitb_2_24 gnd C_bl
Rb_2_25 bit_2_25 bit_2_26 R_bl
Rbb_2_25 bitb_2_25 bitb_2_26 R_bl
Cb_2_25 bit_2_25 gnd C_bl
Cbb_2_25 bitb_2_25 gnd C_bl
Rb_2_26 bit_2_26 bit_2_27 R_bl
Rbb_2_26 bitb_2_26 bitb_2_27 R_bl
Cb_2_26 bit_2_26 gnd C_bl
Cbb_2_26 bitb_2_26 gnd C_bl
Rb_2_27 bit_2_27 bit_2_28 R_bl
Rbb_2_27 bitb_2_27 bitb_2_28 R_bl
Cb_2_27 bit_2_27 gnd C_bl
Cbb_2_27 bitb_2_27 gnd C_bl
Rb_2_28 bit_2_28 bit_2_29 R_bl
Rbb_2_28 bitb_2_28 bitb_2_29 R_bl
Cb_2_28 bit_2_28 gnd C_bl
Cbb_2_28 bitb_2_28 gnd C_bl
Rb_2_29 bit_2_29 bit_2_30 R_bl
Rbb_2_29 bitb_2_29 bitb_2_30 R_bl
Cb_2_29 bit_2_29 gnd C_bl
Cbb_2_29 bitb_2_29 gnd C_bl
Rb_2_30 bit_2_30 bit_2_31 R_bl
Rbb_2_30 bitb_2_30 bitb_2_31 R_bl
Cb_2_30 bit_2_30 gnd C_bl
Cbb_2_30 bitb_2_30 gnd C_bl
Rb_2_31 bit_2_31 bit_2_32 R_bl
Rbb_2_31 bitb_2_31 bitb_2_32 R_bl
Cb_2_31 bit_2_31 gnd C_bl
Cbb_2_31 bitb_2_31 gnd C_bl
Rb_2_32 bit_2_32 bit_2_33 R_bl
Rbb_2_32 bitb_2_32 bitb_2_33 R_bl
Cb_2_32 bit_2_32 gnd C_bl
Cbb_2_32 bitb_2_32 gnd C_bl
Rb_2_33 bit_2_33 bit_2_34 R_bl
Rbb_2_33 bitb_2_33 bitb_2_34 R_bl
Cb_2_33 bit_2_33 gnd C_bl
Cbb_2_33 bitb_2_33 gnd C_bl
Rb_2_34 bit_2_34 bit_2_35 R_bl
Rbb_2_34 bitb_2_34 bitb_2_35 R_bl
Cb_2_34 bit_2_34 gnd C_bl
Cbb_2_34 bitb_2_34 gnd C_bl
Rb_2_35 bit_2_35 bit_2_36 R_bl
Rbb_2_35 bitb_2_35 bitb_2_36 R_bl
Cb_2_35 bit_2_35 gnd C_bl
Cbb_2_35 bitb_2_35 gnd C_bl
Rb_2_36 bit_2_36 bit_2_37 R_bl
Rbb_2_36 bitb_2_36 bitb_2_37 R_bl
Cb_2_36 bit_2_36 gnd C_bl
Cbb_2_36 bitb_2_36 gnd C_bl
Rb_2_37 bit_2_37 bit_2_38 R_bl
Rbb_2_37 bitb_2_37 bitb_2_38 R_bl
Cb_2_37 bit_2_37 gnd C_bl
Cbb_2_37 bitb_2_37 gnd C_bl
Rb_2_38 bit_2_38 bit_2_39 R_bl
Rbb_2_38 bitb_2_38 bitb_2_39 R_bl
Cb_2_38 bit_2_38 gnd C_bl
Cbb_2_38 bitb_2_38 gnd C_bl
Rb_2_39 bit_2_39 bit_2_40 R_bl
Rbb_2_39 bitb_2_39 bitb_2_40 R_bl
Cb_2_39 bit_2_39 gnd C_bl
Cbb_2_39 bitb_2_39 gnd C_bl
Rb_2_40 bit_2_40 bit_2_41 R_bl
Rbb_2_40 bitb_2_40 bitb_2_41 R_bl
Cb_2_40 bit_2_40 gnd C_bl
Cbb_2_40 bitb_2_40 gnd C_bl
Rb_2_41 bit_2_41 bit_2_42 R_bl
Rbb_2_41 bitb_2_41 bitb_2_42 R_bl
Cb_2_41 bit_2_41 gnd C_bl
Cbb_2_41 bitb_2_41 gnd C_bl
Rb_2_42 bit_2_42 bit_2_43 R_bl
Rbb_2_42 bitb_2_42 bitb_2_43 R_bl
Cb_2_42 bit_2_42 gnd C_bl
Cbb_2_42 bitb_2_42 gnd C_bl
Rb_2_43 bit_2_43 bit_2_44 R_bl
Rbb_2_43 bitb_2_43 bitb_2_44 R_bl
Cb_2_43 bit_2_43 gnd C_bl
Cbb_2_43 bitb_2_43 gnd C_bl
Rb_2_44 bit_2_44 bit_2_45 R_bl
Rbb_2_44 bitb_2_44 bitb_2_45 R_bl
Cb_2_44 bit_2_44 gnd C_bl
Cbb_2_44 bitb_2_44 gnd C_bl
Rb_2_45 bit_2_45 bit_2_46 R_bl
Rbb_2_45 bitb_2_45 bitb_2_46 R_bl
Cb_2_45 bit_2_45 gnd C_bl
Cbb_2_45 bitb_2_45 gnd C_bl
Rb_2_46 bit_2_46 bit_2_47 R_bl
Rbb_2_46 bitb_2_46 bitb_2_47 R_bl
Cb_2_46 bit_2_46 gnd C_bl
Cbb_2_46 bitb_2_46 gnd C_bl
Rb_2_47 bit_2_47 bit_2_48 R_bl
Rbb_2_47 bitb_2_47 bitb_2_48 R_bl
Cb_2_47 bit_2_47 gnd C_bl
Cbb_2_47 bitb_2_47 gnd C_bl
Rb_2_48 bit_2_48 bit_2_49 R_bl
Rbb_2_48 bitb_2_48 bitb_2_49 R_bl
Cb_2_48 bit_2_48 gnd C_bl
Cbb_2_48 bitb_2_48 gnd C_bl
Rb_2_49 bit_2_49 bit_2_50 R_bl
Rbb_2_49 bitb_2_49 bitb_2_50 R_bl
Cb_2_49 bit_2_49 gnd C_bl
Cbb_2_49 bitb_2_49 gnd C_bl
Rb_2_50 bit_2_50 bit_2_51 R_bl
Rbb_2_50 bitb_2_50 bitb_2_51 R_bl
Cb_2_50 bit_2_50 gnd C_bl
Cbb_2_50 bitb_2_50 gnd C_bl
Rb_2_51 bit_2_51 bit_2_52 R_bl
Rbb_2_51 bitb_2_51 bitb_2_52 R_bl
Cb_2_51 bit_2_51 gnd C_bl
Cbb_2_51 bitb_2_51 gnd C_bl
Rb_2_52 bit_2_52 bit_2_53 R_bl
Rbb_2_52 bitb_2_52 bitb_2_53 R_bl
Cb_2_52 bit_2_52 gnd C_bl
Cbb_2_52 bitb_2_52 gnd C_bl
Rb_2_53 bit_2_53 bit_2_54 R_bl
Rbb_2_53 bitb_2_53 bitb_2_54 R_bl
Cb_2_53 bit_2_53 gnd C_bl
Cbb_2_53 bitb_2_53 gnd C_bl
Rb_2_54 bit_2_54 bit_2_55 R_bl
Rbb_2_54 bitb_2_54 bitb_2_55 R_bl
Cb_2_54 bit_2_54 gnd C_bl
Cbb_2_54 bitb_2_54 gnd C_bl
Rb_2_55 bit_2_55 bit_2_56 R_bl
Rbb_2_55 bitb_2_55 bitb_2_56 R_bl
Cb_2_55 bit_2_55 gnd C_bl
Cbb_2_55 bitb_2_55 gnd C_bl
Rb_2_56 bit_2_56 bit_2_57 R_bl
Rbb_2_56 bitb_2_56 bitb_2_57 R_bl
Cb_2_56 bit_2_56 gnd C_bl
Cbb_2_56 bitb_2_56 gnd C_bl
Rb_2_57 bit_2_57 bit_2_58 R_bl
Rbb_2_57 bitb_2_57 bitb_2_58 R_bl
Cb_2_57 bit_2_57 gnd C_bl
Cbb_2_57 bitb_2_57 gnd C_bl
Rb_2_58 bit_2_58 bit_2_59 R_bl
Rbb_2_58 bitb_2_58 bitb_2_59 R_bl
Cb_2_58 bit_2_58 gnd C_bl
Cbb_2_58 bitb_2_58 gnd C_bl
Rb_2_59 bit_2_59 bit_2_60 R_bl
Rbb_2_59 bitb_2_59 bitb_2_60 R_bl
Cb_2_59 bit_2_59 gnd C_bl
Cbb_2_59 bitb_2_59 gnd C_bl
Rb_2_60 bit_2_60 bit_2_61 R_bl
Rbb_2_60 bitb_2_60 bitb_2_61 R_bl
Cb_2_60 bit_2_60 gnd C_bl
Cbb_2_60 bitb_2_60 gnd C_bl
Rb_2_61 bit_2_61 bit_2_62 R_bl
Rbb_2_61 bitb_2_61 bitb_2_62 R_bl
Cb_2_61 bit_2_61 gnd C_bl
Cbb_2_61 bitb_2_61 gnd C_bl
Rb_2_62 bit_2_62 bit_2_63 R_bl
Rbb_2_62 bitb_2_62 bitb_2_63 R_bl
Cb_2_62 bit_2_62 gnd C_bl
Cbb_2_62 bitb_2_62 gnd C_bl
Rb_2_63 bit_2_63 bit_2_64 R_bl
Rbb_2_63 bitb_2_63 bitb_2_64 R_bl
Cb_2_63 bit_2_63 gnd C_bl
Cbb_2_63 bitb_2_63 gnd C_bl
Rb_2_64 bit_2_64 bit_2_65 R_bl
Rbb_2_64 bitb_2_64 bitb_2_65 R_bl
Cb_2_64 bit_2_64 gnd C_bl
Cbb_2_64 bitb_2_64 gnd C_bl
Rb_2_65 bit_2_65 bit_2_66 R_bl
Rbb_2_65 bitb_2_65 bitb_2_66 R_bl
Cb_2_65 bit_2_65 gnd C_bl
Cbb_2_65 bitb_2_65 gnd C_bl
Rb_2_66 bit_2_66 bit_2_67 R_bl
Rbb_2_66 bitb_2_66 bitb_2_67 R_bl
Cb_2_66 bit_2_66 gnd C_bl
Cbb_2_66 bitb_2_66 gnd C_bl
Rb_2_67 bit_2_67 bit_2_68 R_bl
Rbb_2_67 bitb_2_67 bitb_2_68 R_bl
Cb_2_67 bit_2_67 gnd C_bl
Cbb_2_67 bitb_2_67 gnd C_bl
Rb_2_68 bit_2_68 bit_2_69 R_bl
Rbb_2_68 bitb_2_68 bitb_2_69 R_bl
Cb_2_68 bit_2_68 gnd C_bl
Cbb_2_68 bitb_2_68 gnd C_bl
Rb_2_69 bit_2_69 bit_2_70 R_bl
Rbb_2_69 bitb_2_69 bitb_2_70 R_bl
Cb_2_69 bit_2_69 gnd C_bl
Cbb_2_69 bitb_2_69 gnd C_bl
Rb_2_70 bit_2_70 bit_2_71 R_bl
Rbb_2_70 bitb_2_70 bitb_2_71 R_bl
Cb_2_70 bit_2_70 gnd C_bl
Cbb_2_70 bitb_2_70 gnd C_bl
Rb_2_71 bit_2_71 bit_2_72 R_bl
Rbb_2_71 bitb_2_71 bitb_2_72 R_bl
Cb_2_71 bit_2_71 gnd C_bl
Cbb_2_71 bitb_2_71 gnd C_bl
Rb_2_72 bit_2_72 bit_2_73 R_bl
Rbb_2_72 bitb_2_72 bitb_2_73 R_bl
Cb_2_72 bit_2_72 gnd C_bl
Cbb_2_72 bitb_2_72 gnd C_bl
Rb_2_73 bit_2_73 bit_2_74 R_bl
Rbb_2_73 bitb_2_73 bitb_2_74 R_bl
Cb_2_73 bit_2_73 gnd C_bl
Cbb_2_73 bitb_2_73 gnd C_bl
Rb_2_74 bit_2_74 bit_2_75 R_bl
Rbb_2_74 bitb_2_74 bitb_2_75 R_bl
Cb_2_74 bit_2_74 gnd C_bl
Cbb_2_74 bitb_2_74 gnd C_bl
Rb_2_75 bit_2_75 bit_2_76 R_bl
Rbb_2_75 bitb_2_75 bitb_2_76 R_bl
Cb_2_75 bit_2_75 gnd C_bl
Cbb_2_75 bitb_2_75 gnd C_bl
Rb_2_76 bit_2_76 bit_2_77 R_bl
Rbb_2_76 bitb_2_76 bitb_2_77 R_bl
Cb_2_76 bit_2_76 gnd C_bl
Cbb_2_76 bitb_2_76 gnd C_bl
Rb_2_77 bit_2_77 bit_2_78 R_bl
Rbb_2_77 bitb_2_77 bitb_2_78 R_bl
Cb_2_77 bit_2_77 gnd C_bl
Cbb_2_77 bitb_2_77 gnd C_bl
Rb_2_78 bit_2_78 bit_2_79 R_bl
Rbb_2_78 bitb_2_78 bitb_2_79 R_bl
Cb_2_78 bit_2_78 gnd C_bl
Cbb_2_78 bitb_2_78 gnd C_bl
Rb_2_79 bit_2_79 bit_2_80 R_bl
Rbb_2_79 bitb_2_79 bitb_2_80 R_bl
Cb_2_79 bit_2_79 gnd C_bl
Cbb_2_79 bitb_2_79 gnd C_bl
Rb_2_80 bit_2_80 bit_2_81 R_bl
Rbb_2_80 bitb_2_80 bitb_2_81 R_bl
Cb_2_80 bit_2_80 gnd C_bl
Cbb_2_80 bitb_2_80 gnd C_bl
Rb_2_81 bit_2_81 bit_2_82 R_bl
Rbb_2_81 bitb_2_81 bitb_2_82 R_bl
Cb_2_81 bit_2_81 gnd C_bl
Cbb_2_81 bitb_2_81 gnd C_bl
Rb_2_82 bit_2_82 bit_2_83 R_bl
Rbb_2_82 bitb_2_82 bitb_2_83 R_bl
Cb_2_82 bit_2_82 gnd C_bl
Cbb_2_82 bitb_2_82 gnd C_bl
Rb_2_83 bit_2_83 bit_2_84 R_bl
Rbb_2_83 bitb_2_83 bitb_2_84 R_bl
Cb_2_83 bit_2_83 gnd C_bl
Cbb_2_83 bitb_2_83 gnd C_bl
Rb_2_84 bit_2_84 bit_2_85 R_bl
Rbb_2_84 bitb_2_84 bitb_2_85 R_bl
Cb_2_84 bit_2_84 gnd C_bl
Cbb_2_84 bitb_2_84 gnd C_bl
Rb_2_85 bit_2_85 bit_2_86 R_bl
Rbb_2_85 bitb_2_85 bitb_2_86 R_bl
Cb_2_85 bit_2_85 gnd C_bl
Cbb_2_85 bitb_2_85 gnd C_bl
Rb_2_86 bit_2_86 bit_2_87 R_bl
Rbb_2_86 bitb_2_86 bitb_2_87 R_bl
Cb_2_86 bit_2_86 gnd C_bl
Cbb_2_86 bitb_2_86 gnd C_bl
Rb_2_87 bit_2_87 bit_2_88 R_bl
Rbb_2_87 bitb_2_87 bitb_2_88 R_bl
Cb_2_87 bit_2_87 gnd C_bl
Cbb_2_87 bitb_2_87 gnd C_bl
Rb_2_88 bit_2_88 bit_2_89 R_bl
Rbb_2_88 bitb_2_88 bitb_2_89 R_bl
Cb_2_88 bit_2_88 gnd C_bl
Cbb_2_88 bitb_2_88 gnd C_bl
Rb_2_89 bit_2_89 bit_2_90 R_bl
Rbb_2_89 bitb_2_89 bitb_2_90 R_bl
Cb_2_89 bit_2_89 gnd C_bl
Cbb_2_89 bitb_2_89 gnd C_bl
Rb_2_90 bit_2_90 bit_2_91 R_bl
Rbb_2_90 bitb_2_90 bitb_2_91 R_bl
Cb_2_90 bit_2_90 gnd C_bl
Cbb_2_90 bitb_2_90 gnd C_bl
Rb_2_91 bit_2_91 bit_2_92 R_bl
Rbb_2_91 bitb_2_91 bitb_2_92 R_bl
Cb_2_91 bit_2_91 gnd C_bl
Cbb_2_91 bitb_2_91 gnd C_bl
Rb_2_92 bit_2_92 bit_2_93 R_bl
Rbb_2_92 bitb_2_92 bitb_2_93 R_bl
Cb_2_92 bit_2_92 gnd C_bl
Cbb_2_92 bitb_2_92 gnd C_bl
Rb_2_93 bit_2_93 bit_2_94 R_bl
Rbb_2_93 bitb_2_93 bitb_2_94 R_bl
Cb_2_93 bit_2_93 gnd C_bl
Cbb_2_93 bitb_2_93 gnd C_bl
Rb_2_94 bit_2_94 bit_2_95 R_bl
Rbb_2_94 bitb_2_94 bitb_2_95 R_bl
Cb_2_94 bit_2_94 gnd C_bl
Cbb_2_94 bitb_2_94 gnd C_bl
Rb_2_95 bit_2_95 bit_2_96 R_bl
Rbb_2_95 bitb_2_95 bitb_2_96 R_bl
Cb_2_95 bit_2_95 gnd C_bl
Cbb_2_95 bitb_2_95 gnd C_bl
Rb_2_96 bit_2_96 bit_2_97 R_bl
Rbb_2_96 bitb_2_96 bitb_2_97 R_bl
Cb_2_96 bit_2_96 gnd C_bl
Cbb_2_96 bitb_2_96 gnd C_bl
Rb_2_97 bit_2_97 bit_2_98 R_bl
Rbb_2_97 bitb_2_97 bitb_2_98 R_bl
Cb_2_97 bit_2_97 gnd C_bl
Cbb_2_97 bitb_2_97 gnd C_bl
Rb_2_98 bit_2_98 bit_2_99 R_bl
Rbb_2_98 bitb_2_98 bitb_2_99 R_bl
Cb_2_98 bit_2_98 gnd C_bl
Cbb_2_98 bitb_2_98 gnd C_bl
Rb_2_99 bit_2_99 bit_2_100 R_bl
Rbb_2_99 bitb_2_99 bitb_2_100 R_bl
Cb_2_99 bit_2_99 gnd C_bl
Cbb_2_99 bitb_2_99 gnd C_bl
Rb_3_0 bit_3_0 bit_3_1 R_bl
Rbb_3_0 bitb_3_0 bitb_3_1 R_bl
Cb_3_0 bit_3_0 gnd C_bl
Cbb_3_0 bitb_3_0 gnd C_bl
Rb_3_1 bit_3_1 bit_3_2 R_bl
Rbb_3_1 bitb_3_1 bitb_3_2 R_bl
Cb_3_1 bit_3_1 gnd C_bl
Cbb_3_1 bitb_3_1 gnd C_bl
Rb_3_2 bit_3_2 bit_3_3 R_bl
Rbb_3_2 bitb_3_2 bitb_3_3 R_bl
Cb_3_2 bit_3_2 gnd C_bl
Cbb_3_2 bitb_3_2 gnd C_bl
Rb_3_3 bit_3_3 bit_3_4 R_bl
Rbb_3_3 bitb_3_3 bitb_3_4 R_bl
Cb_3_3 bit_3_3 gnd C_bl
Cbb_3_3 bitb_3_3 gnd C_bl
Rb_3_4 bit_3_4 bit_3_5 R_bl
Rbb_3_4 bitb_3_4 bitb_3_5 R_bl
Cb_3_4 bit_3_4 gnd C_bl
Cbb_3_4 bitb_3_4 gnd C_bl
Rb_3_5 bit_3_5 bit_3_6 R_bl
Rbb_3_5 bitb_3_5 bitb_3_6 R_bl
Cb_3_5 bit_3_5 gnd C_bl
Cbb_3_5 bitb_3_5 gnd C_bl
Rb_3_6 bit_3_6 bit_3_7 R_bl
Rbb_3_6 bitb_3_6 bitb_3_7 R_bl
Cb_3_6 bit_3_6 gnd C_bl
Cbb_3_6 bitb_3_6 gnd C_bl
Rb_3_7 bit_3_7 bit_3_8 R_bl
Rbb_3_7 bitb_3_7 bitb_3_8 R_bl
Cb_3_7 bit_3_7 gnd C_bl
Cbb_3_7 bitb_3_7 gnd C_bl
Rb_3_8 bit_3_8 bit_3_9 R_bl
Rbb_3_8 bitb_3_8 bitb_3_9 R_bl
Cb_3_8 bit_3_8 gnd C_bl
Cbb_3_8 bitb_3_8 gnd C_bl
Rb_3_9 bit_3_9 bit_3_10 R_bl
Rbb_3_9 bitb_3_9 bitb_3_10 R_bl
Cb_3_9 bit_3_9 gnd C_bl
Cbb_3_9 bitb_3_9 gnd C_bl
Rb_3_10 bit_3_10 bit_3_11 R_bl
Rbb_3_10 bitb_3_10 bitb_3_11 R_bl
Cb_3_10 bit_3_10 gnd C_bl
Cbb_3_10 bitb_3_10 gnd C_bl
Rb_3_11 bit_3_11 bit_3_12 R_bl
Rbb_3_11 bitb_3_11 bitb_3_12 R_bl
Cb_3_11 bit_3_11 gnd C_bl
Cbb_3_11 bitb_3_11 gnd C_bl
Rb_3_12 bit_3_12 bit_3_13 R_bl
Rbb_3_12 bitb_3_12 bitb_3_13 R_bl
Cb_3_12 bit_3_12 gnd C_bl
Cbb_3_12 bitb_3_12 gnd C_bl
Rb_3_13 bit_3_13 bit_3_14 R_bl
Rbb_3_13 bitb_3_13 bitb_3_14 R_bl
Cb_3_13 bit_3_13 gnd C_bl
Cbb_3_13 bitb_3_13 gnd C_bl
Rb_3_14 bit_3_14 bit_3_15 R_bl
Rbb_3_14 bitb_3_14 bitb_3_15 R_bl
Cb_3_14 bit_3_14 gnd C_bl
Cbb_3_14 bitb_3_14 gnd C_bl
Rb_3_15 bit_3_15 bit_3_16 R_bl
Rbb_3_15 bitb_3_15 bitb_3_16 R_bl
Cb_3_15 bit_3_15 gnd C_bl
Cbb_3_15 bitb_3_15 gnd C_bl
Rb_3_16 bit_3_16 bit_3_17 R_bl
Rbb_3_16 bitb_3_16 bitb_3_17 R_bl
Cb_3_16 bit_3_16 gnd C_bl
Cbb_3_16 bitb_3_16 gnd C_bl
Rb_3_17 bit_3_17 bit_3_18 R_bl
Rbb_3_17 bitb_3_17 bitb_3_18 R_bl
Cb_3_17 bit_3_17 gnd C_bl
Cbb_3_17 bitb_3_17 gnd C_bl
Rb_3_18 bit_3_18 bit_3_19 R_bl
Rbb_3_18 bitb_3_18 bitb_3_19 R_bl
Cb_3_18 bit_3_18 gnd C_bl
Cbb_3_18 bitb_3_18 gnd C_bl
Rb_3_19 bit_3_19 bit_3_20 R_bl
Rbb_3_19 bitb_3_19 bitb_3_20 R_bl
Cb_3_19 bit_3_19 gnd C_bl
Cbb_3_19 bitb_3_19 gnd C_bl
Rb_3_20 bit_3_20 bit_3_21 R_bl
Rbb_3_20 bitb_3_20 bitb_3_21 R_bl
Cb_3_20 bit_3_20 gnd C_bl
Cbb_3_20 bitb_3_20 gnd C_bl
Rb_3_21 bit_3_21 bit_3_22 R_bl
Rbb_3_21 bitb_3_21 bitb_3_22 R_bl
Cb_3_21 bit_3_21 gnd C_bl
Cbb_3_21 bitb_3_21 gnd C_bl
Rb_3_22 bit_3_22 bit_3_23 R_bl
Rbb_3_22 bitb_3_22 bitb_3_23 R_bl
Cb_3_22 bit_3_22 gnd C_bl
Cbb_3_22 bitb_3_22 gnd C_bl
Rb_3_23 bit_3_23 bit_3_24 R_bl
Rbb_3_23 bitb_3_23 bitb_3_24 R_bl
Cb_3_23 bit_3_23 gnd C_bl
Cbb_3_23 bitb_3_23 gnd C_bl
Rb_3_24 bit_3_24 bit_3_25 R_bl
Rbb_3_24 bitb_3_24 bitb_3_25 R_bl
Cb_3_24 bit_3_24 gnd C_bl
Cbb_3_24 bitb_3_24 gnd C_bl
Rb_3_25 bit_3_25 bit_3_26 R_bl
Rbb_3_25 bitb_3_25 bitb_3_26 R_bl
Cb_3_25 bit_3_25 gnd C_bl
Cbb_3_25 bitb_3_25 gnd C_bl
Rb_3_26 bit_3_26 bit_3_27 R_bl
Rbb_3_26 bitb_3_26 bitb_3_27 R_bl
Cb_3_26 bit_3_26 gnd C_bl
Cbb_3_26 bitb_3_26 gnd C_bl
Rb_3_27 bit_3_27 bit_3_28 R_bl
Rbb_3_27 bitb_3_27 bitb_3_28 R_bl
Cb_3_27 bit_3_27 gnd C_bl
Cbb_3_27 bitb_3_27 gnd C_bl
Rb_3_28 bit_3_28 bit_3_29 R_bl
Rbb_3_28 bitb_3_28 bitb_3_29 R_bl
Cb_3_28 bit_3_28 gnd C_bl
Cbb_3_28 bitb_3_28 gnd C_bl
Rb_3_29 bit_3_29 bit_3_30 R_bl
Rbb_3_29 bitb_3_29 bitb_3_30 R_bl
Cb_3_29 bit_3_29 gnd C_bl
Cbb_3_29 bitb_3_29 gnd C_bl
Rb_3_30 bit_3_30 bit_3_31 R_bl
Rbb_3_30 bitb_3_30 bitb_3_31 R_bl
Cb_3_30 bit_3_30 gnd C_bl
Cbb_3_30 bitb_3_30 gnd C_bl
Rb_3_31 bit_3_31 bit_3_32 R_bl
Rbb_3_31 bitb_3_31 bitb_3_32 R_bl
Cb_3_31 bit_3_31 gnd C_bl
Cbb_3_31 bitb_3_31 gnd C_bl
Rb_3_32 bit_3_32 bit_3_33 R_bl
Rbb_3_32 bitb_3_32 bitb_3_33 R_bl
Cb_3_32 bit_3_32 gnd C_bl
Cbb_3_32 bitb_3_32 gnd C_bl
Rb_3_33 bit_3_33 bit_3_34 R_bl
Rbb_3_33 bitb_3_33 bitb_3_34 R_bl
Cb_3_33 bit_3_33 gnd C_bl
Cbb_3_33 bitb_3_33 gnd C_bl
Rb_3_34 bit_3_34 bit_3_35 R_bl
Rbb_3_34 bitb_3_34 bitb_3_35 R_bl
Cb_3_34 bit_3_34 gnd C_bl
Cbb_3_34 bitb_3_34 gnd C_bl
Rb_3_35 bit_3_35 bit_3_36 R_bl
Rbb_3_35 bitb_3_35 bitb_3_36 R_bl
Cb_3_35 bit_3_35 gnd C_bl
Cbb_3_35 bitb_3_35 gnd C_bl
Rb_3_36 bit_3_36 bit_3_37 R_bl
Rbb_3_36 bitb_3_36 bitb_3_37 R_bl
Cb_3_36 bit_3_36 gnd C_bl
Cbb_3_36 bitb_3_36 gnd C_bl
Rb_3_37 bit_3_37 bit_3_38 R_bl
Rbb_3_37 bitb_3_37 bitb_3_38 R_bl
Cb_3_37 bit_3_37 gnd C_bl
Cbb_3_37 bitb_3_37 gnd C_bl
Rb_3_38 bit_3_38 bit_3_39 R_bl
Rbb_3_38 bitb_3_38 bitb_3_39 R_bl
Cb_3_38 bit_3_38 gnd C_bl
Cbb_3_38 bitb_3_38 gnd C_bl
Rb_3_39 bit_3_39 bit_3_40 R_bl
Rbb_3_39 bitb_3_39 bitb_3_40 R_bl
Cb_3_39 bit_3_39 gnd C_bl
Cbb_3_39 bitb_3_39 gnd C_bl
Rb_3_40 bit_3_40 bit_3_41 R_bl
Rbb_3_40 bitb_3_40 bitb_3_41 R_bl
Cb_3_40 bit_3_40 gnd C_bl
Cbb_3_40 bitb_3_40 gnd C_bl
Rb_3_41 bit_3_41 bit_3_42 R_bl
Rbb_3_41 bitb_3_41 bitb_3_42 R_bl
Cb_3_41 bit_3_41 gnd C_bl
Cbb_3_41 bitb_3_41 gnd C_bl
Rb_3_42 bit_3_42 bit_3_43 R_bl
Rbb_3_42 bitb_3_42 bitb_3_43 R_bl
Cb_3_42 bit_3_42 gnd C_bl
Cbb_3_42 bitb_3_42 gnd C_bl
Rb_3_43 bit_3_43 bit_3_44 R_bl
Rbb_3_43 bitb_3_43 bitb_3_44 R_bl
Cb_3_43 bit_3_43 gnd C_bl
Cbb_3_43 bitb_3_43 gnd C_bl
Rb_3_44 bit_3_44 bit_3_45 R_bl
Rbb_3_44 bitb_3_44 bitb_3_45 R_bl
Cb_3_44 bit_3_44 gnd C_bl
Cbb_3_44 bitb_3_44 gnd C_bl
Rb_3_45 bit_3_45 bit_3_46 R_bl
Rbb_3_45 bitb_3_45 bitb_3_46 R_bl
Cb_3_45 bit_3_45 gnd C_bl
Cbb_3_45 bitb_3_45 gnd C_bl
Rb_3_46 bit_3_46 bit_3_47 R_bl
Rbb_3_46 bitb_3_46 bitb_3_47 R_bl
Cb_3_46 bit_3_46 gnd C_bl
Cbb_3_46 bitb_3_46 gnd C_bl
Rb_3_47 bit_3_47 bit_3_48 R_bl
Rbb_3_47 bitb_3_47 bitb_3_48 R_bl
Cb_3_47 bit_3_47 gnd C_bl
Cbb_3_47 bitb_3_47 gnd C_bl
Rb_3_48 bit_3_48 bit_3_49 R_bl
Rbb_3_48 bitb_3_48 bitb_3_49 R_bl
Cb_3_48 bit_3_48 gnd C_bl
Cbb_3_48 bitb_3_48 gnd C_bl
Rb_3_49 bit_3_49 bit_3_50 R_bl
Rbb_3_49 bitb_3_49 bitb_3_50 R_bl
Cb_3_49 bit_3_49 gnd C_bl
Cbb_3_49 bitb_3_49 gnd C_bl
Rb_3_50 bit_3_50 bit_3_51 R_bl
Rbb_3_50 bitb_3_50 bitb_3_51 R_bl
Cb_3_50 bit_3_50 gnd C_bl
Cbb_3_50 bitb_3_50 gnd C_bl
Rb_3_51 bit_3_51 bit_3_52 R_bl
Rbb_3_51 bitb_3_51 bitb_3_52 R_bl
Cb_3_51 bit_3_51 gnd C_bl
Cbb_3_51 bitb_3_51 gnd C_bl
Rb_3_52 bit_3_52 bit_3_53 R_bl
Rbb_3_52 bitb_3_52 bitb_3_53 R_bl
Cb_3_52 bit_3_52 gnd C_bl
Cbb_3_52 bitb_3_52 gnd C_bl
Rb_3_53 bit_3_53 bit_3_54 R_bl
Rbb_3_53 bitb_3_53 bitb_3_54 R_bl
Cb_3_53 bit_3_53 gnd C_bl
Cbb_3_53 bitb_3_53 gnd C_bl
Rb_3_54 bit_3_54 bit_3_55 R_bl
Rbb_3_54 bitb_3_54 bitb_3_55 R_bl
Cb_3_54 bit_3_54 gnd C_bl
Cbb_3_54 bitb_3_54 gnd C_bl
Rb_3_55 bit_3_55 bit_3_56 R_bl
Rbb_3_55 bitb_3_55 bitb_3_56 R_bl
Cb_3_55 bit_3_55 gnd C_bl
Cbb_3_55 bitb_3_55 gnd C_bl
Rb_3_56 bit_3_56 bit_3_57 R_bl
Rbb_3_56 bitb_3_56 bitb_3_57 R_bl
Cb_3_56 bit_3_56 gnd C_bl
Cbb_3_56 bitb_3_56 gnd C_bl
Rb_3_57 bit_3_57 bit_3_58 R_bl
Rbb_3_57 bitb_3_57 bitb_3_58 R_bl
Cb_3_57 bit_3_57 gnd C_bl
Cbb_3_57 bitb_3_57 gnd C_bl
Rb_3_58 bit_3_58 bit_3_59 R_bl
Rbb_3_58 bitb_3_58 bitb_3_59 R_bl
Cb_3_58 bit_3_58 gnd C_bl
Cbb_3_58 bitb_3_58 gnd C_bl
Rb_3_59 bit_3_59 bit_3_60 R_bl
Rbb_3_59 bitb_3_59 bitb_3_60 R_bl
Cb_3_59 bit_3_59 gnd C_bl
Cbb_3_59 bitb_3_59 gnd C_bl
Rb_3_60 bit_3_60 bit_3_61 R_bl
Rbb_3_60 bitb_3_60 bitb_3_61 R_bl
Cb_3_60 bit_3_60 gnd C_bl
Cbb_3_60 bitb_3_60 gnd C_bl
Rb_3_61 bit_3_61 bit_3_62 R_bl
Rbb_3_61 bitb_3_61 bitb_3_62 R_bl
Cb_3_61 bit_3_61 gnd C_bl
Cbb_3_61 bitb_3_61 gnd C_bl
Rb_3_62 bit_3_62 bit_3_63 R_bl
Rbb_3_62 bitb_3_62 bitb_3_63 R_bl
Cb_3_62 bit_3_62 gnd C_bl
Cbb_3_62 bitb_3_62 gnd C_bl
Rb_3_63 bit_3_63 bit_3_64 R_bl
Rbb_3_63 bitb_3_63 bitb_3_64 R_bl
Cb_3_63 bit_3_63 gnd C_bl
Cbb_3_63 bitb_3_63 gnd C_bl
Rb_3_64 bit_3_64 bit_3_65 R_bl
Rbb_3_64 bitb_3_64 bitb_3_65 R_bl
Cb_3_64 bit_3_64 gnd C_bl
Cbb_3_64 bitb_3_64 gnd C_bl
Rb_3_65 bit_3_65 bit_3_66 R_bl
Rbb_3_65 bitb_3_65 bitb_3_66 R_bl
Cb_3_65 bit_3_65 gnd C_bl
Cbb_3_65 bitb_3_65 gnd C_bl
Rb_3_66 bit_3_66 bit_3_67 R_bl
Rbb_3_66 bitb_3_66 bitb_3_67 R_bl
Cb_3_66 bit_3_66 gnd C_bl
Cbb_3_66 bitb_3_66 gnd C_bl
Rb_3_67 bit_3_67 bit_3_68 R_bl
Rbb_3_67 bitb_3_67 bitb_3_68 R_bl
Cb_3_67 bit_3_67 gnd C_bl
Cbb_3_67 bitb_3_67 gnd C_bl
Rb_3_68 bit_3_68 bit_3_69 R_bl
Rbb_3_68 bitb_3_68 bitb_3_69 R_bl
Cb_3_68 bit_3_68 gnd C_bl
Cbb_3_68 bitb_3_68 gnd C_bl
Rb_3_69 bit_3_69 bit_3_70 R_bl
Rbb_3_69 bitb_3_69 bitb_3_70 R_bl
Cb_3_69 bit_3_69 gnd C_bl
Cbb_3_69 bitb_3_69 gnd C_bl
Rb_3_70 bit_3_70 bit_3_71 R_bl
Rbb_3_70 bitb_3_70 bitb_3_71 R_bl
Cb_3_70 bit_3_70 gnd C_bl
Cbb_3_70 bitb_3_70 gnd C_bl
Rb_3_71 bit_3_71 bit_3_72 R_bl
Rbb_3_71 bitb_3_71 bitb_3_72 R_bl
Cb_3_71 bit_3_71 gnd C_bl
Cbb_3_71 bitb_3_71 gnd C_bl
Rb_3_72 bit_3_72 bit_3_73 R_bl
Rbb_3_72 bitb_3_72 bitb_3_73 R_bl
Cb_3_72 bit_3_72 gnd C_bl
Cbb_3_72 bitb_3_72 gnd C_bl
Rb_3_73 bit_3_73 bit_3_74 R_bl
Rbb_3_73 bitb_3_73 bitb_3_74 R_bl
Cb_3_73 bit_3_73 gnd C_bl
Cbb_3_73 bitb_3_73 gnd C_bl
Rb_3_74 bit_3_74 bit_3_75 R_bl
Rbb_3_74 bitb_3_74 bitb_3_75 R_bl
Cb_3_74 bit_3_74 gnd C_bl
Cbb_3_74 bitb_3_74 gnd C_bl
Rb_3_75 bit_3_75 bit_3_76 R_bl
Rbb_3_75 bitb_3_75 bitb_3_76 R_bl
Cb_3_75 bit_3_75 gnd C_bl
Cbb_3_75 bitb_3_75 gnd C_bl
Rb_3_76 bit_3_76 bit_3_77 R_bl
Rbb_3_76 bitb_3_76 bitb_3_77 R_bl
Cb_3_76 bit_3_76 gnd C_bl
Cbb_3_76 bitb_3_76 gnd C_bl
Rb_3_77 bit_3_77 bit_3_78 R_bl
Rbb_3_77 bitb_3_77 bitb_3_78 R_bl
Cb_3_77 bit_3_77 gnd C_bl
Cbb_3_77 bitb_3_77 gnd C_bl
Rb_3_78 bit_3_78 bit_3_79 R_bl
Rbb_3_78 bitb_3_78 bitb_3_79 R_bl
Cb_3_78 bit_3_78 gnd C_bl
Cbb_3_78 bitb_3_78 gnd C_bl
Rb_3_79 bit_3_79 bit_3_80 R_bl
Rbb_3_79 bitb_3_79 bitb_3_80 R_bl
Cb_3_79 bit_3_79 gnd C_bl
Cbb_3_79 bitb_3_79 gnd C_bl
Rb_3_80 bit_3_80 bit_3_81 R_bl
Rbb_3_80 bitb_3_80 bitb_3_81 R_bl
Cb_3_80 bit_3_80 gnd C_bl
Cbb_3_80 bitb_3_80 gnd C_bl
Rb_3_81 bit_3_81 bit_3_82 R_bl
Rbb_3_81 bitb_3_81 bitb_3_82 R_bl
Cb_3_81 bit_3_81 gnd C_bl
Cbb_3_81 bitb_3_81 gnd C_bl
Rb_3_82 bit_3_82 bit_3_83 R_bl
Rbb_3_82 bitb_3_82 bitb_3_83 R_bl
Cb_3_82 bit_3_82 gnd C_bl
Cbb_3_82 bitb_3_82 gnd C_bl
Rb_3_83 bit_3_83 bit_3_84 R_bl
Rbb_3_83 bitb_3_83 bitb_3_84 R_bl
Cb_3_83 bit_3_83 gnd C_bl
Cbb_3_83 bitb_3_83 gnd C_bl
Rb_3_84 bit_3_84 bit_3_85 R_bl
Rbb_3_84 bitb_3_84 bitb_3_85 R_bl
Cb_3_84 bit_3_84 gnd C_bl
Cbb_3_84 bitb_3_84 gnd C_bl
Rb_3_85 bit_3_85 bit_3_86 R_bl
Rbb_3_85 bitb_3_85 bitb_3_86 R_bl
Cb_3_85 bit_3_85 gnd C_bl
Cbb_3_85 bitb_3_85 gnd C_bl
Rb_3_86 bit_3_86 bit_3_87 R_bl
Rbb_3_86 bitb_3_86 bitb_3_87 R_bl
Cb_3_86 bit_3_86 gnd C_bl
Cbb_3_86 bitb_3_86 gnd C_bl
Rb_3_87 bit_3_87 bit_3_88 R_bl
Rbb_3_87 bitb_3_87 bitb_3_88 R_bl
Cb_3_87 bit_3_87 gnd C_bl
Cbb_3_87 bitb_3_87 gnd C_bl
Rb_3_88 bit_3_88 bit_3_89 R_bl
Rbb_3_88 bitb_3_88 bitb_3_89 R_bl
Cb_3_88 bit_3_88 gnd C_bl
Cbb_3_88 bitb_3_88 gnd C_bl
Rb_3_89 bit_3_89 bit_3_90 R_bl
Rbb_3_89 bitb_3_89 bitb_3_90 R_bl
Cb_3_89 bit_3_89 gnd C_bl
Cbb_3_89 bitb_3_89 gnd C_bl
Rb_3_90 bit_3_90 bit_3_91 R_bl
Rbb_3_90 bitb_3_90 bitb_3_91 R_bl
Cb_3_90 bit_3_90 gnd C_bl
Cbb_3_90 bitb_3_90 gnd C_bl
Rb_3_91 bit_3_91 bit_3_92 R_bl
Rbb_3_91 bitb_3_91 bitb_3_92 R_bl
Cb_3_91 bit_3_91 gnd C_bl
Cbb_3_91 bitb_3_91 gnd C_bl
Rb_3_92 bit_3_92 bit_3_93 R_bl
Rbb_3_92 bitb_3_92 bitb_3_93 R_bl
Cb_3_92 bit_3_92 gnd C_bl
Cbb_3_92 bitb_3_92 gnd C_bl
Rb_3_93 bit_3_93 bit_3_94 R_bl
Rbb_3_93 bitb_3_93 bitb_3_94 R_bl
Cb_3_93 bit_3_93 gnd C_bl
Cbb_3_93 bitb_3_93 gnd C_bl
Rb_3_94 bit_3_94 bit_3_95 R_bl
Rbb_3_94 bitb_3_94 bitb_3_95 R_bl
Cb_3_94 bit_3_94 gnd C_bl
Cbb_3_94 bitb_3_94 gnd C_bl
Rb_3_95 bit_3_95 bit_3_96 R_bl
Rbb_3_95 bitb_3_95 bitb_3_96 R_bl
Cb_3_95 bit_3_95 gnd C_bl
Cbb_3_95 bitb_3_95 gnd C_bl
Rb_3_96 bit_3_96 bit_3_97 R_bl
Rbb_3_96 bitb_3_96 bitb_3_97 R_bl
Cb_3_96 bit_3_96 gnd C_bl
Cbb_3_96 bitb_3_96 gnd C_bl
Rb_3_97 bit_3_97 bit_3_98 R_bl
Rbb_3_97 bitb_3_97 bitb_3_98 R_bl
Cb_3_97 bit_3_97 gnd C_bl
Cbb_3_97 bitb_3_97 gnd C_bl
Rb_3_98 bit_3_98 bit_3_99 R_bl
Rbb_3_98 bitb_3_98 bitb_3_99 R_bl
Cb_3_98 bit_3_98 gnd C_bl
Cbb_3_98 bitb_3_98 gnd C_bl
Rb_3_99 bit_3_99 bit_3_100 R_bl
Rbb_3_99 bitb_3_99 bitb_3_100 R_bl
Cb_3_99 bit_3_99 gnd C_bl
Cbb_3_99 bitb_3_99 gnd C_bl
Rb_4_0 bit_4_0 bit_4_1 R_bl
Rbb_4_0 bitb_4_0 bitb_4_1 R_bl
Cb_4_0 bit_4_0 gnd C_bl
Cbb_4_0 bitb_4_0 gnd C_bl
Rb_4_1 bit_4_1 bit_4_2 R_bl
Rbb_4_1 bitb_4_1 bitb_4_2 R_bl
Cb_4_1 bit_4_1 gnd C_bl
Cbb_4_1 bitb_4_1 gnd C_bl
Rb_4_2 bit_4_2 bit_4_3 R_bl
Rbb_4_2 bitb_4_2 bitb_4_3 R_bl
Cb_4_2 bit_4_2 gnd C_bl
Cbb_4_2 bitb_4_2 gnd C_bl
Rb_4_3 bit_4_3 bit_4_4 R_bl
Rbb_4_3 bitb_4_3 bitb_4_4 R_bl
Cb_4_3 bit_4_3 gnd C_bl
Cbb_4_3 bitb_4_3 gnd C_bl
Rb_4_4 bit_4_4 bit_4_5 R_bl
Rbb_4_4 bitb_4_4 bitb_4_5 R_bl
Cb_4_4 bit_4_4 gnd C_bl
Cbb_4_4 bitb_4_4 gnd C_bl
Rb_4_5 bit_4_5 bit_4_6 R_bl
Rbb_4_5 bitb_4_5 bitb_4_6 R_bl
Cb_4_5 bit_4_5 gnd C_bl
Cbb_4_5 bitb_4_5 gnd C_bl
Rb_4_6 bit_4_6 bit_4_7 R_bl
Rbb_4_6 bitb_4_6 bitb_4_7 R_bl
Cb_4_6 bit_4_6 gnd C_bl
Cbb_4_6 bitb_4_6 gnd C_bl
Rb_4_7 bit_4_7 bit_4_8 R_bl
Rbb_4_7 bitb_4_7 bitb_4_8 R_bl
Cb_4_7 bit_4_7 gnd C_bl
Cbb_4_7 bitb_4_7 gnd C_bl
Rb_4_8 bit_4_8 bit_4_9 R_bl
Rbb_4_8 bitb_4_8 bitb_4_9 R_bl
Cb_4_8 bit_4_8 gnd C_bl
Cbb_4_8 bitb_4_8 gnd C_bl
Rb_4_9 bit_4_9 bit_4_10 R_bl
Rbb_4_9 bitb_4_9 bitb_4_10 R_bl
Cb_4_9 bit_4_9 gnd C_bl
Cbb_4_9 bitb_4_9 gnd C_bl
Rb_4_10 bit_4_10 bit_4_11 R_bl
Rbb_4_10 bitb_4_10 bitb_4_11 R_bl
Cb_4_10 bit_4_10 gnd C_bl
Cbb_4_10 bitb_4_10 gnd C_bl
Rb_4_11 bit_4_11 bit_4_12 R_bl
Rbb_4_11 bitb_4_11 bitb_4_12 R_bl
Cb_4_11 bit_4_11 gnd C_bl
Cbb_4_11 bitb_4_11 gnd C_bl
Rb_4_12 bit_4_12 bit_4_13 R_bl
Rbb_4_12 bitb_4_12 bitb_4_13 R_bl
Cb_4_12 bit_4_12 gnd C_bl
Cbb_4_12 bitb_4_12 gnd C_bl
Rb_4_13 bit_4_13 bit_4_14 R_bl
Rbb_4_13 bitb_4_13 bitb_4_14 R_bl
Cb_4_13 bit_4_13 gnd C_bl
Cbb_4_13 bitb_4_13 gnd C_bl
Rb_4_14 bit_4_14 bit_4_15 R_bl
Rbb_4_14 bitb_4_14 bitb_4_15 R_bl
Cb_4_14 bit_4_14 gnd C_bl
Cbb_4_14 bitb_4_14 gnd C_bl
Rb_4_15 bit_4_15 bit_4_16 R_bl
Rbb_4_15 bitb_4_15 bitb_4_16 R_bl
Cb_4_15 bit_4_15 gnd C_bl
Cbb_4_15 bitb_4_15 gnd C_bl
Rb_4_16 bit_4_16 bit_4_17 R_bl
Rbb_4_16 bitb_4_16 bitb_4_17 R_bl
Cb_4_16 bit_4_16 gnd C_bl
Cbb_4_16 bitb_4_16 gnd C_bl
Rb_4_17 bit_4_17 bit_4_18 R_bl
Rbb_4_17 bitb_4_17 bitb_4_18 R_bl
Cb_4_17 bit_4_17 gnd C_bl
Cbb_4_17 bitb_4_17 gnd C_bl
Rb_4_18 bit_4_18 bit_4_19 R_bl
Rbb_4_18 bitb_4_18 bitb_4_19 R_bl
Cb_4_18 bit_4_18 gnd C_bl
Cbb_4_18 bitb_4_18 gnd C_bl
Rb_4_19 bit_4_19 bit_4_20 R_bl
Rbb_4_19 bitb_4_19 bitb_4_20 R_bl
Cb_4_19 bit_4_19 gnd C_bl
Cbb_4_19 bitb_4_19 gnd C_bl
Rb_4_20 bit_4_20 bit_4_21 R_bl
Rbb_4_20 bitb_4_20 bitb_4_21 R_bl
Cb_4_20 bit_4_20 gnd C_bl
Cbb_4_20 bitb_4_20 gnd C_bl
Rb_4_21 bit_4_21 bit_4_22 R_bl
Rbb_4_21 bitb_4_21 bitb_4_22 R_bl
Cb_4_21 bit_4_21 gnd C_bl
Cbb_4_21 bitb_4_21 gnd C_bl
Rb_4_22 bit_4_22 bit_4_23 R_bl
Rbb_4_22 bitb_4_22 bitb_4_23 R_bl
Cb_4_22 bit_4_22 gnd C_bl
Cbb_4_22 bitb_4_22 gnd C_bl
Rb_4_23 bit_4_23 bit_4_24 R_bl
Rbb_4_23 bitb_4_23 bitb_4_24 R_bl
Cb_4_23 bit_4_23 gnd C_bl
Cbb_4_23 bitb_4_23 gnd C_bl
Rb_4_24 bit_4_24 bit_4_25 R_bl
Rbb_4_24 bitb_4_24 bitb_4_25 R_bl
Cb_4_24 bit_4_24 gnd C_bl
Cbb_4_24 bitb_4_24 gnd C_bl
Rb_4_25 bit_4_25 bit_4_26 R_bl
Rbb_4_25 bitb_4_25 bitb_4_26 R_bl
Cb_4_25 bit_4_25 gnd C_bl
Cbb_4_25 bitb_4_25 gnd C_bl
Rb_4_26 bit_4_26 bit_4_27 R_bl
Rbb_4_26 bitb_4_26 bitb_4_27 R_bl
Cb_4_26 bit_4_26 gnd C_bl
Cbb_4_26 bitb_4_26 gnd C_bl
Rb_4_27 bit_4_27 bit_4_28 R_bl
Rbb_4_27 bitb_4_27 bitb_4_28 R_bl
Cb_4_27 bit_4_27 gnd C_bl
Cbb_4_27 bitb_4_27 gnd C_bl
Rb_4_28 bit_4_28 bit_4_29 R_bl
Rbb_4_28 bitb_4_28 bitb_4_29 R_bl
Cb_4_28 bit_4_28 gnd C_bl
Cbb_4_28 bitb_4_28 gnd C_bl
Rb_4_29 bit_4_29 bit_4_30 R_bl
Rbb_4_29 bitb_4_29 bitb_4_30 R_bl
Cb_4_29 bit_4_29 gnd C_bl
Cbb_4_29 bitb_4_29 gnd C_bl
Rb_4_30 bit_4_30 bit_4_31 R_bl
Rbb_4_30 bitb_4_30 bitb_4_31 R_bl
Cb_4_30 bit_4_30 gnd C_bl
Cbb_4_30 bitb_4_30 gnd C_bl
Rb_4_31 bit_4_31 bit_4_32 R_bl
Rbb_4_31 bitb_4_31 bitb_4_32 R_bl
Cb_4_31 bit_4_31 gnd C_bl
Cbb_4_31 bitb_4_31 gnd C_bl
Rb_4_32 bit_4_32 bit_4_33 R_bl
Rbb_4_32 bitb_4_32 bitb_4_33 R_bl
Cb_4_32 bit_4_32 gnd C_bl
Cbb_4_32 bitb_4_32 gnd C_bl
Rb_4_33 bit_4_33 bit_4_34 R_bl
Rbb_4_33 bitb_4_33 bitb_4_34 R_bl
Cb_4_33 bit_4_33 gnd C_bl
Cbb_4_33 bitb_4_33 gnd C_bl
Rb_4_34 bit_4_34 bit_4_35 R_bl
Rbb_4_34 bitb_4_34 bitb_4_35 R_bl
Cb_4_34 bit_4_34 gnd C_bl
Cbb_4_34 bitb_4_34 gnd C_bl
Rb_4_35 bit_4_35 bit_4_36 R_bl
Rbb_4_35 bitb_4_35 bitb_4_36 R_bl
Cb_4_35 bit_4_35 gnd C_bl
Cbb_4_35 bitb_4_35 gnd C_bl
Rb_4_36 bit_4_36 bit_4_37 R_bl
Rbb_4_36 bitb_4_36 bitb_4_37 R_bl
Cb_4_36 bit_4_36 gnd C_bl
Cbb_4_36 bitb_4_36 gnd C_bl
Rb_4_37 bit_4_37 bit_4_38 R_bl
Rbb_4_37 bitb_4_37 bitb_4_38 R_bl
Cb_4_37 bit_4_37 gnd C_bl
Cbb_4_37 bitb_4_37 gnd C_bl
Rb_4_38 bit_4_38 bit_4_39 R_bl
Rbb_4_38 bitb_4_38 bitb_4_39 R_bl
Cb_4_38 bit_4_38 gnd C_bl
Cbb_4_38 bitb_4_38 gnd C_bl
Rb_4_39 bit_4_39 bit_4_40 R_bl
Rbb_4_39 bitb_4_39 bitb_4_40 R_bl
Cb_4_39 bit_4_39 gnd C_bl
Cbb_4_39 bitb_4_39 gnd C_bl
Rb_4_40 bit_4_40 bit_4_41 R_bl
Rbb_4_40 bitb_4_40 bitb_4_41 R_bl
Cb_4_40 bit_4_40 gnd C_bl
Cbb_4_40 bitb_4_40 gnd C_bl
Rb_4_41 bit_4_41 bit_4_42 R_bl
Rbb_4_41 bitb_4_41 bitb_4_42 R_bl
Cb_4_41 bit_4_41 gnd C_bl
Cbb_4_41 bitb_4_41 gnd C_bl
Rb_4_42 bit_4_42 bit_4_43 R_bl
Rbb_4_42 bitb_4_42 bitb_4_43 R_bl
Cb_4_42 bit_4_42 gnd C_bl
Cbb_4_42 bitb_4_42 gnd C_bl
Rb_4_43 bit_4_43 bit_4_44 R_bl
Rbb_4_43 bitb_4_43 bitb_4_44 R_bl
Cb_4_43 bit_4_43 gnd C_bl
Cbb_4_43 bitb_4_43 gnd C_bl
Rb_4_44 bit_4_44 bit_4_45 R_bl
Rbb_4_44 bitb_4_44 bitb_4_45 R_bl
Cb_4_44 bit_4_44 gnd C_bl
Cbb_4_44 bitb_4_44 gnd C_bl
Rb_4_45 bit_4_45 bit_4_46 R_bl
Rbb_4_45 bitb_4_45 bitb_4_46 R_bl
Cb_4_45 bit_4_45 gnd C_bl
Cbb_4_45 bitb_4_45 gnd C_bl
Rb_4_46 bit_4_46 bit_4_47 R_bl
Rbb_4_46 bitb_4_46 bitb_4_47 R_bl
Cb_4_46 bit_4_46 gnd C_bl
Cbb_4_46 bitb_4_46 gnd C_bl
Rb_4_47 bit_4_47 bit_4_48 R_bl
Rbb_4_47 bitb_4_47 bitb_4_48 R_bl
Cb_4_47 bit_4_47 gnd C_bl
Cbb_4_47 bitb_4_47 gnd C_bl
Rb_4_48 bit_4_48 bit_4_49 R_bl
Rbb_4_48 bitb_4_48 bitb_4_49 R_bl
Cb_4_48 bit_4_48 gnd C_bl
Cbb_4_48 bitb_4_48 gnd C_bl
Rb_4_49 bit_4_49 bit_4_50 R_bl
Rbb_4_49 bitb_4_49 bitb_4_50 R_bl
Cb_4_49 bit_4_49 gnd C_bl
Cbb_4_49 bitb_4_49 gnd C_bl
Rb_4_50 bit_4_50 bit_4_51 R_bl
Rbb_4_50 bitb_4_50 bitb_4_51 R_bl
Cb_4_50 bit_4_50 gnd C_bl
Cbb_4_50 bitb_4_50 gnd C_bl
Rb_4_51 bit_4_51 bit_4_52 R_bl
Rbb_4_51 bitb_4_51 bitb_4_52 R_bl
Cb_4_51 bit_4_51 gnd C_bl
Cbb_4_51 bitb_4_51 gnd C_bl
Rb_4_52 bit_4_52 bit_4_53 R_bl
Rbb_4_52 bitb_4_52 bitb_4_53 R_bl
Cb_4_52 bit_4_52 gnd C_bl
Cbb_4_52 bitb_4_52 gnd C_bl
Rb_4_53 bit_4_53 bit_4_54 R_bl
Rbb_4_53 bitb_4_53 bitb_4_54 R_bl
Cb_4_53 bit_4_53 gnd C_bl
Cbb_4_53 bitb_4_53 gnd C_bl
Rb_4_54 bit_4_54 bit_4_55 R_bl
Rbb_4_54 bitb_4_54 bitb_4_55 R_bl
Cb_4_54 bit_4_54 gnd C_bl
Cbb_4_54 bitb_4_54 gnd C_bl
Rb_4_55 bit_4_55 bit_4_56 R_bl
Rbb_4_55 bitb_4_55 bitb_4_56 R_bl
Cb_4_55 bit_4_55 gnd C_bl
Cbb_4_55 bitb_4_55 gnd C_bl
Rb_4_56 bit_4_56 bit_4_57 R_bl
Rbb_4_56 bitb_4_56 bitb_4_57 R_bl
Cb_4_56 bit_4_56 gnd C_bl
Cbb_4_56 bitb_4_56 gnd C_bl
Rb_4_57 bit_4_57 bit_4_58 R_bl
Rbb_4_57 bitb_4_57 bitb_4_58 R_bl
Cb_4_57 bit_4_57 gnd C_bl
Cbb_4_57 bitb_4_57 gnd C_bl
Rb_4_58 bit_4_58 bit_4_59 R_bl
Rbb_4_58 bitb_4_58 bitb_4_59 R_bl
Cb_4_58 bit_4_58 gnd C_bl
Cbb_4_58 bitb_4_58 gnd C_bl
Rb_4_59 bit_4_59 bit_4_60 R_bl
Rbb_4_59 bitb_4_59 bitb_4_60 R_bl
Cb_4_59 bit_4_59 gnd C_bl
Cbb_4_59 bitb_4_59 gnd C_bl
Rb_4_60 bit_4_60 bit_4_61 R_bl
Rbb_4_60 bitb_4_60 bitb_4_61 R_bl
Cb_4_60 bit_4_60 gnd C_bl
Cbb_4_60 bitb_4_60 gnd C_bl
Rb_4_61 bit_4_61 bit_4_62 R_bl
Rbb_4_61 bitb_4_61 bitb_4_62 R_bl
Cb_4_61 bit_4_61 gnd C_bl
Cbb_4_61 bitb_4_61 gnd C_bl
Rb_4_62 bit_4_62 bit_4_63 R_bl
Rbb_4_62 bitb_4_62 bitb_4_63 R_bl
Cb_4_62 bit_4_62 gnd C_bl
Cbb_4_62 bitb_4_62 gnd C_bl
Rb_4_63 bit_4_63 bit_4_64 R_bl
Rbb_4_63 bitb_4_63 bitb_4_64 R_bl
Cb_4_63 bit_4_63 gnd C_bl
Cbb_4_63 bitb_4_63 gnd C_bl
Rb_4_64 bit_4_64 bit_4_65 R_bl
Rbb_4_64 bitb_4_64 bitb_4_65 R_bl
Cb_4_64 bit_4_64 gnd C_bl
Cbb_4_64 bitb_4_64 gnd C_bl
Rb_4_65 bit_4_65 bit_4_66 R_bl
Rbb_4_65 bitb_4_65 bitb_4_66 R_bl
Cb_4_65 bit_4_65 gnd C_bl
Cbb_4_65 bitb_4_65 gnd C_bl
Rb_4_66 bit_4_66 bit_4_67 R_bl
Rbb_4_66 bitb_4_66 bitb_4_67 R_bl
Cb_4_66 bit_4_66 gnd C_bl
Cbb_4_66 bitb_4_66 gnd C_bl
Rb_4_67 bit_4_67 bit_4_68 R_bl
Rbb_4_67 bitb_4_67 bitb_4_68 R_bl
Cb_4_67 bit_4_67 gnd C_bl
Cbb_4_67 bitb_4_67 gnd C_bl
Rb_4_68 bit_4_68 bit_4_69 R_bl
Rbb_4_68 bitb_4_68 bitb_4_69 R_bl
Cb_4_68 bit_4_68 gnd C_bl
Cbb_4_68 bitb_4_68 gnd C_bl
Rb_4_69 bit_4_69 bit_4_70 R_bl
Rbb_4_69 bitb_4_69 bitb_4_70 R_bl
Cb_4_69 bit_4_69 gnd C_bl
Cbb_4_69 bitb_4_69 gnd C_bl
Rb_4_70 bit_4_70 bit_4_71 R_bl
Rbb_4_70 bitb_4_70 bitb_4_71 R_bl
Cb_4_70 bit_4_70 gnd C_bl
Cbb_4_70 bitb_4_70 gnd C_bl
Rb_4_71 bit_4_71 bit_4_72 R_bl
Rbb_4_71 bitb_4_71 bitb_4_72 R_bl
Cb_4_71 bit_4_71 gnd C_bl
Cbb_4_71 bitb_4_71 gnd C_bl
Rb_4_72 bit_4_72 bit_4_73 R_bl
Rbb_4_72 bitb_4_72 bitb_4_73 R_bl
Cb_4_72 bit_4_72 gnd C_bl
Cbb_4_72 bitb_4_72 gnd C_bl
Rb_4_73 bit_4_73 bit_4_74 R_bl
Rbb_4_73 bitb_4_73 bitb_4_74 R_bl
Cb_4_73 bit_4_73 gnd C_bl
Cbb_4_73 bitb_4_73 gnd C_bl
Rb_4_74 bit_4_74 bit_4_75 R_bl
Rbb_4_74 bitb_4_74 bitb_4_75 R_bl
Cb_4_74 bit_4_74 gnd C_bl
Cbb_4_74 bitb_4_74 gnd C_bl
Rb_4_75 bit_4_75 bit_4_76 R_bl
Rbb_4_75 bitb_4_75 bitb_4_76 R_bl
Cb_4_75 bit_4_75 gnd C_bl
Cbb_4_75 bitb_4_75 gnd C_bl
Rb_4_76 bit_4_76 bit_4_77 R_bl
Rbb_4_76 bitb_4_76 bitb_4_77 R_bl
Cb_4_76 bit_4_76 gnd C_bl
Cbb_4_76 bitb_4_76 gnd C_bl
Rb_4_77 bit_4_77 bit_4_78 R_bl
Rbb_4_77 bitb_4_77 bitb_4_78 R_bl
Cb_4_77 bit_4_77 gnd C_bl
Cbb_4_77 bitb_4_77 gnd C_bl
Rb_4_78 bit_4_78 bit_4_79 R_bl
Rbb_4_78 bitb_4_78 bitb_4_79 R_bl
Cb_4_78 bit_4_78 gnd C_bl
Cbb_4_78 bitb_4_78 gnd C_bl
Rb_4_79 bit_4_79 bit_4_80 R_bl
Rbb_4_79 bitb_4_79 bitb_4_80 R_bl
Cb_4_79 bit_4_79 gnd C_bl
Cbb_4_79 bitb_4_79 gnd C_bl
Rb_4_80 bit_4_80 bit_4_81 R_bl
Rbb_4_80 bitb_4_80 bitb_4_81 R_bl
Cb_4_80 bit_4_80 gnd C_bl
Cbb_4_80 bitb_4_80 gnd C_bl
Rb_4_81 bit_4_81 bit_4_82 R_bl
Rbb_4_81 bitb_4_81 bitb_4_82 R_bl
Cb_4_81 bit_4_81 gnd C_bl
Cbb_4_81 bitb_4_81 gnd C_bl
Rb_4_82 bit_4_82 bit_4_83 R_bl
Rbb_4_82 bitb_4_82 bitb_4_83 R_bl
Cb_4_82 bit_4_82 gnd C_bl
Cbb_4_82 bitb_4_82 gnd C_bl
Rb_4_83 bit_4_83 bit_4_84 R_bl
Rbb_4_83 bitb_4_83 bitb_4_84 R_bl
Cb_4_83 bit_4_83 gnd C_bl
Cbb_4_83 bitb_4_83 gnd C_bl
Rb_4_84 bit_4_84 bit_4_85 R_bl
Rbb_4_84 bitb_4_84 bitb_4_85 R_bl
Cb_4_84 bit_4_84 gnd C_bl
Cbb_4_84 bitb_4_84 gnd C_bl
Rb_4_85 bit_4_85 bit_4_86 R_bl
Rbb_4_85 bitb_4_85 bitb_4_86 R_bl
Cb_4_85 bit_4_85 gnd C_bl
Cbb_4_85 bitb_4_85 gnd C_bl
Rb_4_86 bit_4_86 bit_4_87 R_bl
Rbb_4_86 bitb_4_86 bitb_4_87 R_bl
Cb_4_86 bit_4_86 gnd C_bl
Cbb_4_86 bitb_4_86 gnd C_bl
Rb_4_87 bit_4_87 bit_4_88 R_bl
Rbb_4_87 bitb_4_87 bitb_4_88 R_bl
Cb_4_87 bit_4_87 gnd C_bl
Cbb_4_87 bitb_4_87 gnd C_bl
Rb_4_88 bit_4_88 bit_4_89 R_bl
Rbb_4_88 bitb_4_88 bitb_4_89 R_bl
Cb_4_88 bit_4_88 gnd C_bl
Cbb_4_88 bitb_4_88 gnd C_bl
Rb_4_89 bit_4_89 bit_4_90 R_bl
Rbb_4_89 bitb_4_89 bitb_4_90 R_bl
Cb_4_89 bit_4_89 gnd C_bl
Cbb_4_89 bitb_4_89 gnd C_bl
Rb_4_90 bit_4_90 bit_4_91 R_bl
Rbb_4_90 bitb_4_90 bitb_4_91 R_bl
Cb_4_90 bit_4_90 gnd C_bl
Cbb_4_90 bitb_4_90 gnd C_bl
Rb_4_91 bit_4_91 bit_4_92 R_bl
Rbb_4_91 bitb_4_91 bitb_4_92 R_bl
Cb_4_91 bit_4_91 gnd C_bl
Cbb_4_91 bitb_4_91 gnd C_bl
Rb_4_92 bit_4_92 bit_4_93 R_bl
Rbb_4_92 bitb_4_92 bitb_4_93 R_bl
Cb_4_92 bit_4_92 gnd C_bl
Cbb_4_92 bitb_4_92 gnd C_bl
Rb_4_93 bit_4_93 bit_4_94 R_bl
Rbb_4_93 bitb_4_93 bitb_4_94 R_bl
Cb_4_93 bit_4_93 gnd C_bl
Cbb_4_93 bitb_4_93 gnd C_bl
Rb_4_94 bit_4_94 bit_4_95 R_bl
Rbb_4_94 bitb_4_94 bitb_4_95 R_bl
Cb_4_94 bit_4_94 gnd C_bl
Cbb_4_94 bitb_4_94 gnd C_bl
Rb_4_95 bit_4_95 bit_4_96 R_bl
Rbb_4_95 bitb_4_95 bitb_4_96 R_bl
Cb_4_95 bit_4_95 gnd C_bl
Cbb_4_95 bitb_4_95 gnd C_bl
Rb_4_96 bit_4_96 bit_4_97 R_bl
Rbb_4_96 bitb_4_96 bitb_4_97 R_bl
Cb_4_96 bit_4_96 gnd C_bl
Cbb_4_96 bitb_4_96 gnd C_bl
Rb_4_97 bit_4_97 bit_4_98 R_bl
Rbb_4_97 bitb_4_97 bitb_4_98 R_bl
Cb_4_97 bit_4_97 gnd C_bl
Cbb_4_97 bitb_4_97 gnd C_bl
Rb_4_98 bit_4_98 bit_4_99 R_bl
Rbb_4_98 bitb_4_98 bitb_4_99 R_bl
Cb_4_98 bit_4_98 gnd C_bl
Cbb_4_98 bitb_4_98 gnd C_bl
Rb_4_99 bit_4_99 bit_4_100 R_bl
Rbb_4_99 bitb_4_99 bitb_4_100 R_bl
Cb_4_99 bit_4_99 gnd C_bl
Cbb_4_99 bitb_4_99 gnd C_bl
Rb_5_0 bit_5_0 bit_5_1 R_bl
Rbb_5_0 bitb_5_0 bitb_5_1 R_bl
Cb_5_0 bit_5_0 gnd C_bl
Cbb_5_0 bitb_5_0 gnd C_bl
Rb_5_1 bit_5_1 bit_5_2 R_bl
Rbb_5_1 bitb_5_1 bitb_5_2 R_bl
Cb_5_1 bit_5_1 gnd C_bl
Cbb_5_1 bitb_5_1 gnd C_bl
Rb_5_2 bit_5_2 bit_5_3 R_bl
Rbb_5_2 bitb_5_2 bitb_5_3 R_bl
Cb_5_2 bit_5_2 gnd C_bl
Cbb_5_2 bitb_5_2 gnd C_bl
Rb_5_3 bit_5_3 bit_5_4 R_bl
Rbb_5_3 bitb_5_3 bitb_5_4 R_bl
Cb_5_3 bit_5_3 gnd C_bl
Cbb_5_3 bitb_5_3 gnd C_bl
Rb_5_4 bit_5_4 bit_5_5 R_bl
Rbb_5_4 bitb_5_4 bitb_5_5 R_bl
Cb_5_4 bit_5_4 gnd C_bl
Cbb_5_4 bitb_5_4 gnd C_bl
Rb_5_5 bit_5_5 bit_5_6 R_bl
Rbb_5_5 bitb_5_5 bitb_5_6 R_bl
Cb_5_5 bit_5_5 gnd C_bl
Cbb_5_5 bitb_5_5 gnd C_bl
Rb_5_6 bit_5_6 bit_5_7 R_bl
Rbb_5_6 bitb_5_6 bitb_5_7 R_bl
Cb_5_6 bit_5_6 gnd C_bl
Cbb_5_6 bitb_5_6 gnd C_bl
Rb_5_7 bit_5_7 bit_5_8 R_bl
Rbb_5_7 bitb_5_7 bitb_5_8 R_bl
Cb_5_7 bit_5_7 gnd C_bl
Cbb_5_7 bitb_5_7 gnd C_bl
Rb_5_8 bit_5_8 bit_5_9 R_bl
Rbb_5_8 bitb_5_8 bitb_5_9 R_bl
Cb_5_8 bit_5_8 gnd C_bl
Cbb_5_8 bitb_5_8 gnd C_bl
Rb_5_9 bit_5_9 bit_5_10 R_bl
Rbb_5_9 bitb_5_9 bitb_5_10 R_bl
Cb_5_9 bit_5_9 gnd C_bl
Cbb_5_9 bitb_5_9 gnd C_bl
Rb_5_10 bit_5_10 bit_5_11 R_bl
Rbb_5_10 bitb_5_10 bitb_5_11 R_bl
Cb_5_10 bit_5_10 gnd C_bl
Cbb_5_10 bitb_5_10 gnd C_bl
Rb_5_11 bit_5_11 bit_5_12 R_bl
Rbb_5_11 bitb_5_11 bitb_5_12 R_bl
Cb_5_11 bit_5_11 gnd C_bl
Cbb_5_11 bitb_5_11 gnd C_bl
Rb_5_12 bit_5_12 bit_5_13 R_bl
Rbb_5_12 bitb_5_12 bitb_5_13 R_bl
Cb_5_12 bit_5_12 gnd C_bl
Cbb_5_12 bitb_5_12 gnd C_bl
Rb_5_13 bit_5_13 bit_5_14 R_bl
Rbb_5_13 bitb_5_13 bitb_5_14 R_bl
Cb_5_13 bit_5_13 gnd C_bl
Cbb_5_13 bitb_5_13 gnd C_bl
Rb_5_14 bit_5_14 bit_5_15 R_bl
Rbb_5_14 bitb_5_14 bitb_5_15 R_bl
Cb_5_14 bit_5_14 gnd C_bl
Cbb_5_14 bitb_5_14 gnd C_bl
Rb_5_15 bit_5_15 bit_5_16 R_bl
Rbb_5_15 bitb_5_15 bitb_5_16 R_bl
Cb_5_15 bit_5_15 gnd C_bl
Cbb_5_15 bitb_5_15 gnd C_bl
Rb_5_16 bit_5_16 bit_5_17 R_bl
Rbb_5_16 bitb_5_16 bitb_5_17 R_bl
Cb_5_16 bit_5_16 gnd C_bl
Cbb_5_16 bitb_5_16 gnd C_bl
Rb_5_17 bit_5_17 bit_5_18 R_bl
Rbb_5_17 bitb_5_17 bitb_5_18 R_bl
Cb_5_17 bit_5_17 gnd C_bl
Cbb_5_17 bitb_5_17 gnd C_bl
Rb_5_18 bit_5_18 bit_5_19 R_bl
Rbb_5_18 bitb_5_18 bitb_5_19 R_bl
Cb_5_18 bit_5_18 gnd C_bl
Cbb_5_18 bitb_5_18 gnd C_bl
Rb_5_19 bit_5_19 bit_5_20 R_bl
Rbb_5_19 bitb_5_19 bitb_5_20 R_bl
Cb_5_19 bit_5_19 gnd C_bl
Cbb_5_19 bitb_5_19 gnd C_bl
Rb_5_20 bit_5_20 bit_5_21 R_bl
Rbb_5_20 bitb_5_20 bitb_5_21 R_bl
Cb_5_20 bit_5_20 gnd C_bl
Cbb_5_20 bitb_5_20 gnd C_bl
Rb_5_21 bit_5_21 bit_5_22 R_bl
Rbb_5_21 bitb_5_21 bitb_5_22 R_bl
Cb_5_21 bit_5_21 gnd C_bl
Cbb_5_21 bitb_5_21 gnd C_bl
Rb_5_22 bit_5_22 bit_5_23 R_bl
Rbb_5_22 bitb_5_22 bitb_5_23 R_bl
Cb_5_22 bit_5_22 gnd C_bl
Cbb_5_22 bitb_5_22 gnd C_bl
Rb_5_23 bit_5_23 bit_5_24 R_bl
Rbb_5_23 bitb_5_23 bitb_5_24 R_bl
Cb_5_23 bit_5_23 gnd C_bl
Cbb_5_23 bitb_5_23 gnd C_bl
Rb_5_24 bit_5_24 bit_5_25 R_bl
Rbb_5_24 bitb_5_24 bitb_5_25 R_bl
Cb_5_24 bit_5_24 gnd C_bl
Cbb_5_24 bitb_5_24 gnd C_bl
Rb_5_25 bit_5_25 bit_5_26 R_bl
Rbb_5_25 bitb_5_25 bitb_5_26 R_bl
Cb_5_25 bit_5_25 gnd C_bl
Cbb_5_25 bitb_5_25 gnd C_bl
Rb_5_26 bit_5_26 bit_5_27 R_bl
Rbb_5_26 bitb_5_26 bitb_5_27 R_bl
Cb_5_26 bit_5_26 gnd C_bl
Cbb_5_26 bitb_5_26 gnd C_bl
Rb_5_27 bit_5_27 bit_5_28 R_bl
Rbb_5_27 bitb_5_27 bitb_5_28 R_bl
Cb_5_27 bit_5_27 gnd C_bl
Cbb_5_27 bitb_5_27 gnd C_bl
Rb_5_28 bit_5_28 bit_5_29 R_bl
Rbb_5_28 bitb_5_28 bitb_5_29 R_bl
Cb_5_28 bit_5_28 gnd C_bl
Cbb_5_28 bitb_5_28 gnd C_bl
Rb_5_29 bit_5_29 bit_5_30 R_bl
Rbb_5_29 bitb_5_29 bitb_5_30 R_bl
Cb_5_29 bit_5_29 gnd C_bl
Cbb_5_29 bitb_5_29 gnd C_bl
Rb_5_30 bit_5_30 bit_5_31 R_bl
Rbb_5_30 bitb_5_30 bitb_5_31 R_bl
Cb_5_30 bit_5_30 gnd C_bl
Cbb_5_30 bitb_5_30 gnd C_bl
Rb_5_31 bit_5_31 bit_5_32 R_bl
Rbb_5_31 bitb_5_31 bitb_5_32 R_bl
Cb_5_31 bit_5_31 gnd C_bl
Cbb_5_31 bitb_5_31 gnd C_bl
Rb_5_32 bit_5_32 bit_5_33 R_bl
Rbb_5_32 bitb_5_32 bitb_5_33 R_bl
Cb_5_32 bit_5_32 gnd C_bl
Cbb_5_32 bitb_5_32 gnd C_bl
Rb_5_33 bit_5_33 bit_5_34 R_bl
Rbb_5_33 bitb_5_33 bitb_5_34 R_bl
Cb_5_33 bit_5_33 gnd C_bl
Cbb_5_33 bitb_5_33 gnd C_bl
Rb_5_34 bit_5_34 bit_5_35 R_bl
Rbb_5_34 bitb_5_34 bitb_5_35 R_bl
Cb_5_34 bit_5_34 gnd C_bl
Cbb_5_34 bitb_5_34 gnd C_bl
Rb_5_35 bit_5_35 bit_5_36 R_bl
Rbb_5_35 bitb_5_35 bitb_5_36 R_bl
Cb_5_35 bit_5_35 gnd C_bl
Cbb_5_35 bitb_5_35 gnd C_bl
Rb_5_36 bit_5_36 bit_5_37 R_bl
Rbb_5_36 bitb_5_36 bitb_5_37 R_bl
Cb_5_36 bit_5_36 gnd C_bl
Cbb_5_36 bitb_5_36 gnd C_bl
Rb_5_37 bit_5_37 bit_5_38 R_bl
Rbb_5_37 bitb_5_37 bitb_5_38 R_bl
Cb_5_37 bit_5_37 gnd C_bl
Cbb_5_37 bitb_5_37 gnd C_bl
Rb_5_38 bit_5_38 bit_5_39 R_bl
Rbb_5_38 bitb_5_38 bitb_5_39 R_bl
Cb_5_38 bit_5_38 gnd C_bl
Cbb_5_38 bitb_5_38 gnd C_bl
Rb_5_39 bit_5_39 bit_5_40 R_bl
Rbb_5_39 bitb_5_39 bitb_5_40 R_bl
Cb_5_39 bit_5_39 gnd C_bl
Cbb_5_39 bitb_5_39 gnd C_bl
Rb_5_40 bit_5_40 bit_5_41 R_bl
Rbb_5_40 bitb_5_40 bitb_5_41 R_bl
Cb_5_40 bit_5_40 gnd C_bl
Cbb_5_40 bitb_5_40 gnd C_bl
Rb_5_41 bit_5_41 bit_5_42 R_bl
Rbb_5_41 bitb_5_41 bitb_5_42 R_bl
Cb_5_41 bit_5_41 gnd C_bl
Cbb_5_41 bitb_5_41 gnd C_bl
Rb_5_42 bit_5_42 bit_5_43 R_bl
Rbb_5_42 bitb_5_42 bitb_5_43 R_bl
Cb_5_42 bit_5_42 gnd C_bl
Cbb_5_42 bitb_5_42 gnd C_bl
Rb_5_43 bit_5_43 bit_5_44 R_bl
Rbb_5_43 bitb_5_43 bitb_5_44 R_bl
Cb_5_43 bit_5_43 gnd C_bl
Cbb_5_43 bitb_5_43 gnd C_bl
Rb_5_44 bit_5_44 bit_5_45 R_bl
Rbb_5_44 bitb_5_44 bitb_5_45 R_bl
Cb_5_44 bit_5_44 gnd C_bl
Cbb_5_44 bitb_5_44 gnd C_bl
Rb_5_45 bit_5_45 bit_5_46 R_bl
Rbb_5_45 bitb_5_45 bitb_5_46 R_bl
Cb_5_45 bit_5_45 gnd C_bl
Cbb_5_45 bitb_5_45 gnd C_bl
Rb_5_46 bit_5_46 bit_5_47 R_bl
Rbb_5_46 bitb_5_46 bitb_5_47 R_bl
Cb_5_46 bit_5_46 gnd C_bl
Cbb_5_46 bitb_5_46 gnd C_bl
Rb_5_47 bit_5_47 bit_5_48 R_bl
Rbb_5_47 bitb_5_47 bitb_5_48 R_bl
Cb_5_47 bit_5_47 gnd C_bl
Cbb_5_47 bitb_5_47 gnd C_bl
Rb_5_48 bit_5_48 bit_5_49 R_bl
Rbb_5_48 bitb_5_48 bitb_5_49 R_bl
Cb_5_48 bit_5_48 gnd C_bl
Cbb_5_48 bitb_5_48 gnd C_bl
Rb_5_49 bit_5_49 bit_5_50 R_bl
Rbb_5_49 bitb_5_49 bitb_5_50 R_bl
Cb_5_49 bit_5_49 gnd C_bl
Cbb_5_49 bitb_5_49 gnd C_bl
Rb_5_50 bit_5_50 bit_5_51 R_bl
Rbb_5_50 bitb_5_50 bitb_5_51 R_bl
Cb_5_50 bit_5_50 gnd C_bl
Cbb_5_50 bitb_5_50 gnd C_bl
Rb_5_51 bit_5_51 bit_5_52 R_bl
Rbb_5_51 bitb_5_51 bitb_5_52 R_bl
Cb_5_51 bit_5_51 gnd C_bl
Cbb_5_51 bitb_5_51 gnd C_bl
Rb_5_52 bit_5_52 bit_5_53 R_bl
Rbb_5_52 bitb_5_52 bitb_5_53 R_bl
Cb_5_52 bit_5_52 gnd C_bl
Cbb_5_52 bitb_5_52 gnd C_bl
Rb_5_53 bit_5_53 bit_5_54 R_bl
Rbb_5_53 bitb_5_53 bitb_5_54 R_bl
Cb_5_53 bit_5_53 gnd C_bl
Cbb_5_53 bitb_5_53 gnd C_bl
Rb_5_54 bit_5_54 bit_5_55 R_bl
Rbb_5_54 bitb_5_54 bitb_5_55 R_bl
Cb_5_54 bit_5_54 gnd C_bl
Cbb_5_54 bitb_5_54 gnd C_bl
Rb_5_55 bit_5_55 bit_5_56 R_bl
Rbb_5_55 bitb_5_55 bitb_5_56 R_bl
Cb_5_55 bit_5_55 gnd C_bl
Cbb_5_55 bitb_5_55 gnd C_bl
Rb_5_56 bit_5_56 bit_5_57 R_bl
Rbb_5_56 bitb_5_56 bitb_5_57 R_bl
Cb_5_56 bit_5_56 gnd C_bl
Cbb_5_56 bitb_5_56 gnd C_bl
Rb_5_57 bit_5_57 bit_5_58 R_bl
Rbb_5_57 bitb_5_57 bitb_5_58 R_bl
Cb_5_57 bit_5_57 gnd C_bl
Cbb_5_57 bitb_5_57 gnd C_bl
Rb_5_58 bit_5_58 bit_5_59 R_bl
Rbb_5_58 bitb_5_58 bitb_5_59 R_bl
Cb_5_58 bit_5_58 gnd C_bl
Cbb_5_58 bitb_5_58 gnd C_bl
Rb_5_59 bit_5_59 bit_5_60 R_bl
Rbb_5_59 bitb_5_59 bitb_5_60 R_bl
Cb_5_59 bit_5_59 gnd C_bl
Cbb_5_59 bitb_5_59 gnd C_bl
Rb_5_60 bit_5_60 bit_5_61 R_bl
Rbb_5_60 bitb_5_60 bitb_5_61 R_bl
Cb_5_60 bit_5_60 gnd C_bl
Cbb_5_60 bitb_5_60 gnd C_bl
Rb_5_61 bit_5_61 bit_5_62 R_bl
Rbb_5_61 bitb_5_61 bitb_5_62 R_bl
Cb_5_61 bit_5_61 gnd C_bl
Cbb_5_61 bitb_5_61 gnd C_bl
Rb_5_62 bit_5_62 bit_5_63 R_bl
Rbb_5_62 bitb_5_62 bitb_5_63 R_bl
Cb_5_62 bit_5_62 gnd C_bl
Cbb_5_62 bitb_5_62 gnd C_bl
Rb_5_63 bit_5_63 bit_5_64 R_bl
Rbb_5_63 bitb_5_63 bitb_5_64 R_bl
Cb_5_63 bit_5_63 gnd C_bl
Cbb_5_63 bitb_5_63 gnd C_bl
Rb_5_64 bit_5_64 bit_5_65 R_bl
Rbb_5_64 bitb_5_64 bitb_5_65 R_bl
Cb_5_64 bit_5_64 gnd C_bl
Cbb_5_64 bitb_5_64 gnd C_bl
Rb_5_65 bit_5_65 bit_5_66 R_bl
Rbb_5_65 bitb_5_65 bitb_5_66 R_bl
Cb_5_65 bit_5_65 gnd C_bl
Cbb_5_65 bitb_5_65 gnd C_bl
Rb_5_66 bit_5_66 bit_5_67 R_bl
Rbb_5_66 bitb_5_66 bitb_5_67 R_bl
Cb_5_66 bit_5_66 gnd C_bl
Cbb_5_66 bitb_5_66 gnd C_bl
Rb_5_67 bit_5_67 bit_5_68 R_bl
Rbb_5_67 bitb_5_67 bitb_5_68 R_bl
Cb_5_67 bit_5_67 gnd C_bl
Cbb_5_67 bitb_5_67 gnd C_bl
Rb_5_68 bit_5_68 bit_5_69 R_bl
Rbb_5_68 bitb_5_68 bitb_5_69 R_bl
Cb_5_68 bit_5_68 gnd C_bl
Cbb_5_68 bitb_5_68 gnd C_bl
Rb_5_69 bit_5_69 bit_5_70 R_bl
Rbb_5_69 bitb_5_69 bitb_5_70 R_bl
Cb_5_69 bit_5_69 gnd C_bl
Cbb_5_69 bitb_5_69 gnd C_bl
Rb_5_70 bit_5_70 bit_5_71 R_bl
Rbb_5_70 bitb_5_70 bitb_5_71 R_bl
Cb_5_70 bit_5_70 gnd C_bl
Cbb_5_70 bitb_5_70 gnd C_bl
Rb_5_71 bit_5_71 bit_5_72 R_bl
Rbb_5_71 bitb_5_71 bitb_5_72 R_bl
Cb_5_71 bit_5_71 gnd C_bl
Cbb_5_71 bitb_5_71 gnd C_bl
Rb_5_72 bit_5_72 bit_5_73 R_bl
Rbb_5_72 bitb_5_72 bitb_5_73 R_bl
Cb_5_72 bit_5_72 gnd C_bl
Cbb_5_72 bitb_5_72 gnd C_bl
Rb_5_73 bit_5_73 bit_5_74 R_bl
Rbb_5_73 bitb_5_73 bitb_5_74 R_bl
Cb_5_73 bit_5_73 gnd C_bl
Cbb_5_73 bitb_5_73 gnd C_bl
Rb_5_74 bit_5_74 bit_5_75 R_bl
Rbb_5_74 bitb_5_74 bitb_5_75 R_bl
Cb_5_74 bit_5_74 gnd C_bl
Cbb_5_74 bitb_5_74 gnd C_bl
Rb_5_75 bit_5_75 bit_5_76 R_bl
Rbb_5_75 bitb_5_75 bitb_5_76 R_bl
Cb_5_75 bit_5_75 gnd C_bl
Cbb_5_75 bitb_5_75 gnd C_bl
Rb_5_76 bit_5_76 bit_5_77 R_bl
Rbb_5_76 bitb_5_76 bitb_5_77 R_bl
Cb_5_76 bit_5_76 gnd C_bl
Cbb_5_76 bitb_5_76 gnd C_bl
Rb_5_77 bit_5_77 bit_5_78 R_bl
Rbb_5_77 bitb_5_77 bitb_5_78 R_bl
Cb_5_77 bit_5_77 gnd C_bl
Cbb_5_77 bitb_5_77 gnd C_bl
Rb_5_78 bit_5_78 bit_5_79 R_bl
Rbb_5_78 bitb_5_78 bitb_5_79 R_bl
Cb_5_78 bit_5_78 gnd C_bl
Cbb_5_78 bitb_5_78 gnd C_bl
Rb_5_79 bit_5_79 bit_5_80 R_bl
Rbb_5_79 bitb_5_79 bitb_5_80 R_bl
Cb_5_79 bit_5_79 gnd C_bl
Cbb_5_79 bitb_5_79 gnd C_bl
Rb_5_80 bit_5_80 bit_5_81 R_bl
Rbb_5_80 bitb_5_80 bitb_5_81 R_bl
Cb_5_80 bit_5_80 gnd C_bl
Cbb_5_80 bitb_5_80 gnd C_bl
Rb_5_81 bit_5_81 bit_5_82 R_bl
Rbb_5_81 bitb_5_81 bitb_5_82 R_bl
Cb_5_81 bit_5_81 gnd C_bl
Cbb_5_81 bitb_5_81 gnd C_bl
Rb_5_82 bit_5_82 bit_5_83 R_bl
Rbb_5_82 bitb_5_82 bitb_5_83 R_bl
Cb_5_82 bit_5_82 gnd C_bl
Cbb_5_82 bitb_5_82 gnd C_bl
Rb_5_83 bit_5_83 bit_5_84 R_bl
Rbb_5_83 bitb_5_83 bitb_5_84 R_bl
Cb_5_83 bit_5_83 gnd C_bl
Cbb_5_83 bitb_5_83 gnd C_bl
Rb_5_84 bit_5_84 bit_5_85 R_bl
Rbb_5_84 bitb_5_84 bitb_5_85 R_bl
Cb_5_84 bit_5_84 gnd C_bl
Cbb_5_84 bitb_5_84 gnd C_bl
Rb_5_85 bit_5_85 bit_5_86 R_bl
Rbb_5_85 bitb_5_85 bitb_5_86 R_bl
Cb_5_85 bit_5_85 gnd C_bl
Cbb_5_85 bitb_5_85 gnd C_bl
Rb_5_86 bit_5_86 bit_5_87 R_bl
Rbb_5_86 bitb_5_86 bitb_5_87 R_bl
Cb_5_86 bit_5_86 gnd C_bl
Cbb_5_86 bitb_5_86 gnd C_bl
Rb_5_87 bit_5_87 bit_5_88 R_bl
Rbb_5_87 bitb_5_87 bitb_5_88 R_bl
Cb_5_87 bit_5_87 gnd C_bl
Cbb_5_87 bitb_5_87 gnd C_bl
Rb_5_88 bit_5_88 bit_5_89 R_bl
Rbb_5_88 bitb_5_88 bitb_5_89 R_bl
Cb_5_88 bit_5_88 gnd C_bl
Cbb_5_88 bitb_5_88 gnd C_bl
Rb_5_89 bit_5_89 bit_5_90 R_bl
Rbb_5_89 bitb_5_89 bitb_5_90 R_bl
Cb_5_89 bit_5_89 gnd C_bl
Cbb_5_89 bitb_5_89 gnd C_bl
Rb_5_90 bit_5_90 bit_5_91 R_bl
Rbb_5_90 bitb_5_90 bitb_5_91 R_bl
Cb_5_90 bit_5_90 gnd C_bl
Cbb_5_90 bitb_5_90 gnd C_bl
Rb_5_91 bit_5_91 bit_5_92 R_bl
Rbb_5_91 bitb_5_91 bitb_5_92 R_bl
Cb_5_91 bit_5_91 gnd C_bl
Cbb_5_91 bitb_5_91 gnd C_bl
Rb_5_92 bit_5_92 bit_5_93 R_bl
Rbb_5_92 bitb_5_92 bitb_5_93 R_bl
Cb_5_92 bit_5_92 gnd C_bl
Cbb_5_92 bitb_5_92 gnd C_bl
Rb_5_93 bit_5_93 bit_5_94 R_bl
Rbb_5_93 bitb_5_93 bitb_5_94 R_bl
Cb_5_93 bit_5_93 gnd C_bl
Cbb_5_93 bitb_5_93 gnd C_bl
Rb_5_94 bit_5_94 bit_5_95 R_bl
Rbb_5_94 bitb_5_94 bitb_5_95 R_bl
Cb_5_94 bit_5_94 gnd C_bl
Cbb_5_94 bitb_5_94 gnd C_bl
Rb_5_95 bit_5_95 bit_5_96 R_bl
Rbb_5_95 bitb_5_95 bitb_5_96 R_bl
Cb_5_95 bit_5_95 gnd C_bl
Cbb_5_95 bitb_5_95 gnd C_bl
Rb_5_96 bit_5_96 bit_5_97 R_bl
Rbb_5_96 bitb_5_96 bitb_5_97 R_bl
Cb_5_96 bit_5_96 gnd C_bl
Cbb_5_96 bitb_5_96 gnd C_bl
Rb_5_97 bit_5_97 bit_5_98 R_bl
Rbb_5_97 bitb_5_97 bitb_5_98 R_bl
Cb_5_97 bit_5_97 gnd C_bl
Cbb_5_97 bitb_5_97 gnd C_bl
Rb_5_98 bit_5_98 bit_5_99 R_bl
Rbb_5_98 bitb_5_98 bitb_5_99 R_bl
Cb_5_98 bit_5_98 gnd C_bl
Cbb_5_98 bitb_5_98 gnd C_bl
Rb_5_99 bit_5_99 bit_5_100 R_bl
Rbb_5_99 bitb_5_99 bitb_5_100 R_bl
Cb_5_99 bit_5_99 gnd C_bl
Cbb_5_99 bitb_5_99 gnd C_bl
Rb_6_0 bit_6_0 bit_6_1 R_bl
Rbb_6_0 bitb_6_0 bitb_6_1 R_bl
Cb_6_0 bit_6_0 gnd C_bl
Cbb_6_0 bitb_6_0 gnd C_bl
Rb_6_1 bit_6_1 bit_6_2 R_bl
Rbb_6_1 bitb_6_1 bitb_6_2 R_bl
Cb_6_1 bit_6_1 gnd C_bl
Cbb_6_1 bitb_6_1 gnd C_bl
Rb_6_2 bit_6_2 bit_6_3 R_bl
Rbb_6_2 bitb_6_2 bitb_6_3 R_bl
Cb_6_2 bit_6_2 gnd C_bl
Cbb_6_2 bitb_6_2 gnd C_bl
Rb_6_3 bit_6_3 bit_6_4 R_bl
Rbb_6_3 bitb_6_3 bitb_6_4 R_bl
Cb_6_3 bit_6_3 gnd C_bl
Cbb_6_3 bitb_6_3 gnd C_bl
Rb_6_4 bit_6_4 bit_6_5 R_bl
Rbb_6_4 bitb_6_4 bitb_6_5 R_bl
Cb_6_4 bit_6_4 gnd C_bl
Cbb_6_4 bitb_6_4 gnd C_bl
Rb_6_5 bit_6_5 bit_6_6 R_bl
Rbb_6_5 bitb_6_5 bitb_6_6 R_bl
Cb_6_5 bit_6_5 gnd C_bl
Cbb_6_5 bitb_6_5 gnd C_bl
Rb_6_6 bit_6_6 bit_6_7 R_bl
Rbb_6_6 bitb_6_6 bitb_6_7 R_bl
Cb_6_6 bit_6_6 gnd C_bl
Cbb_6_6 bitb_6_6 gnd C_bl
Rb_6_7 bit_6_7 bit_6_8 R_bl
Rbb_6_7 bitb_6_7 bitb_6_8 R_bl
Cb_6_7 bit_6_7 gnd C_bl
Cbb_6_7 bitb_6_7 gnd C_bl
Rb_6_8 bit_6_8 bit_6_9 R_bl
Rbb_6_8 bitb_6_8 bitb_6_9 R_bl
Cb_6_8 bit_6_8 gnd C_bl
Cbb_6_8 bitb_6_8 gnd C_bl
Rb_6_9 bit_6_9 bit_6_10 R_bl
Rbb_6_9 bitb_6_9 bitb_6_10 R_bl
Cb_6_9 bit_6_9 gnd C_bl
Cbb_6_9 bitb_6_9 gnd C_bl
Rb_6_10 bit_6_10 bit_6_11 R_bl
Rbb_6_10 bitb_6_10 bitb_6_11 R_bl
Cb_6_10 bit_6_10 gnd C_bl
Cbb_6_10 bitb_6_10 gnd C_bl
Rb_6_11 bit_6_11 bit_6_12 R_bl
Rbb_6_11 bitb_6_11 bitb_6_12 R_bl
Cb_6_11 bit_6_11 gnd C_bl
Cbb_6_11 bitb_6_11 gnd C_bl
Rb_6_12 bit_6_12 bit_6_13 R_bl
Rbb_6_12 bitb_6_12 bitb_6_13 R_bl
Cb_6_12 bit_6_12 gnd C_bl
Cbb_6_12 bitb_6_12 gnd C_bl
Rb_6_13 bit_6_13 bit_6_14 R_bl
Rbb_6_13 bitb_6_13 bitb_6_14 R_bl
Cb_6_13 bit_6_13 gnd C_bl
Cbb_6_13 bitb_6_13 gnd C_bl
Rb_6_14 bit_6_14 bit_6_15 R_bl
Rbb_6_14 bitb_6_14 bitb_6_15 R_bl
Cb_6_14 bit_6_14 gnd C_bl
Cbb_6_14 bitb_6_14 gnd C_bl
Rb_6_15 bit_6_15 bit_6_16 R_bl
Rbb_6_15 bitb_6_15 bitb_6_16 R_bl
Cb_6_15 bit_6_15 gnd C_bl
Cbb_6_15 bitb_6_15 gnd C_bl
Rb_6_16 bit_6_16 bit_6_17 R_bl
Rbb_6_16 bitb_6_16 bitb_6_17 R_bl
Cb_6_16 bit_6_16 gnd C_bl
Cbb_6_16 bitb_6_16 gnd C_bl
Rb_6_17 bit_6_17 bit_6_18 R_bl
Rbb_6_17 bitb_6_17 bitb_6_18 R_bl
Cb_6_17 bit_6_17 gnd C_bl
Cbb_6_17 bitb_6_17 gnd C_bl
Rb_6_18 bit_6_18 bit_6_19 R_bl
Rbb_6_18 bitb_6_18 bitb_6_19 R_bl
Cb_6_18 bit_6_18 gnd C_bl
Cbb_6_18 bitb_6_18 gnd C_bl
Rb_6_19 bit_6_19 bit_6_20 R_bl
Rbb_6_19 bitb_6_19 bitb_6_20 R_bl
Cb_6_19 bit_6_19 gnd C_bl
Cbb_6_19 bitb_6_19 gnd C_bl
Rb_6_20 bit_6_20 bit_6_21 R_bl
Rbb_6_20 bitb_6_20 bitb_6_21 R_bl
Cb_6_20 bit_6_20 gnd C_bl
Cbb_6_20 bitb_6_20 gnd C_bl
Rb_6_21 bit_6_21 bit_6_22 R_bl
Rbb_6_21 bitb_6_21 bitb_6_22 R_bl
Cb_6_21 bit_6_21 gnd C_bl
Cbb_6_21 bitb_6_21 gnd C_bl
Rb_6_22 bit_6_22 bit_6_23 R_bl
Rbb_6_22 bitb_6_22 bitb_6_23 R_bl
Cb_6_22 bit_6_22 gnd C_bl
Cbb_6_22 bitb_6_22 gnd C_bl
Rb_6_23 bit_6_23 bit_6_24 R_bl
Rbb_6_23 bitb_6_23 bitb_6_24 R_bl
Cb_6_23 bit_6_23 gnd C_bl
Cbb_6_23 bitb_6_23 gnd C_bl
Rb_6_24 bit_6_24 bit_6_25 R_bl
Rbb_6_24 bitb_6_24 bitb_6_25 R_bl
Cb_6_24 bit_6_24 gnd C_bl
Cbb_6_24 bitb_6_24 gnd C_bl
Rb_6_25 bit_6_25 bit_6_26 R_bl
Rbb_6_25 bitb_6_25 bitb_6_26 R_bl
Cb_6_25 bit_6_25 gnd C_bl
Cbb_6_25 bitb_6_25 gnd C_bl
Rb_6_26 bit_6_26 bit_6_27 R_bl
Rbb_6_26 bitb_6_26 bitb_6_27 R_bl
Cb_6_26 bit_6_26 gnd C_bl
Cbb_6_26 bitb_6_26 gnd C_bl
Rb_6_27 bit_6_27 bit_6_28 R_bl
Rbb_6_27 bitb_6_27 bitb_6_28 R_bl
Cb_6_27 bit_6_27 gnd C_bl
Cbb_6_27 bitb_6_27 gnd C_bl
Rb_6_28 bit_6_28 bit_6_29 R_bl
Rbb_6_28 bitb_6_28 bitb_6_29 R_bl
Cb_6_28 bit_6_28 gnd C_bl
Cbb_6_28 bitb_6_28 gnd C_bl
Rb_6_29 bit_6_29 bit_6_30 R_bl
Rbb_6_29 bitb_6_29 bitb_6_30 R_bl
Cb_6_29 bit_6_29 gnd C_bl
Cbb_6_29 bitb_6_29 gnd C_bl
Rb_6_30 bit_6_30 bit_6_31 R_bl
Rbb_6_30 bitb_6_30 bitb_6_31 R_bl
Cb_6_30 bit_6_30 gnd C_bl
Cbb_6_30 bitb_6_30 gnd C_bl
Rb_6_31 bit_6_31 bit_6_32 R_bl
Rbb_6_31 bitb_6_31 bitb_6_32 R_bl
Cb_6_31 bit_6_31 gnd C_bl
Cbb_6_31 bitb_6_31 gnd C_bl
Rb_6_32 bit_6_32 bit_6_33 R_bl
Rbb_6_32 bitb_6_32 bitb_6_33 R_bl
Cb_6_32 bit_6_32 gnd C_bl
Cbb_6_32 bitb_6_32 gnd C_bl
Rb_6_33 bit_6_33 bit_6_34 R_bl
Rbb_6_33 bitb_6_33 bitb_6_34 R_bl
Cb_6_33 bit_6_33 gnd C_bl
Cbb_6_33 bitb_6_33 gnd C_bl
Rb_6_34 bit_6_34 bit_6_35 R_bl
Rbb_6_34 bitb_6_34 bitb_6_35 R_bl
Cb_6_34 bit_6_34 gnd C_bl
Cbb_6_34 bitb_6_34 gnd C_bl
Rb_6_35 bit_6_35 bit_6_36 R_bl
Rbb_6_35 bitb_6_35 bitb_6_36 R_bl
Cb_6_35 bit_6_35 gnd C_bl
Cbb_6_35 bitb_6_35 gnd C_bl
Rb_6_36 bit_6_36 bit_6_37 R_bl
Rbb_6_36 bitb_6_36 bitb_6_37 R_bl
Cb_6_36 bit_6_36 gnd C_bl
Cbb_6_36 bitb_6_36 gnd C_bl
Rb_6_37 bit_6_37 bit_6_38 R_bl
Rbb_6_37 bitb_6_37 bitb_6_38 R_bl
Cb_6_37 bit_6_37 gnd C_bl
Cbb_6_37 bitb_6_37 gnd C_bl
Rb_6_38 bit_6_38 bit_6_39 R_bl
Rbb_6_38 bitb_6_38 bitb_6_39 R_bl
Cb_6_38 bit_6_38 gnd C_bl
Cbb_6_38 bitb_6_38 gnd C_bl
Rb_6_39 bit_6_39 bit_6_40 R_bl
Rbb_6_39 bitb_6_39 bitb_6_40 R_bl
Cb_6_39 bit_6_39 gnd C_bl
Cbb_6_39 bitb_6_39 gnd C_bl
Rb_6_40 bit_6_40 bit_6_41 R_bl
Rbb_6_40 bitb_6_40 bitb_6_41 R_bl
Cb_6_40 bit_6_40 gnd C_bl
Cbb_6_40 bitb_6_40 gnd C_bl
Rb_6_41 bit_6_41 bit_6_42 R_bl
Rbb_6_41 bitb_6_41 bitb_6_42 R_bl
Cb_6_41 bit_6_41 gnd C_bl
Cbb_6_41 bitb_6_41 gnd C_bl
Rb_6_42 bit_6_42 bit_6_43 R_bl
Rbb_6_42 bitb_6_42 bitb_6_43 R_bl
Cb_6_42 bit_6_42 gnd C_bl
Cbb_6_42 bitb_6_42 gnd C_bl
Rb_6_43 bit_6_43 bit_6_44 R_bl
Rbb_6_43 bitb_6_43 bitb_6_44 R_bl
Cb_6_43 bit_6_43 gnd C_bl
Cbb_6_43 bitb_6_43 gnd C_bl
Rb_6_44 bit_6_44 bit_6_45 R_bl
Rbb_6_44 bitb_6_44 bitb_6_45 R_bl
Cb_6_44 bit_6_44 gnd C_bl
Cbb_6_44 bitb_6_44 gnd C_bl
Rb_6_45 bit_6_45 bit_6_46 R_bl
Rbb_6_45 bitb_6_45 bitb_6_46 R_bl
Cb_6_45 bit_6_45 gnd C_bl
Cbb_6_45 bitb_6_45 gnd C_bl
Rb_6_46 bit_6_46 bit_6_47 R_bl
Rbb_6_46 bitb_6_46 bitb_6_47 R_bl
Cb_6_46 bit_6_46 gnd C_bl
Cbb_6_46 bitb_6_46 gnd C_bl
Rb_6_47 bit_6_47 bit_6_48 R_bl
Rbb_6_47 bitb_6_47 bitb_6_48 R_bl
Cb_6_47 bit_6_47 gnd C_bl
Cbb_6_47 bitb_6_47 gnd C_bl
Rb_6_48 bit_6_48 bit_6_49 R_bl
Rbb_6_48 bitb_6_48 bitb_6_49 R_bl
Cb_6_48 bit_6_48 gnd C_bl
Cbb_6_48 bitb_6_48 gnd C_bl
Rb_6_49 bit_6_49 bit_6_50 R_bl
Rbb_6_49 bitb_6_49 bitb_6_50 R_bl
Cb_6_49 bit_6_49 gnd C_bl
Cbb_6_49 bitb_6_49 gnd C_bl
Rb_6_50 bit_6_50 bit_6_51 R_bl
Rbb_6_50 bitb_6_50 bitb_6_51 R_bl
Cb_6_50 bit_6_50 gnd C_bl
Cbb_6_50 bitb_6_50 gnd C_bl
Rb_6_51 bit_6_51 bit_6_52 R_bl
Rbb_6_51 bitb_6_51 bitb_6_52 R_bl
Cb_6_51 bit_6_51 gnd C_bl
Cbb_6_51 bitb_6_51 gnd C_bl
Rb_6_52 bit_6_52 bit_6_53 R_bl
Rbb_6_52 bitb_6_52 bitb_6_53 R_bl
Cb_6_52 bit_6_52 gnd C_bl
Cbb_6_52 bitb_6_52 gnd C_bl
Rb_6_53 bit_6_53 bit_6_54 R_bl
Rbb_6_53 bitb_6_53 bitb_6_54 R_bl
Cb_6_53 bit_6_53 gnd C_bl
Cbb_6_53 bitb_6_53 gnd C_bl
Rb_6_54 bit_6_54 bit_6_55 R_bl
Rbb_6_54 bitb_6_54 bitb_6_55 R_bl
Cb_6_54 bit_6_54 gnd C_bl
Cbb_6_54 bitb_6_54 gnd C_bl
Rb_6_55 bit_6_55 bit_6_56 R_bl
Rbb_6_55 bitb_6_55 bitb_6_56 R_bl
Cb_6_55 bit_6_55 gnd C_bl
Cbb_6_55 bitb_6_55 gnd C_bl
Rb_6_56 bit_6_56 bit_6_57 R_bl
Rbb_6_56 bitb_6_56 bitb_6_57 R_bl
Cb_6_56 bit_6_56 gnd C_bl
Cbb_6_56 bitb_6_56 gnd C_bl
Rb_6_57 bit_6_57 bit_6_58 R_bl
Rbb_6_57 bitb_6_57 bitb_6_58 R_bl
Cb_6_57 bit_6_57 gnd C_bl
Cbb_6_57 bitb_6_57 gnd C_bl
Rb_6_58 bit_6_58 bit_6_59 R_bl
Rbb_6_58 bitb_6_58 bitb_6_59 R_bl
Cb_6_58 bit_6_58 gnd C_bl
Cbb_6_58 bitb_6_58 gnd C_bl
Rb_6_59 bit_6_59 bit_6_60 R_bl
Rbb_6_59 bitb_6_59 bitb_6_60 R_bl
Cb_6_59 bit_6_59 gnd C_bl
Cbb_6_59 bitb_6_59 gnd C_bl
Rb_6_60 bit_6_60 bit_6_61 R_bl
Rbb_6_60 bitb_6_60 bitb_6_61 R_bl
Cb_6_60 bit_6_60 gnd C_bl
Cbb_6_60 bitb_6_60 gnd C_bl
Rb_6_61 bit_6_61 bit_6_62 R_bl
Rbb_6_61 bitb_6_61 bitb_6_62 R_bl
Cb_6_61 bit_6_61 gnd C_bl
Cbb_6_61 bitb_6_61 gnd C_bl
Rb_6_62 bit_6_62 bit_6_63 R_bl
Rbb_6_62 bitb_6_62 bitb_6_63 R_bl
Cb_6_62 bit_6_62 gnd C_bl
Cbb_6_62 bitb_6_62 gnd C_bl
Rb_6_63 bit_6_63 bit_6_64 R_bl
Rbb_6_63 bitb_6_63 bitb_6_64 R_bl
Cb_6_63 bit_6_63 gnd C_bl
Cbb_6_63 bitb_6_63 gnd C_bl
Rb_6_64 bit_6_64 bit_6_65 R_bl
Rbb_6_64 bitb_6_64 bitb_6_65 R_bl
Cb_6_64 bit_6_64 gnd C_bl
Cbb_6_64 bitb_6_64 gnd C_bl
Rb_6_65 bit_6_65 bit_6_66 R_bl
Rbb_6_65 bitb_6_65 bitb_6_66 R_bl
Cb_6_65 bit_6_65 gnd C_bl
Cbb_6_65 bitb_6_65 gnd C_bl
Rb_6_66 bit_6_66 bit_6_67 R_bl
Rbb_6_66 bitb_6_66 bitb_6_67 R_bl
Cb_6_66 bit_6_66 gnd C_bl
Cbb_6_66 bitb_6_66 gnd C_bl
Rb_6_67 bit_6_67 bit_6_68 R_bl
Rbb_6_67 bitb_6_67 bitb_6_68 R_bl
Cb_6_67 bit_6_67 gnd C_bl
Cbb_6_67 bitb_6_67 gnd C_bl
Rb_6_68 bit_6_68 bit_6_69 R_bl
Rbb_6_68 bitb_6_68 bitb_6_69 R_bl
Cb_6_68 bit_6_68 gnd C_bl
Cbb_6_68 bitb_6_68 gnd C_bl
Rb_6_69 bit_6_69 bit_6_70 R_bl
Rbb_6_69 bitb_6_69 bitb_6_70 R_bl
Cb_6_69 bit_6_69 gnd C_bl
Cbb_6_69 bitb_6_69 gnd C_bl
Rb_6_70 bit_6_70 bit_6_71 R_bl
Rbb_6_70 bitb_6_70 bitb_6_71 R_bl
Cb_6_70 bit_6_70 gnd C_bl
Cbb_6_70 bitb_6_70 gnd C_bl
Rb_6_71 bit_6_71 bit_6_72 R_bl
Rbb_6_71 bitb_6_71 bitb_6_72 R_bl
Cb_6_71 bit_6_71 gnd C_bl
Cbb_6_71 bitb_6_71 gnd C_bl
Rb_6_72 bit_6_72 bit_6_73 R_bl
Rbb_6_72 bitb_6_72 bitb_6_73 R_bl
Cb_6_72 bit_6_72 gnd C_bl
Cbb_6_72 bitb_6_72 gnd C_bl
Rb_6_73 bit_6_73 bit_6_74 R_bl
Rbb_6_73 bitb_6_73 bitb_6_74 R_bl
Cb_6_73 bit_6_73 gnd C_bl
Cbb_6_73 bitb_6_73 gnd C_bl
Rb_6_74 bit_6_74 bit_6_75 R_bl
Rbb_6_74 bitb_6_74 bitb_6_75 R_bl
Cb_6_74 bit_6_74 gnd C_bl
Cbb_6_74 bitb_6_74 gnd C_bl
Rb_6_75 bit_6_75 bit_6_76 R_bl
Rbb_6_75 bitb_6_75 bitb_6_76 R_bl
Cb_6_75 bit_6_75 gnd C_bl
Cbb_6_75 bitb_6_75 gnd C_bl
Rb_6_76 bit_6_76 bit_6_77 R_bl
Rbb_6_76 bitb_6_76 bitb_6_77 R_bl
Cb_6_76 bit_6_76 gnd C_bl
Cbb_6_76 bitb_6_76 gnd C_bl
Rb_6_77 bit_6_77 bit_6_78 R_bl
Rbb_6_77 bitb_6_77 bitb_6_78 R_bl
Cb_6_77 bit_6_77 gnd C_bl
Cbb_6_77 bitb_6_77 gnd C_bl
Rb_6_78 bit_6_78 bit_6_79 R_bl
Rbb_6_78 bitb_6_78 bitb_6_79 R_bl
Cb_6_78 bit_6_78 gnd C_bl
Cbb_6_78 bitb_6_78 gnd C_bl
Rb_6_79 bit_6_79 bit_6_80 R_bl
Rbb_6_79 bitb_6_79 bitb_6_80 R_bl
Cb_6_79 bit_6_79 gnd C_bl
Cbb_6_79 bitb_6_79 gnd C_bl
Rb_6_80 bit_6_80 bit_6_81 R_bl
Rbb_6_80 bitb_6_80 bitb_6_81 R_bl
Cb_6_80 bit_6_80 gnd C_bl
Cbb_6_80 bitb_6_80 gnd C_bl
Rb_6_81 bit_6_81 bit_6_82 R_bl
Rbb_6_81 bitb_6_81 bitb_6_82 R_bl
Cb_6_81 bit_6_81 gnd C_bl
Cbb_6_81 bitb_6_81 gnd C_bl
Rb_6_82 bit_6_82 bit_6_83 R_bl
Rbb_6_82 bitb_6_82 bitb_6_83 R_bl
Cb_6_82 bit_6_82 gnd C_bl
Cbb_6_82 bitb_6_82 gnd C_bl
Rb_6_83 bit_6_83 bit_6_84 R_bl
Rbb_6_83 bitb_6_83 bitb_6_84 R_bl
Cb_6_83 bit_6_83 gnd C_bl
Cbb_6_83 bitb_6_83 gnd C_bl
Rb_6_84 bit_6_84 bit_6_85 R_bl
Rbb_6_84 bitb_6_84 bitb_6_85 R_bl
Cb_6_84 bit_6_84 gnd C_bl
Cbb_6_84 bitb_6_84 gnd C_bl
Rb_6_85 bit_6_85 bit_6_86 R_bl
Rbb_6_85 bitb_6_85 bitb_6_86 R_bl
Cb_6_85 bit_6_85 gnd C_bl
Cbb_6_85 bitb_6_85 gnd C_bl
Rb_6_86 bit_6_86 bit_6_87 R_bl
Rbb_6_86 bitb_6_86 bitb_6_87 R_bl
Cb_6_86 bit_6_86 gnd C_bl
Cbb_6_86 bitb_6_86 gnd C_bl
Rb_6_87 bit_6_87 bit_6_88 R_bl
Rbb_6_87 bitb_6_87 bitb_6_88 R_bl
Cb_6_87 bit_6_87 gnd C_bl
Cbb_6_87 bitb_6_87 gnd C_bl
Rb_6_88 bit_6_88 bit_6_89 R_bl
Rbb_6_88 bitb_6_88 bitb_6_89 R_bl
Cb_6_88 bit_6_88 gnd C_bl
Cbb_6_88 bitb_6_88 gnd C_bl
Rb_6_89 bit_6_89 bit_6_90 R_bl
Rbb_6_89 bitb_6_89 bitb_6_90 R_bl
Cb_6_89 bit_6_89 gnd C_bl
Cbb_6_89 bitb_6_89 gnd C_bl
Rb_6_90 bit_6_90 bit_6_91 R_bl
Rbb_6_90 bitb_6_90 bitb_6_91 R_bl
Cb_6_90 bit_6_90 gnd C_bl
Cbb_6_90 bitb_6_90 gnd C_bl
Rb_6_91 bit_6_91 bit_6_92 R_bl
Rbb_6_91 bitb_6_91 bitb_6_92 R_bl
Cb_6_91 bit_6_91 gnd C_bl
Cbb_6_91 bitb_6_91 gnd C_bl
Rb_6_92 bit_6_92 bit_6_93 R_bl
Rbb_6_92 bitb_6_92 bitb_6_93 R_bl
Cb_6_92 bit_6_92 gnd C_bl
Cbb_6_92 bitb_6_92 gnd C_bl
Rb_6_93 bit_6_93 bit_6_94 R_bl
Rbb_6_93 bitb_6_93 bitb_6_94 R_bl
Cb_6_93 bit_6_93 gnd C_bl
Cbb_6_93 bitb_6_93 gnd C_bl
Rb_6_94 bit_6_94 bit_6_95 R_bl
Rbb_6_94 bitb_6_94 bitb_6_95 R_bl
Cb_6_94 bit_6_94 gnd C_bl
Cbb_6_94 bitb_6_94 gnd C_bl
Rb_6_95 bit_6_95 bit_6_96 R_bl
Rbb_6_95 bitb_6_95 bitb_6_96 R_bl
Cb_6_95 bit_6_95 gnd C_bl
Cbb_6_95 bitb_6_95 gnd C_bl
Rb_6_96 bit_6_96 bit_6_97 R_bl
Rbb_6_96 bitb_6_96 bitb_6_97 R_bl
Cb_6_96 bit_6_96 gnd C_bl
Cbb_6_96 bitb_6_96 gnd C_bl
Rb_6_97 bit_6_97 bit_6_98 R_bl
Rbb_6_97 bitb_6_97 bitb_6_98 R_bl
Cb_6_97 bit_6_97 gnd C_bl
Cbb_6_97 bitb_6_97 gnd C_bl
Rb_6_98 bit_6_98 bit_6_99 R_bl
Rbb_6_98 bitb_6_98 bitb_6_99 R_bl
Cb_6_98 bit_6_98 gnd C_bl
Cbb_6_98 bitb_6_98 gnd C_bl
Rb_6_99 bit_6_99 bit_6_100 R_bl
Rbb_6_99 bitb_6_99 bitb_6_100 R_bl
Cb_6_99 bit_6_99 gnd C_bl
Cbb_6_99 bitb_6_99 gnd C_bl
Rb_7_0 bit_7_0 bit_7_1 R_bl
Rbb_7_0 bitb_7_0 bitb_7_1 R_bl
Cb_7_0 bit_7_0 gnd C_bl
Cbb_7_0 bitb_7_0 gnd C_bl
Rb_7_1 bit_7_1 bit_7_2 R_bl
Rbb_7_1 bitb_7_1 bitb_7_2 R_bl
Cb_7_1 bit_7_1 gnd C_bl
Cbb_7_1 bitb_7_1 gnd C_bl
Rb_7_2 bit_7_2 bit_7_3 R_bl
Rbb_7_2 bitb_7_2 bitb_7_3 R_bl
Cb_7_2 bit_7_2 gnd C_bl
Cbb_7_2 bitb_7_2 gnd C_bl
Rb_7_3 bit_7_3 bit_7_4 R_bl
Rbb_7_3 bitb_7_3 bitb_7_4 R_bl
Cb_7_3 bit_7_3 gnd C_bl
Cbb_7_3 bitb_7_3 gnd C_bl
Rb_7_4 bit_7_4 bit_7_5 R_bl
Rbb_7_4 bitb_7_4 bitb_7_5 R_bl
Cb_7_4 bit_7_4 gnd C_bl
Cbb_7_4 bitb_7_4 gnd C_bl
Rb_7_5 bit_7_5 bit_7_6 R_bl
Rbb_7_5 bitb_7_5 bitb_7_6 R_bl
Cb_7_5 bit_7_5 gnd C_bl
Cbb_7_5 bitb_7_5 gnd C_bl
Rb_7_6 bit_7_6 bit_7_7 R_bl
Rbb_7_6 bitb_7_6 bitb_7_7 R_bl
Cb_7_6 bit_7_6 gnd C_bl
Cbb_7_6 bitb_7_6 gnd C_bl
Rb_7_7 bit_7_7 bit_7_8 R_bl
Rbb_7_7 bitb_7_7 bitb_7_8 R_bl
Cb_7_7 bit_7_7 gnd C_bl
Cbb_7_7 bitb_7_7 gnd C_bl
Rb_7_8 bit_7_8 bit_7_9 R_bl
Rbb_7_8 bitb_7_8 bitb_7_9 R_bl
Cb_7_8 bit_7_8 gnd C_bl
Cbb_7_8 bitb_7_8 gnd C_bl
Rb_7_9 bit_7_9 bit_7_10 R_bl
Rbb_7_9 bitb_7_9 bitb_7_10 R_bl
Cb_7_9 bit_7_9 gnd C_bl
Cbb_7_9 bitb_7_9 gnd C_bl
Rb_7_10 bit_7_10 bit_7_11 R_bl
Rbb_7_10 bitb_7_10 bitb_7_11 R_bl
Cb_7_10 bit_7_10 gnd C_bl
Cbb_7_10 bitb_7_10 gnd C_bl
Rb_7_11 bit_7_11 bit_7_12 R_bl
Rbb_7_11 bitb_7_11 bitb_7_12 R_bl
Cb_7_11 bit_7_11 gnd C_bl
Cbb_7_11 bitb_7_11 gnd C_bl
Rb_7_12 bit_7_12 bit_7_13 R_bl
Rbb_7_12 bitb_7_12 bitb_7_13 R_bl
Cb_7_12 bit_7_12 gnd C_bl
Cbb_7_12 bitb_7_12 gnd C_bl
Rb_7_13 bit_7_13 bit_7_14 R_bl
Rbb_7_13 bitb_7_13 bitb_7_14 R_bl
Cb_7_13 bit_7_13 gnd C_bl
Cbb_7_13 bitb_7_13 gnd C_bl
Rb_7_14 bit_7_14 bit_7_15 R_bl
Rbb_7_14 bitb_7_14 bitb_7_15 R_bl
Cb_7_14 bit_7_14 gnd C_bl
Cbb_7_14 bitb_7_14 gnd C_bl
Rb_7_15 bit_7_15 bit_7_16 R_bl
Rbb_7_15 bitb_7_15 bitb_7_16 R_bl
Cb_7_15 bit_7_15 gnd C_bl
Cbb_7_15 bitb_7_15 gnd C_bl
Rb_7_16 bit_7_16 bit_7_17 R_bl
Rbb_7_16 bitb_7_16 bitb_7_17 R_bl
Cb_7_16 bit_7_16 gnd C_bl
Cbb_7_16 bitb_7_16 gnd C_bl
Rb_7_17 bit_7_17 bit_7_18 R_bl
Rbb_7_17 bitb_7_17 bitb_7_18 R_bl
Cb_7_17 bit_7_17 gnd C_bl
Cbb_7_17 bitb_7_17 gnd C_bl
Rb_7_18 bit_7_18 bit_7_19 R_bl
Rbb_7_18 bitb_7_18 bitb_7_19 R_bl
Cb_7_18 bit_7_18 gnd C_bl
Cbb_7_18 bitb_7_18 gnd C_bl
Rb_7_19 bit_7_19 bit_7_20 R_bl
Rbb_7_19 bitb_7_19 bitb_7_20 R_bl
Cb_7_19 bit_7_19 gnd C_bl
Cbb_7_19 bitb_7_19 gnd C_bl
Rb_7_20 bit_7_20 bit_7_21 R_bl
Rbb_7_20 bitb_7_20 bitb_7_21 R_bl
Cb_7_20 bit_7_20 gnd C_bl
Cbb_7_20 bitb_7_20 gnd C_bl
Rb_7_21 bit_7_21 bit_7_22 R_bl
Rbb_7_21 bitb_7_21 bitb_7_22 R_bl
Cb_7_21 bit_7_21 gnd C_bl
Cbb_7_21 bitb_7_21 gnd C_bl
Rb_7_22 bit_7_22 bit_7_23 R_bl
Rbb_7_22 bitb_7_22 bitb_7_23 R_bl
Cb_7_22 bit_7_22 gnd C_bl
Cbb_7_22 bitb_7_22 gnd C_bl
Rb_7_23 bit_7_23 bit_7_24 R_bl
Rbb_7_23 bitb_7_23 bitb_7_24 R_bl
Cb_7_23 bit_7_23 gnd C_bl
Cbb_7_23 bitb_7_23 gnd C_bl
Rb_7_24 bit_7_24 bit_7_25 R_bl
Rbb_7_24 bitb_7_24 bitb_7_25 R_bl
Cb_7_24 bit_7_24 gnd C_bl
Cbb_7_24 bitb_7_24 gnd C_bl
Rb_7_25 bit_7_25 bit_7_26 R_bl
Rbb_7_25 bitb_7_25 bitb_7_26 R_bl
Cb_7_25 bit_7_25 gnd C_bl
Cbb_7_25 bitb_7_25 gnd C_bl
Rb_7_26 bit_7_26 bit_7_27 R_bl
Rbb_7_26 bitb_7_26 bitb_7_27 R_bl
Cb_7_26 bit_7_26 gnd C_bl
Cbb_7_26 bitb_7_26 gnd C_bl
Rb_7_27 bit_7_27 bit_7_28 R_bl
Rbb_7_27 bitb_7_27 bitb_7_28 R_bl
Cb_7_27 bit_7_27 gnd C_bl
Cbb_7_27 bitb_7_27 gnd C_bl
Rb_7_28 bit_7_28 bit_7_29 R_bl
Rbb_7_28 bitb_7_28 bitb_7_29 R_bl
Cb_7_28 bit_7_28 gnd C_bl
Cbb_7_28 bitb_7_28 gnd C_bl
Rb_7_29 bit_7_29 bit_7_30 R_bl
Rbb_7_29 bitb_7_29 bitb_7_30 R_bl
Cb_7_29 bit_7_29 gnd C_bl
Cbb_7_29 bitb_7_29 gnd C_bl
Rb_7_30 bit_7_30 bit_7_31 R_bl
Rbb_7_30 bitb_7_30 bitb_7_31 R_bl
Cb_7_30 bit_7_30 gnd C_bl
Cbb_7_30 bitb_7_30 gnd C_bl
Rb_7_31 bit_7_31 bit_7_32 R_bl
Rbb_7_31 bitb_7_31 bitb_7_32 R_bl
Cb_7_31 bit_7_31 gnd C_bl
Cbb_7_31 bitb_7_31 gnd C_bl
Rb_7_32 bit_7_32 bit_7_33 R_bl
Rbb_7_32 bitb_7_32 bitb_7_33 R_bl
Cb_7_32 bit_7_32 gnd C_bl
Cbb_7_32 bitb_7_32 gnd C_bl
Rb_7_33 bit_7_33 bit_7_34 R_bl
Rbb_7_33 bitb_7_33 bitb_7_34 R_bl
Cb_7_33 bit_7_33 gnd C_bl
Cbb_7_33 bitb_7_33 gnd C_bl
Rb_7_34 bit_7_34 bit_7_35 R_bl
Rbb_7_34 bitb_7_34 bitb_7_35 R_bl
Cb_7_34 bit_7_34 gnd C_bl
Cbb_7_34 bitb_7_34 gnd C_bl
Rb_7_35 bit_7_35 bit_7_36 R_bl
Rbb_7_35 bitb_7_35 bitb_7_36 R_bl
Cb_7_35 bit_7_35 gnd C_bl
Cbb_7_35 bitb_7_35 gnd C_bl
Rb_7_36 bit_7_36 bit_7_37 R_bl
Rbb_7_36 bitb_7_36 bitb_7_37 R_bl
Cb_7_36 bit_7_36 gnd C_bl
Cbb_7_36 bitb_7_36 gnd C_bl
Rb_7_37 bit_7_37 bit_7_38 R_bl
Rbb_7_37 bitb_7_37 bitb_7_38 R_bl
Cb_7_37 bit_7_37 gnd C_bl
Cbb_7_37 bitb_7_37 gnd C_bl
Rb_7_38 bit_7_38 bit_7_39 R_bl
Rbb_7_38 bitb_7_38 bitb_7_39 R_bl
Cb_7_38 bit_7_38 gnd C_bl
Cbb_7_38 bitb_7_38 gnd C_bl
Rb_7_39 bit_7_39 bit_7_40 R_bl
Rbb_7_39 bitb_7_39 bitb_7_40 R_bl
Cb_7_39 bit_7_39 gnd C_bl
Cbb_7_39 bitb_7_39 gnd C_bl
Rb_7_40 bit_7_40 bit_7_41 R_bl
Rbb_7_40 bitb_7_40 bitb_7_41 R_bl
Cb_7_40 bit_7_40 gnd C_bl
Cbb_7_40 bitb_7_40 gnd C_bl
Rb_7_41 bit_7_41 bit_7_42 R_bl
Rbb_7_41 bitb_7_41 bitb_7_42 R_bl
Cb_7_41 bit_7_41 gnd C_bl
Cbb_7_41 bitb_7_41 gnd C_bl
Rb_7_42 bit_7_42 bit_7_43 R_bl
Rbb_7_42 bitb_7_42 bitb_7_43 R_bl
Cb_7_42 bit_7_42 gnd C_bl
Cbb_7_42 bitb_7_42 gnd C_bl
Rb_7_43 bit_7_43 bit_7_44 R_bl
Rbb_7_43 bitb_7_43 bitb_7_44 R_bl
Cb_7_43 bit_7_43 gnd C_bl
Cbb_7_43 bitb_7_43 gnd C_bl
Rb_7_44 bit_7_44 bit_7_45 R_bl
Rbb_7_44 bitb_7_44 bitb_7_45 R_bl
Cb_7_44 bit_7_44 gnd C_bl
Cbb_7_44 bitb_7_44 gnd C_bl
Rb_7_45 bit_7_45 bit_7_46 R_bl
Rbb_7_45 bitb_7_45 bitb_7_46 R_bl
Cb_7_45 bit_7_45 gnd C_bl
Cbb_7_45 bitb_7_45 gnd C_bl
Rb_7_46 bit_7_46 bit_7_47 R_bl
Rbb_7_46 bitb_7_46 bitb_7_47 R_bl
Cb_7_46 bit_7_46 gnd C_bl
Cbb_7_46 bitb_7_46 gnd C_bl
Rb_7_47 bit_7_47 bit_7_48 R_bl
Rbb_7_47 bitb_7_47 bitb_7_48 R_bl
Cb_7_47 bit_7_47 gnd C_bl
Cbb_7_47 bitb_7_47 gnd C_bl
Rb_7_48 bit_7_48 bit_7_49 R_bl
Rbb_7_48 bitb_7_48 bitb_7_49 R_bl
Cb_7_48 bit_7_48 gnd C_bl
Cbb_7_48 bitb_7_48 gnd C_bl
Rb_7_49 bit_7_49 bit_7_50 R_bl
Rbb_7_49 bitb_7_49 bitb_7_50 R_bl
Cb_7_49 bit_7_49 gnd C_bl
Cbb_7_49 bitb_7_49 gnd C_bl
Rb_7_50 bit_7_50 bit_7_51 R_bl
Rbb_7_50 bitb_7_50 bitb_7_51 R_bl
Cb_7_50 bit_7_50 gnd C_bl
Cbb_7_50 bitb_7_50 gnd C_bl
Rb_7_51 bit_7_51 bit_7_52 R_bl
Rbb_7_51 bitb_7_51 bitb_7_52 R_bl
Cb_7_51 bit_7_51 gnd C_bl
Cbb_7_51 bitb_7_51 gnd C_bl
Rb_7_52 bit_7_52 bit_7_53 R_bl
Rbb_7_52 bitb_7_52 bitb_7_53 R_bl
Cb_7_52 bit_7_52 gnd C_bl
Cbb_7_52 bitb_7_52 gnd C_bl
Rb_7_53 bit_7_53 bit_7_54 R_bl
Rbb_7_53 bitb_7_53 bitb_7_54 R_bl
Cb_7_53 bit_7_53 gnd C_bl
Cbb_7_53 bitb_7_53 gnd C_bl
Rb_7_54 bit_7_54 bit_7_55 R_bl
Rbb_7_54 bitb_7_54 bitb_7_55 R_bl
Cb_7_54 bit_7_54 gnd C_bl
Cbb_7_54 bitb_7_54 gnd C_bl
Rb_7_55 bit_7_55 bit_7_56 R_bl
Rbb_7_55 bitb_7_55 bitb_7_56 R_bl
Cb_7_55 bit_7_55 gnd C_bl
Cbb_7_55 bitb_7_55 gnd C_bl
Rb_7_56 bit_7_56 bit_7_57 R_bl
Rbb_7_56 bitb_7_56 bitb_7_57 R_bl
Cb_7_56 bit_7_56 gnd C_bl
Cbb_7_56 bitb_7_56 gnd C_bl
Rb_7_57 bit_7_57 bit_7_58 R_bl
Rbb_7_57 bitb_7_57 bitb_7_58 R_bl
Cb_7_57 bit_7_57 gnd C_bl
Cbb_7_57 bitb_7_57 gnd C_bl
Rb_7_58 bit_7_58 bit_7_59 R_bl
Rbb_7_58 bitb_7_58 bitb_7_59 R_bl
Cb_7_58 bit_7_58 gnd C_bl
Cbb_7_58 bitb_7_58 gnd C_bl
Rb_7_59 bit_7_59 bit_7_60 R_bl
Rbb_7_59 bitb_7_59 bitb_7_60 R_bl
Cb_7_59 bit_7_59 gnd C_bl
Cbb_7_59 bitb_7_59 gnd C_bl
Rb_7_60 bit_7_60 bit_7_61 R_bl
Rbb_7_60 bitb_7_60 bitb_7_61 R_bl
Cb_7_60 bit_7_60 gnd C_bl
Cbb_7_60 bitb_7_60 gnd C_bl
Rb_7_61 bit_7_61 bit_7_62 R_bl
Rbb_7_61 bitb_7_61 bitb_7_62 R_bl
Cb_7_61 bit_7_61 gnd C_bl
Cbb_7_61 bitb_7_61 gnd C_bl
Rb_7_62 bit_7_62 bit_7_63 R_bl
Rbb_7_62 bitb_7_62 bitb_7_63 R_bl
Cb_7_62 bit_7_62 gnd C_bl
Cbb_7_62 bitb_7_62 gnd C_bl
Rb_7_63 bit_7_63 bit_7_64 R_bl
Rbb_7_63 bitb_7_63 bitb_7_64 R_bl
Cb_7_63 bit_7_63 gnd C_bl
Cbb_7_63 bitb_7_63 gnd C_bl
Rb_7_64 bit_7_64 bit_7_65 R_bl
Rbb_7_64 bitb_7_64 bitb_7_65 R_bl
Cb_7_64 bit_7_64 gnd C_bl
Cbb_7_64 bitb_7_64 gnd C_bl
Rb_7_65 bit_7_65 bit_7_66 R_bl
Rbb_7_65 bitb_7_65 bitb_7_66 R_bl
Cb_7_65 bit_7_65 gnd C_bl
Cbb_7_65 bitb_7_65 gnd C_bl
Rb_7_66 bit_7_66 bit_7_67 R_bl
Rbb_7_66 bitb_7_66 bitb_7_67 R_bl
Cb_7_66 bit_7_66 gnd C_bl
Cbb_7_66 bitb_7_66 gnd C_bl
Rb_7_67 bit_7_67 bit_7_68 R_bl
Rbb_7_67 bitb_7_67 bitb_7_68 R_bl
Cb_7_67 bit_7_67 gnd C_bl
Cbb_7_67 bitb_7_67 gnd C_bl
Rb_7_68 bit_7_68 bit_7_69 R_bl
Rbb_7_68 bitb_7_68 bitb_7_69 R_bl
Cb_7_68 bit_7_68 gnd C_bl
Cbb_7_68 bitb_7_68 gnd C_bl
Rb_7_69 bit_7_69 bit_7_70 R_bl
Rbb_7_69 bitb_7_69 bitb_7_70 R_bl
Cb_7_69 bit_7_69 gnd C_bl
Cbb_7_69 bitb_7_69 gnd C_bl
Rb_7_70 bit_7_70 bit_7_71 R_bl
Rbb_7_70 bitb_7_70 bitb_7_71 R_bl
Cb_7_70 bit_7_70 gnd C_bl
Cbb_7_70 bitb_7_70 gnd C_bl
Rb_7_71 bit_7_71 bit_7_72 R_bl
Rbb_7_71 bitb_7_71 bitb_7_72 R_bl
Cb_7_71 bit_7_71 gnd C_bl
Cbb_7_71 bitb_7_71 gnd C_bl
Rb_7_72 bit_7_72 bit_7_73 R_bl
Rbb_7_72 bitb_7_72 bitb_7_73 R_bl
Cb_7_72 bit_7_72 gnd C_bl
Cbb_7_72 bitb_7_72 gnd C_bl
Rb_7_73 bit_7_73 bit_7_74 R_bl
Rbb_7_73 bitb_7_73 bitb_7_74 R_bl
Cb_7_73 bit_7_73 gnd C_bl
Cbb_7_73 bitb_7_73 gnd C_bl
Rb_7_74 bit_7_74 bit_7_75 R_bl
Rbb_7_74 bitb_7_74 bitb_7_75 R_bl
Cb_7_74 bit_7_74 gnd C_bl
Cbb_7_74 bitb_7_74 gnd C_bl
Rb_7_75 bit_7_75 bit_7_76 R_bl
Rbb_7_75 bitb_7_75 bitb_7_76 R_bl
Cb_7_75 bit_7_75 gnd C_bl
Cbb_7_75 bitb_7_75 gnd C_bl
Rb_7_76 bit_7_76 bit_7_77 R_bl
Rbb_7_76 bitb_7_76 bitb_7_77 R_bl
Cb_7_76 bit_7_76 gnd C_bl
Cbb_7_76 bitb_7_76 gnd C_bl
Rb_7_77 bit_7_77 bit_7_78 R_bl
Rbb_7_77 bitb_7_77 bitb_7_78 R_bl
Cb_7_77 bit_7_77 gnd C_bl
Cbb_7_77 bitb_7_77 gnd C_bl
Rb_7_78 bit_7_78 bit_7_79 R_bl
Rbb_7_78 bitb_7_78 bitb_7_79 R_bl
Cb_7_78 bit_7_78 gnd C_bl
Cbb_7_78 bitb_7_78 gnd C_bl
Rb_7_79 bit_7_79 bit_7_80 R_bl
Rbb_7_79 bitb_7_79 bitb_7_80 R_bl
Cb_7_79 bit_7_79 gnd C_bl
Cbb_7_79 bitb_7_79 gnd C_bl
Rb_7_80 bit_7_80 bit_7_81 R_bl
Rbb_7_80 bitb_7_80 bitb_7_81 R_bl
Cb_7_80 bit_7_80 gnd C_bl
Cbb_7_80 bitb_7_80 gnd C_bl
Rb_7_81 bit_7_81 bit_7_82 R_bl
Rbb_7_81 bitb_7_81 bitb_7_82 R_bl
Cb_7_81 bit_7_81 gnd C_bl
Cbb_7_81 bitb_7_81 gnd C_bl
Rb_7_82 bit_7_82 bit_7_83 R_bl
Rbb_7_82 bitb_7_82 bitb_7_83 R_bl
Cb_7_82 bit_7_82 gnd C_bl
Cbb_7_82 bitb_7_82 gnd C_bl
Rb_7_83 bit_7_83 bit_7_84 R_bl
Rbb_7_83 bitb_7_83 bitb_7_84 R_bl
Cb_7_83 bit_7_83 gnd C_bl
Cbb_7_83 bitb_7_83 gnd C_bl
Rb_7_84 bit_7_84 bit_7_85 R_bl
Rbb_7_84 bitb_7_84 bitb_7_85 R_bl
Cb_7_84 bit_7_84 gnd C_bl
Cbb_7_84 bitb_7_84 gnd C_bl
Rb_7_85 bit_7_85 bit_7_86 R_bl
Rbb_7_85 bitb_7_85 bitb_7_86 R_bl
Cb_7_85 bit_7_85 gnd C_bl
Cbb_7_85 bitb_7_85 gnd C_bl
Rb_7_86 bit_7_86 bit_7_87 R_bl
Rbb_7_86 bitb_7_86 bitb_7_87 R_bl
Cb_7_86 bit_7_86 gnd C_bl
Cbb_7_86 bitb_7_86 gnd C_bl
Rb_7_87 bit_7_87 bit_7_88 R_bl
Rbb_7_87 bitb_7_87 bitb_7_88 R_bl
Cb_7_87 bit_7_87 gnd C_bl
Cbb_7_87 bitb_7_87 gnd C_bl
Rb_7_88 bit_7_88 bit_7_89 R_bl
Rbb_7_88 bitb_7_88 bitb_7_89 R_bl
Cb_7_88 bit_7_88 gnd C_bl
Cbb_7_88 bitb_7_88 gnd C_bl
Rb_7_89 bit_7_89 bit_7_90 R_bl
Rbb_7_89 bitb_7_89 bitb_7_90 R_bl
Cb_7_89 bit_7_89 gnd C_bl
Cbb_7_89 bitb_7_89 gnd C_bl
Rb_7_90 bit_7_90 bit_7_91 R_bl
Rbb_7_90 bitb_7_90 bitb_7_91 R_bl
Cb_7_90 bit_7_90 gnd C_bl
Cbb_7_90 bitb_7_90 gnd C_bl
Rb_7_91 bit_7_91 bit_7_92 R_bl
Rbb_7_91 bitb_7_91 bitb_7_92 R_bl
Cb_7_91 bit_7_91 gnd C_bl
Cbb_7_91 bitb_7_91 gnd C_bl
Rb_7_92 bit_7_92 bit_7_93 R_bl
Rbb_7_92 bitb_7_92 bitb_7_93 R_bl
Cb_7_92 bit_7_92 gnd C_bl
Cbb_7_92 bitb_7_92 gnd C_bl
Rb_7_93 bit_7_93 bit_7_94 R_bl
Rbb_7_93 bitb_7_93 bitb_7_94 R_bl
Cb_7_93 bit_7_93 gnd C_bl
Cbb_7_93 bitb_7_93 gnd C_bl
Rb_7_94 bit_7_94 bit_7_95 R_bl
Rbb_7_94 bitb_7_94 bitb_7_95 R_bl
Cb_7_94 bit_7_94 gnd C_bl
Cbb_7_94 bitb_7_94 gnd C_bl
Rb_7_95 bit_7_95 bit_7_96 R_bl
Rbb_7_95 bitb_7_95 bitb_7_96 R_bl
Cb_7_95 bit_7_95 gnd C_bl
Cbb_7_95 bitb_7_95 gnd C_bl
Rb_7_96 bit_7_96 bit_7_97 R_bl
Rbb_7_96 bitb_7_96 bitb_7_97 R_bl
Cb_7_96 bit_7_96 gnd C_bl
Cbb_7_96 bitb_7_96 gnd C_bl
Rb_7_97 bit_7_97 bit_7_98 R_bl
Rbb_7_97 bitb_7_97 bitb_7_98 R_bl
Cb_7_97 bit_7_97 gnd C_bl
Cbb_7_97 bitb_7_97 gnd C_bl
Rb_7_98 bit_7_98 bit_7_99 R_bl
Rbb_7_98 bitb_7_98 bitb_7_99 R_bl
Cb_7_98 bit_7_98 gnd C_bl
Cbb_7_98 bitb_7_98 gnd C_bl
Rb_7_99 bit_7_99 bit_7_100 R_bl
Rbb_7_99 bitb_7_99 bitb_7_100 R_bl
Cb_7_99 bit_7_99 gnd C_bl
Cbb_7_99 bitb_7_99 gnd C_bl
Rb_8_0 bit_8_0 bit_8_1 R_bl
Rbb_8_0 bitb_8_0 bitb_8_1 R_bl
Cb_8_0 bit_8_0 gnd C_bl
Cbb_8_0 bitb_8_0 gnd C_bl
Rb_8_1 bit_8_1 bit_8_2 R_bl
Rbb_8_1 bitb_8_1 bitb_8_2 R_bl
Cb_8_1 bit_8_1 gnd C_bl
Cbb_8_1 bitb_8_1 gnd C_bl
Rb_8_2 bit_8_2 bit_8_3 R_bl
Rbb_8_2 bitb_8_2 bitb_8_3 R_bl
Cb_8_2 bit_8_2 gnd C_bl
Cbb_8_2 bitb_8_2 gnd C_bl
Rb_8_3 bit_8_3 bit_8_4 R_bl
Rbb_8_3 bitb_8_3 bitb_8_4 R_bl
Cb_8_3 bit_8_3 gnd C_bl
Cbb_8_3 bitb_8_3 gnd C_bl
Rb_8_4 bit_8_4 bit_8_5 R_bl
Rbb_8_4 bitb_8_4 bitb_8_5 R_bl
Cb_8_4 bit_8_4 gnd C_bl
Cbb_8_4 bitb_8_4 gnd C_bl
Rb_8_5 bit_8_5 bit_8_6 R_bl
Rbb_8_5 bitb_8_5 bitb_8_6 R_bl
Cb_8_5 bit_8_5 gnd C_bl
Cbb_8_5 bitb_8_5 gnd C_bl
Rb_8_6 bit_8_6 bit_8_7 R_bl
Rbb_8_6 bitb_8_6 bitb_8_7 R_bl
Cb_8_6 bit_8_6 gnd C_bl
Cbb_8_6 bitb_8_6 gnd C_bl
Rb_8_7 bit_8_7 bit_8_8 R_bl
Rbb_8_7 bitb_8_7 bitb_8_8 R_bl
Cb_8_7 bit_8_7 gnd C_bl
Cbb_8_7 bitb_8_7 gnd C_bl
Rb_8_8 bit_8_8 bit_8_9 R_bl
Rbb_8_8 bitb_8_8 bitb_8_9 R_bl
Cb_8_8 bit_8_8 gnd C_bl
Cbb_8_8 bitb_8_8 gnd C_bl
Rb_8_9 bit_8_9 bit_8_10 R_bl
Rbb_8_9 bitb_8_9 bitb_8_10 R_bl
Cb_8_9 bit_8_9 gnd C_bl
Cbb_8_9 bitb_8_9 gnd C_bl
Rb_8_10 bit_8_10 bit_8_11 R_bl
Rbb_8_10 bitb_8_10 bitb_8_11 R_bl
Cb_8_10 bit_8_10 gnd C_bl
Cbb_8_10 bitb_8_10 gnd C_bl
Rb_8_11 bit_8_11 bit_8_12 R_bl
Rbb_8_11 bitb_8_11 bitb_8_12 R_bl
Cb_8_11 bit_8_11 gnd C_bl
Cbb_8_11 bitb_8_11 gnd C_bl
Rb_8_12 bit_8_12 bit_8_13 R_bl
Rbb_8_12 bitb_8_12 bitb_8_13 R_bl
Cb_8_12 bit_8_12 gnd C_bl
Cbb_8_12 bitb_8_12 gnd C_bl
Rb_8_13 bit_8_13 bit_8_14 R_bl
Rbb_8_13 bitb_8_13 bitb_8_14 R_bl
Cb_8_13 bit_8_13 gnd C_bl
Cbb_8_13 bitb_8_13 gnd C_bl
Rb_8_14 bit_8_14 bit_8_15 R_bl
Rbb_8_14 bitb_8_14 bitb_8_15 R_bl
Cb_8_14 bit_8_14 gnd C_bl
Cbb_8_14 bitb_8_14 gnd C_bl
Rb_8_15 bit_8_15 bit_8_16 R_bl
Rbb_8_15 bitb_8_15 bitb_8_16 R_bl
Cb_8_15 bit_8_15 gnd C_bl
Cbb_8_15 bitb_8_15 gnd C_bl
Rb_8_16 bit_8_16 bit_8_17 R_bl
Rbb_8_16 bitb_8_16 bitb_8_17 R_bl
Cb_8_16 bit_8_16 gnd C_bl
Cbb_8_16 bitb_8_16 gnd C_bl
Rb_8_17 bit_8_17 bit_8_18 R_bl
Rbb_8_17 bitb_8_17 bitb_8_18 R_bl
Cb_8_17 bit_8_17 gnd C_bl
Cbb_8_17 bitb_8_17 gnd C_bl
Rb_8_18 bit_8_18 bit_8_19 R_bl
Rbb_8_18 bitb_8_18 bitb_8_19 R_bl
Cb_8_18 bit_8_18 gnd C_bl
Cbb_8_18 bitb_8_18 gnd C_bl
Rb_8_19 bit_8_19 bit_8_20 R_bl
Rbb_8_19 bitb_8_19 bitb_8_20 R_bl
Cb_8_19 bit_8_19 gnd C_bl
Cbb_8_19 bitb_8_19 gnd C_bl
Rb_8_20 bit_8_20 bit_8_21 R_bl
Rbb_8_20 bitb_8_20 bitb_8_21 R_bl
Cb_8_20 bit_8_20 gnd C_bl
Cbb_8_20 bitb_8_20 gnd C_bl
Rb_8_21 bit_8_21 bit_8_22 R_bl
Rbb_8_21 bitb_8_21 bitb_8_22 R_bl
Cb_8_21 bit_8_21 gnd C_bl
Cbb_8_21 bitb_8_21 gnd C_bl
Rb_8_22 bit_8_22 bit_8_23 R_bl
Rbb_8_22 bitb_8_22 bitb_8_23 R_bl
Cb_8_22 bit_8_22 gnd C_bl
Cbb_8_22 bitb_8_22 gnd C_bl
Rb_8_23 bit_8_23 bit_8_24 R_bl
Rbb_8_23 bitb_8_23 bitb_8_24 R_bl
Cb_8_23 bit_8_23 gnd C_bl
Cbb_8_23 bitb_8_23 gnd C_bl
Rb_8_24 bit_8_24 bit_8_25 R_bl
Rbb_8_24 bitb_8_24 bitb_8_25 R_bl
Cb_8_24 bit_8_24 gnd C_bl
Cbb_8_24 bitb_8_24 gnd C_bl
Rb_8_25 bit_8_25 bit_8_26 R_bl
Rbb_8_25 bitb_8_25 bitb_8_26 R_bl
Cb_8_25 bit_8_25 gnd C_bl
Cbb_8_25 bitb_8_25 gnd C_bl
Rb_8_26 bit_8_26 bit_8_27 R_bl
Rbb_8_26 bitb_8_26 bitb_8_27 R_bl
Cb_8_26 bit_8_26 gnd C_bl
Cbb_8_26 bitb_8_26 gnd C_bl
Rb_8_27 bit_8_27 bit_8_28 R_bl
Rbb_8_27 bitb_8_27 bitb_8_28 R_bl
Cb_8_27 bit_8_27 gnd C_bl
Cbb_8_27 bitb_8_27 gnd C_bl
Rb_8_28 bit_8_28 bit_8_29 R_bl
Rbb_8_28 bitb_8_28 bitb_8_29 R_bl
Cb_8_28 bit_8_28 gnd C_bl
Cbb_8_28 bitb_8_28 gnd C_bl
Rb_8_29 bit_8_29 bit_8_30 R_bl
Rbb_8_29 bitb_8_29 bitb_8_30 R_bl
Cb_8_29 bit_8_29 gnd C_bl
Cbb_8_29 bitb_8_29 gnd C_bl
Rb_8_30 bit_8_30 bit_8_31 R_bl
Rbb_8_30 bitb_8_30 bitb_8_31 R_bl
Cb_8_30 bit_8_30 gnd C_bl
Cbb_8_30 bitb_8_30 gnd C_bl
Rb_8_31 bit_8_31 bit_8_32 R_bl
Rbb_8_31 bitb_8_31 bitb_8_32 R_bl
Cb_8_31 bit_8_31 gnd C_bl
Cbb_8_31 bitb_8_31 gnd C_bl
Rb_8_32 bit_8_32 bit_8_33 R_bl
Rbb_8_32 bitb_8_32 bitb_8_33 R_bl
Cb_8_32 bit_8_32 gnd C_bl
Cbb_8_32 bitb_8_32 gnd C_bl
Rb_8_33 bit_8_33 bit_8_34 R_bl
Rbb_8_33 bitb_8_33 bitb_8_34 R_bl
Cb_8_33 bit_8_33 gnd C_bl
Cbb_8_33 bitb_8_33 gnd C_bl
Rb_8_34 bit_8_34 bit_8_35 R_bl
Rbb_8_34 bitb_8_34 bitb_8_35 R_bl
Cb_8_34 bit_8_34 gnd C_bl
Cbb_8_34 bitb_8_34 gnd C_bl
Rb_8_35 bit_8_35 bit_8_36 R_bl
Rbb_8_35 bitb_8_35 bitb_8_36 R_bl
Cb_8_35 bit_8_35 gnd C_bl
Cbb_8_35 bitb_8_35 gnd C_bl
Rb_8_36 bit_8_36 bit_8_37 R_bl
Rbb_8_36 bitb_8_36 bitb_8_37 R_bl
Cb_8_36 bit_8_36 gnd C_bl
Cbb_8_36 bitb_8_36 gnd C_bl
Rb_8_37 bit_8_37 bit_8_38 R_bl
Rbb_8_37 bitb_8_37 bitb_8_38 R_bl
Cb_8_37 bit_8_37 gnd C_bl
Cbb_8_37 bitb_8_37 gnd C_bl
Rb_8_38 bit_8_38 bit_8_39 R_bl
Rbb_8_38 bitb_8_38 bitb_8_39 R_bl
Cb_8_38 bit_8_38 gnd C_bl
Cbb_8_38 bitb_8_38 gnd C_bl
Rb_8_39 bit_8_39 bit_8_40 R_bl
Rbb_8_39 bitb_8_39 bitb_8_40 R_bl
Cb_8_39 bit_8_39 gnd C_bl
Cbb_8_39 bitb_8_39 gnd C_bl
Rb_8_40 bit_8_40 bit_8_41 R_bl
Rbb_8_40 bitb_8_40 bitb_8_41 R_bl
Cb_8_40 bit_8_40 gnd C_bl
Cbb_8_40 bitb_8_40 gnd C_bl
Rb_8_41 bit_8_41 bit_8_42 R_bl
Rbb_8_41 bitb_8_41 bitb_8_42 R_bl
Cb_8_41 bit_8_41 gnd C_bl
Cbb_8_41 bitb_8_41 gnd C_bl
Rb_8_42 bit_8_42 bit_8_43 R_bl
Rbb_8_42 bitb_8_42 bitb_8_43 R_bl
Cb_8_42 bit_8_42 gnd C_bl
Cbb_8_42 bitb_8_42 gnd C_bl
Rb_8_43 bit_8_43 bit_8_44 R_bl
Rbb_8_43 bitb_8_43 bitb_8_44 R_bl
Cb_8_43 bit_8_43 gnd C_bl
Cbb_8_43 bitb_8_43 gnd C_bl
Rb_8_44 bit_8_44 bit_8_45 R_bl
Rbb_8_44 bitb_8_44 bitb_8_45 R_bl
Cb_8_44 bit_8_44 gnd C_bl
Cbb_8_44 bitb_8_44 gnd C_bl
Rb_8_45 bit_8_45 bit_8_46 R_bl
Rbb_8_45 bitb_8_45 bitb_8_46 R_bl
Cb_8_45 bit_8_45 gnd C_bl
Cbb_8_45 bitb_8_45 gnd C_bl
Rb_8_46 bit_8_46 bit_8_47 R_bl
Rbb_8_46 bitb_8_46 bitb_8_47 R_bl
Cb_8_46 bit_8_46 gnd C_bl
Cbb_8_46 bitb_8_46 gnd C_bl
Rb_8_47 bit_8_47 bit_8_48 R_bl
Rbb_8_47 bitb_8_47 bitb_8_48 R_bl
Cb_8_47 bit_8_47 gnd C_bl
Cbb_8_47 bitb_8_47 gnd C_bl
Rb_8_48 bit_8_48 bit_8_49 R_bl
Rbb_8_48 bitb_8_48 bitb_8_49 R_bl
Cb_8_48 bit_8_48 gnd C_bl
Cbb_8_48 bitb_8_48 gnd C_bl
Rb_8_49 bit_8_49 bit_8_50 R_bl
Rbb_8_49 bitb_8_49 bitb_8_50 R_bl
Cb_8_49 bit_8_49 gnd C_bl
Cbb_8_49 bitb_8_49 gnd C_bl
Rb_8_50 bit_8_50 bit_8_51 R_bl
Rbb_8_50 bitb_8_50 bitb_8_51 R_bl
Cb_8_50 bit_8_50 gnd C_bl
Cbb_8_50 bitb_8_50 gnd C_bl
Rb_8_51 bit_8_51 bit_8_52 R_bl
Rbb_8_51 bitb_8_51 bitb_8_52 R_bl
Cb_8_51 bit_8_51 gnd C_bl
Cbb_8_51 bitb_8_51 gnd C_bl
Rb_8_52 bit_8_52 bit_8_53 R_bl
Rbb_8_52 bitb_8_52 bitb_8_53 R_bl
Cb_8_52 bit_8_52 gnd C_bl
Cbb_8_52 bitb_8_52 gnd C_bl
Rb_8_53 bit_8_53 bit_8_54 R_bl
Rbb_8_53 bitb_8_53 bitb_8_54 R_bl
Cb_8_53 bit_8_53 gnd C_bl
Cbb_8_53 bitb_8_53 gnd C_bl
Rb_8_54 bit_8_54 bit_8_55 R_bl
Rbb_8_54 bitb_8_54 bitb_8_55 R_bl
Cb_8_54 bit_8_54 gnd C_bl
Cbb_8_54 bitb_8_54 gnd C_bl
Rb_8_55 bit_8_55 bit_8_56 R_bl
Rbb_8_55 bitb_8_55 bitb_8_56 R_bl
Cb_8_55 bit_8_55 gnd C_bl
Cbb_8_55 bitb_8_55 gnd C_bl
Rb_8_56 bit_8_56 bit_8_57 R_bl
Rbb_8_56 bitb_8_56 bitb_8_57 R_bl
Cb_8_56 bit_8_56 gnd C_bl
Cbb_8_56 bitb_8_56 gnd C_bl
Rb_8_57 bit_8_57 bit_8_58 R_bl
Rbb_8_57 bitb_8_57 bitb_8_58 R_bl
Cb_8_57 bit_8_57 gnd C_bl
Cbb_8_57 bitb_8_57 gnd C_bl
Rb_8_58 bit_8_58 bit_8_59 R_bl
Rbb_8_58 bitb_8_58 bitb_8_59 R_bl
Cb_8_58 bit_8_58 gnd C_bl
Cbb_8_58 bitb_8_58 gnd C_bl
Rb_8_59 bit_8_59 bit_8_60 R_bl
Rbb_8_59 bitb_8_59 bitb_8_60 R_bl
Cb_8_59 bit_8_59 gnd C_bl
Cbb_8_59 bitb_8_59 gnd C_bl
Rb_8_60 bit_8_60 bit_8_61 R_bl
Rbb_8_60 bitb_8_60 bitb_8_61 R_bl
Cb_8_60 bit_8_60 gnd C_bl
Cbb_8_60 bitb_8_60 gnd C_bl
Rb_8_61 bit_8_61 bit_8_62 R_bl
Rbb_8_61 bitb_8_61 bitb_8_62 R_bl
Cb_8_61 bit_8_61 gnd C_bl
Cbb_8_61 bitb_8_61 gnd C_bl
Rb_8_62 bit_8_62 bit_8_63 R_bl
Rbb_8_62 bitb_8_62 bitb_8_63 R_bl
Cb_8_62 bit_8_62 gnd C_bl
Cbb_8_62 bitb_8_62 gnd C_bl
Rb_8_63 bit_8_63 bit_8_64 R_bl
Rbb_8_63 bitb_8_63 bitb_8_64 R_bl
Cb_8_63 bit_8_63 gnd C_bl
Cbb_8_63 bitb_8_63 gnd C_bl
Rb_8_64 bit_8_64 bit_8_65 R_bl
Rbb_8_64 bitb_8_64 bitb_8_65 R_bl
Cb_8_64 bit_8_64 gnd C_bl
Cbb_8_64 bitb_8_64 gnd C_bl
Rb_8_65 bit_8_65 bit_8_66 R_bl
Rbb_8_65 bitb_8_65 bitb_8_66 R_bl
Cb_8_65 bit_8_65 gnd C_bl
Cbb_8_65 bitb_8_65 gnd C_bl
Rb_8_66 bit_8_66 bit_8_67 R_bl
Rbb_8_66 bitb_8_66 bitb_8_67 R_bl
Cb_8_66 bit_8_66 gnd C_bl
Cbb_8_66 bitb_8_66 gnd C_bl
Rb_8_67 bit_8_67 bit_8_68 R_bl
Rbb_8_67 bitb_8_67 bitb_8_68 R_bl
Cb_8_67 bit_8_67 gnd C_bl
Cbb_8_67 bitb_8_67 gnd C_bl
Rb_8_68 bit_8_68 bit_8_69 R_bl
Rbb_8_68 bitb_8_68 bitb_8_69 R_bl
Cb_8_68 bit_8_68 gnd C_bl
Cbb_8_68 bitb_8_68 gnd C_bl
Rb_8_69 bit_8_69 bit_8_70 R_bl
Rbb_8_69 bitb_8_69 bitb_8_70 R_bl
Cb_8_69 bit_8_69 gnd C_bl
Cbb_8_69 bitb_8_69 gnd C_bl
Rb_8_70 bit_8_70 bit_8_71 R_bl
Rbb_8_70 bitb_8_70 bitb_8_71 R_bl
Cb_8_70 bit_8_70 gnd C_bl
Cbb_8_70 bitb_8_70 gnd C_bl
Rb_8_71 bit_8_71 bit_8_72 R_bl
Rbb_8_71 bitb_8_71 bitb_8_72 R_bl
Cb_8_71 bit_8_71 gnd C_bl
Cbb_8_71 bitb_8_71 gnd C_bl
Rb_8_72 bit_8_72 bit_8_73 R_bl
Rbb_8_72 bitb_8_72 bitb_8_73 R_bl
Cb_8_72 bit_8_72 gnd C_bl
Cbb_8_72 bitb_8_72 gnd C_bl
Rb_8_73 bit_8_73 bit_8_74 R_bl
Rbb_8_73 bitb_8_73 bitb_8_74 R_bl
Cb_8_73 bit_8_73 gnd C_bl
Cbb_8_73 bitb_8_73 gnd C_bl
Rb_8_74 bit_8_74 bit_8_75 R_bl
Rbb_8_74 bitb_8_74 bitb_8_75 R_bl
Cb_8_74 bit_8_74 gnd C_bl
Cbb_8_74 bitb_8_74 gnd C_bl
Rb_8_75 bit_8_75 bit_8_76 R_bl
Rbb_8_75 bitb_8_75 bitb_8_76 R_bl
Cb_8_75 bit_8_75 gnd C_bl
Cbb_8_75 bitb_8_75 gnd C_bl
Rb_8_76 bit_8_76 bit_8_77 R_bl
Rbb_8_76 bitb_8_76 bitb_8_77 R_bl
Cb_8_76 bit_8_76 gnd C_bl
Cbb_8_76 bitb_8_76 gnd C_bl
Rb_8_77 bit_8_77 bit_8_78 R_bl
Rbb_8_77 bitb_8_77 bitb_8_78 R_bl
Cb_8_77 bit_8_77 gnd C_bl
Cbb_8_77 bitb_8_77 gnd C_bl
Rb_8_78 bit_8_78 bit_8_79 R_bl
Rbb_8_78 bitb_8_78 bitb_8_79 R_bl
Cb_8_78 bit_8_78 gnd C_bl
Cbb_8_78 bitb_8_78 gnd C_bl
Rb_8_79 bit_8_79 bit_8_80 R_bl
Rbb_8_79 bitb_8_79 bitb_8_80 R_bl
Cb_8_79 bit_8_79 gnd C_bl
Cbb_8_79 bitb_8_79 gnd C_bl
Rb_8_80 bit_8_80 bit_8_81 R_bl
Rbb_8_80 bitb_8_80 bitb_8_81 R_bl
Cb_8_80 bit_8_80 gnd C_bl
Cbb_8_80 bitb_8_80 gnd C_bl
Rb_8_81 bit_8_81 bit_8_82 R_bl
Rbb_8_81 bitb_8_81 bitb_8_82 R_bl
Cb_8_81 bit_8_81 gnd C_bl
Cbb_8_81 bitb_8_81 gnd C_bl
Rb_8_82 bit_8_82 bit_8_83 R_bl
Rbb_8_82 bitb_8_82 bitb_8_83 R_bl
Cb_8_82 bit_8_82 gnd C_bl
Cbb_8_82 bitb_8_82 gnd C_bl
Rb_8_83 bit_8_83 bit_8_84 R_bl
Rbb_8_83 bitb_8_83 bitb_8_84 R_bl
Cb_8_83 bit_8_83 gnd C_bl
Cbb_8_83 bitb_8_83 gnd C_bl
Rb_8_84 bit_8_84 bit_8_85 R_bl
Rbb_8_84 bitb_8_84 bitb_8_85 R_bl
Cb_8_84 bit_8_84 gnd C_bl
Cbb_8_84 bitb_8_84 gnd C_bl
Rb_8_85 bit_8_85 bit_8_86 R_bl
Rbb_8_85 bitb_8_85 bitb_8_86 R_bl
Cb_8_85 bit_8_85 gnd C_bl
Cbb_8_85 bitb_8_85 gnd C_bl
Rb_8_86 bit_8_86 bit_8_87 R_bl
Rbb_8_86 bitb_8_86 bitb_8_87 R_bl
Cb_8_86 bit_8_86 gnd C_bl
Cbb_8_86 bitb_8_86 gnd C_bl
Rb_8_87 bit_8_87 bit_8_88 R_bl
Rbb_8_87 bitb_8_87 bitb_8_88 R_bl
Cb_8_87 bit_8_87 gnd C_bl
Cbb_8_87 bitb_8_87 gnd C_bl
Rb_8_88 bit_8_88 bit_8_89 R_bl
Rbb_8_88 bitb_8_88 bitb_8_89 R_bl
Cb_8_88 bit_8_88 gnd C_bl
Cbb_8_88 bitb_8_88 gnd C_bl
Rb_8_89 bit_8_89 bit_8_90 R_bl
Rbb_8_89 bitb_8_89 bitb_8_90 R_bl
Cb_8_89 bit_8_89 gnd C_bl
Cbb_8_89 bitb_8_89 gnd C_bl
Rb_8_90 bit_8_90 bit_8_91 R_bl
Rbb_8_90 bitb_8_90 bitb_8_91 R_bl
Cb_8_90 bit_8_90 gnd C_bl
Cbb_8_90 bitb_8_90 gnd C_bl
Rb_8_91 bit_8_91 bit_8_92 R_bl
Rbb_8_91 bitb_8_91 bitb_8_92 R_bl
Cb_8_91 bit_8_91 gnd C_bl
Cbb_8_91 bitb_8_91 gnd C_bl
Rb_8_92 bit_8_92 bit_8_93 R_bl
Rbb_8_92 bitb_8_92 bitb_8_93 R_bl
Cb_8_92 bit_8_92 gnd C_bl
Cbb_8_92 bitb_8_92 gnd C_bl
Rb_8_93 bit_8_93 bit_8_94 R_bl
Rbb_8_93 bitb_8_93 bitb_8_94 R_bl
Cb_8_93 bit_8_93 gnd C_bl
Cbb_8_93 bitb_8_93 gnd C_bl
Rb_8_94 bit_8_94 bit_8_95 R_bl
Rbb_8_94 bitb_8_94 bitb_8_95 R_bl
Cb_8_94 bit_8_94 gnd C_bl
Cbb_8_94 bitb_8_94 gnd C_bl
Rb_8_95 bit_8_95 bit_8_96 R_bl
Rbb_8_95 bitb_8_95 bitb_8_96 R_bl
Cb_8_95 bit_8_95 gnd C_bl
Cbb_8_95 bitb_8_95 gnd C_bl
Rb_8_96 bit_8_96 bit_8_97 R_bl
Rbb_8_96 bitb_8_96 bitb_8_97 R_bl
Cb_8_96 bit_8_96 gnd C_bl
Cbb_8_96 bitb_8_96 gnd C_bl
Rb_8_97 bit_8_97 bit_8_98 R_bl
Rbb_8_97 bitb_8_97 bitb_8_98 R_bl
Cb_8_97 bit_8_97 gnd C_bl
Cbb_8_97 bitb_8_97 gnd C_bl
Rb_8_98 bit_8_98 bit_8_99 R_bl
Rbb_8_98 bitb_8_98 bitb_8_99 R_bl
Cb_8_98 bit_8_98 gnd C_bl
Cbb_8_98 bitb_8_98 gnd C_bl
Rb_8_99 bit_8_99 bit_8_100 R_bl
Rbb_8_99 bitb_8_99 bitb_8_100 R_bl
Cb_8_99 bit_8_99 gnd C_bl
Cbb_8_99 bitb_8_99 gnd C_bl
Rb_9_0 bit_9_0 bit_9_1 R_bl
Rbb_9_0 bitb_9_0 bitb_9_1 R_bl
Cb_9_0 bit_9_0 gnd C_bl
Cbb_9_0 bitb_9_0 gnd C_bl
Rb_9_1 bit_9_1 bit_9_2 R_bl
Rbb_9_1 bitb_9_1 bitb_9_2 R_bl
Cb_9_1 bit_9_1 gnd C_bl
Cbb_9_1 bitb_9_1 gnd C_bl
Rb_9_2 bit_9_2 bit_9_3 R_bl
Rbb_9_2 bitb_9_2 bitb_9_3 R_bl
Cb_9_2 bit_9_2 gnd C_bl
Cbb_9_2 bitb_9_2 gnd C_bl
Rb_9_3 bit_9_3 bit_9_4 R_bl
Rbb_9_3 bitb_9_3 bitb_9_4 R_bl
Cb_9_3 bit_9_3 gnd C_bl
Cbb_9_3 bitb_9_3 gnd C_bl
Rb_9_4 bit_9_4 bit_9_5 R_bl
Rbb_9_4 bitb_9_4 bitb_9_5 R_bl
Cb_9_4 bit_9_4 gnd C_bl
Cbb_9_4 bitb_9_4 gnd C_bl
Rb_9_5 bit_9_5 bit_9_6 R_bl
Rbb_9_5 bitb_9_5 bitb_9_6 R_bl
Cb_9_5 bit_9_5 gnd C_bl
Cbb_9_5 bitb_9_5 gnd C_bl
Rb_9_6 bit_9_6 bit_9_7 R_bl
Rbb_9_6 bitb_9_6 bitb_9_7 R_bl
Cb_9_6 bit_9_6 gnd C_bl
Cbb_9_6 bitb_9_6 gnd C_bl
Rb_9_7 bit_9_7 bit_9_8 R_bl
Rbb_9_7 bitb_9_7 bitb_9_8 R_bl
Cb_9_7 bit_9_7 gnd C_bl
Cbb_9_7 bitb_9_7 gnd C_bl
Rb_9_8 bit_9_8 bit_9_9 R_bl
Rbb_9_8 bitb_9_8 bitb_9_9 R_bl
Cb_9_8 bit_9_8 gnd C_bl
Cbb_9_8 bitb_9_8 gnd C_bl
Rb_9_9 bit_9_9 bit_9_10 R_bl
Rbb_9_9 bitb_9_9 bitb_9_10 R_bl
Cb_9_9 bit_9_9 gnd C_bl
Cbb_9_9 bitb_9_9 gnd C_bl
Rb_9_10 bit_9_10 bit_9_11 R_bl
Rbb_9_10 bitb_9_10 bitb_9_11 R_bl
Cb_9_10 bit_9_10 gnd C_bl
Cbb_9_10 bitb_9_10 gnd C_bl
Rb_9_11 bit_9_11 bit_9_12 R_bl
Rbb_9_11 bitb_9_11 bitb_9_12 R_bl
Cb_9_11 bit_9_11 gnd C_bl
Cbb_9_11 bitb_9_11 gnd C_bl
Rb_9_12 bit_9_12 bit_9_13 R_bl
Rbb_9_12 bitb_9_12 bitb_9_13 R_bl
Cb_9_12 bit_9_12 gnd C_bl
Cbb_9_12 bitb_9_12 gnd C_bl
Rb_9_13 bit_9_13 bit_9_14 R_bl
Rbb_9_13 bitb_9_13 bitb_9_14 R_bl
Cb_9_13 bit_9_13 gnd C_bl
Cbb_9_13 bitb_9_13 gnd C_bl
Rb_9_14 bit_9_14 bit_9_15 R_bl
Rbb_9_14 bitb_9_14 bitb_9_15 R_bl
Cb_9_14 bit_9_14 gnd C_bl
Cbb_9_14 bitb_9_14 gnd C_bl
Rb_9_15 bit_9_15 bit_9_16 R_bl
Rbb_9_15 bitb_9_15 bitb_9_16 R_bl
Cb_9_15 bit_9_15 gnd C_bl
Cbb_9_15 bitb_9_15 gnd C_bl
Rb_9_16 bit_9_16 bit_9_17 R_bl
Rbb_9_16 bitb_9_16 bitb_9_17 R_bl
Cb_9_16 bit_9_16 gnd C_bl
Cbb_9_16 bitb_9_16 gnd C_bl
Rb_9_17 bit_9_17 bit_9_18 R_bl
Rbb_9_17 bitb_9_17 bitb_9_18 R_bl
Cb_9_17 bit_9_17 gnd C_bl
Cbb_9_17 bitb_9_17 gnd C_bl
Rb_9_18 bit_9_18 bit_9_19 R_bl
Rbb_9_18 bitb_9_18 bitb_9_19 R_bl
Cb_9_18 bit_9_18 gnd C_bl
Cbb_9_18 bitb_9_18 gnd C_bl
Rb_9_19 bit_9_19 bit_9_20 R_bl
Rbb_9_19 bitb_9_19 bitb_9_20 R_bl
Cb_9_19 bit_9_19 gnd C_bl
Cbb_9_19 bitb_9_19 gnd C_bl
Rb_9_20 bit_9_20 bit_9_21 R_bl
Rbb_9_20 bitb_9_20 bitb_9_21 R_bl
Cb_9_20 bit_9_20 gnd C_bl
Cbb_9_20 bitb_9_20 gnd C_bl
Rb_9_21 bit_9_21 bit_9_22 R_bl
Rbb_9_21 bitb_9_21 bitb_9_22 R_bl
Cb_9_21 bit_9_21 gnd C_bl
Cbb_9_21 bitb_9_21 gnd C_bl
Rb_9_22 bit_9_22 bit_9_23 R_bl
Rbb_9_22 bitb_9_22 bitb_9_23 R_bl
Cb_9_22 bit_9_22 gnd C_bl
Cbb_9_22 bitb_9_22 gnd C_bl
Rb_9_23 bit_9_23 bit_9_24 R_bl
Rbb_9_23 bitb_9_23 bitb_9_24 R_bl
Cb_9_23 bit_9_23 gnd C_bl
Cbb_9_23 bitb_9_23 gnd C_bl
Rb_9_24 bit_9_24 bit_9_25 R_bl
Rbb_9_24 bitb_9_24 bitb_9_25 R_bl
Cb_9_24 bit_9_24 gnd C_bl
Cbb_9_24 bitb_9_24 gnd C_bl
Rb_9_25 bit_9_25 bit_9_26 R_bl
Rbb_9_25 bitb_9_25 bitb_9_26 R_bl
Cb_9_25 bit_9_25 gnd C_bl
Cbb_9_25 bitb_9_25 gnd C_bl
Rb_9_26 bit_9_26 bit_9_27 R_bl
Rbb_9_26 bitb_9_26 bitb_9_27 R_bl
Cb_9_26 bit_9_26 gnd C_bl
Cbb_9_26 bitb_9_26 gnd C_bl
Rb_9_27 bit_9_27 bit_9_28 R_bl
Rbb_9_27 bitb_9_27 bitb_9_28 R_bl
Cb_9_27 bit_9_27 gnd C_bl
Cbb_9_27 bitb_9_27 gnd C_bl
Rb_9_28 bit_9_28 bit_9_29 R_bl
Rbb_9_28 bitb_9_28 bitb_9_29 R_bl
Cb_9_28 bit_9_28 gnd C_bl
Cbb_9_28 bitb_9_28 gnd C_bl
Rb_9_29 bit_9_29 bit_9_30 R_bl
Rbb_9_29 bitb_9_29 bitb_9_30 R_bl
Cb_9_29 bit_9_29 gnd C_bl
Cbb_9_29 bitb_9_29 gnd C_bl
Rb_9_30 bit_9_30 bit_9_31 R_bl
Rbb_9_30 bitb_9_30 bitb_9_31 R_bl
Cb_9_30 bit_9_30 gnd C_bl
Cbb_9_30 bitb_9_30 gnd C_bl
Rb_9_31 bit_9_31 bit_9_32 R_bl
Rbb_9_31 bitb_9_31 bitb_9_32 R_bl
Cb_9_31 bit_9_31 gnd C_bl
Cbb_9_31 bitb_9_31 gnd C_bl
Rb_9_32 bit_9_32 bit_9_33 R_bl
Rbb_9_32 bitb_9_32 bitb_9_33 R_bl
Cb_9_32 bit_9_32 gnd C_bl
Cbb_9_32 bitb_9_32 gnd C_bl
Rb_9_33 bit_9_33 bit_9_34 R_bl
Rbb_9_33 bitb_9_33 bitb_9_34 R_bl
Cb_9_33 bit_9_33 gnd C_bl
Cbb_9_33 bitb_9_33 gnd C_bl
Rb_9_34 bit_9_34 bit_9_35 R_bl
Rbb_9_34 bitb_9_34 bitb_9_35 R_bl
Cb_9_34 bit_9_34 gnd C_bl
Cbb_9_34 bitb_9_34 gnd C_bl
Rb_9_35 bit_9_35 bit_9_36 R_bl
Rbb_9_35 bitb_9_35 bitb_9_36 R_bl
Cb_9_35 bit_9_35 gnd C_bl
Cbb_9_35 bitb_9_35 gnd C_bl
Rb_9_36 bit_9_36 bit_9_37 R_bl
Rbb_9_36 bitb_9_36 bitb_9_37 R_bl
Cb_9_36 bit_9_36 gnd C_bl
Cbb_9_36 bitb_9_36 gnd C_bl
Rb_9_37 bit_9_37 bit_9_38 R_bl
Rbb_9_37 bitb_9_37 bitb_9_38 R_bl
Cb_9_37 bit_9_37 gnd C_bl
Cbb_9_37 bitb_9_37 gnd C_bl
Rb_9_38 bit_9_38 bit_9_39 R_bl
Rbb_9_38 bitb_9_38 bitb_9_39 R_bl
Cb_9_38 bit_9_38 gnd C_bl
Cbb_9_38 bitb_9_38 gnd C_bl
Rb_9_39 bit_9_39 bit_9_40 R_bl
Rbb_9_39 bitb_9_39 bitb_9_40 R_bl
Cb_9_39 bit_9_39 gnd C_bl
Cbb_9_39 bitb_9_39 gnd C_bl
Rb_9_40 bit_9_40 bit_9_41 R_bl
Rbb_9_40 bitb_9_40 bitb_9_41 R_bl
Cb_9_40 bit_9_40 gnd C_bl
Cbb_9_40 bitb_9_40 gnd C_bl
Rb_9_41 bit_9_41 bit_9_42 R_bl
Rbb_9_41 bitb_9_41 bitb_9_42 R_bl
Cb_9_41 bit_9_41 gnd C_bl
Cbb_9_41 bitb_9_41 gnd C_bl
Rb_9_42 bit_9_42 bit_9_43 R_bl
Rbb_9_42 bitb_9_42 bitb_9_43 R_bl
Cb_9_42 bit_9_42 gnd C_bl
Cbb_9_42 bitb_9_42 gnd C_bl
Rb_9_43 bit_9_43 bit_9_44 R_bl
Rbb_9_43 bitb_9_43 bitb_9_44 R_bl
Cb_9_43 bit_9_43 gnd C_bl
Cbb_9_43 bitb_9_43 gnd C_bl
Rb_9_44 bit_9_44 bit_9_45 R_bl
Rbb_9_44 bitb_9_44 bitb_9_45 R_bl
Cb_9_44 bit_9_44 gnd C_bl
Cbb_9_44 bitb_9_44 gnd C_bl
Rb_9_45 bit_9_45 bit_9_46 R_bl
Rbb_9_45 bitb_9_45 bitb_9_46 R_bl
Cb_9_45 bit_9_45 gnd C_bl
Cbb_9_45 bitb_9_45 gnd C_bl
Rb_9_46 bit_9_46 bit_9_47 R_bl
Rbb_9_46 bitb_9_46 bitb_9_47 R_bl
Cb_9_46 bit_9_46 gnd C_bl
Cbb_9_46 bitb_9_46 gnd C_bl
Rb_9_47 bit_9_47 bit_9_48 R_bl
Rbb_9_47 bitb_9_47 bitb_9_48 R_bl
Cb_9_47 bit_9_47 gnd C_bl
Cbb_9_47 bitb_9_47 gnd C_bl
Rb_9_48 bit_9_48 bit_9_49 R_bl
Rbb_9_48 bitb_9_48 bitb_9_49 R_bl
Cb_9_48 bit_9_48 gnd C_bl
Cbb_9_48 bitb_9_48 gnd C_bl
Rb_9_49 bit_9_49 bit_9_50 R_bl
Rbb_9_49 bitb_9_49 bitb_9_50 R_bl
Cb_9_49 bit_9_49 gnd C_bl
Cbb_9_49 bitb_9_49 gnd C_bl
Rb_9_50 bit_9_50 bit_9_51 R_bl
Rbb_9_50 bitb_9_50 bitb_9_51 R_bl
Cb_9_50 bit_9_50 gnd C_bl
Cbb_9_50 bitb_9_50 gnd C_bl
Rb_9_51 bit_9_51 bit_9_52 R_bl
Rbb_9_51 bitb_9_51 bitb_9_52 R_bl
Cb_9_51 bit_9_51 gnd C_bl
Cbb_9_51 bitb_9_51 gnd C_bl
Rb_9_52 bit_9_52 bit_9_53 R_bl
Rbb_9_52 bitb_9_52 bitb_9_53 R_bl
Cb_9_52 bit_9_52 gnd C_bl
Cbb_9_52 bitb_9_52 gnd C_bl
Rb_9_53 bit_9_53 bit_9_54 R_bl
Rbb_9_53 bitb_9_53 bitb_9_54 R_bl
Cb_9_53 bit_9_53 gnd C_bl
Cbb_9_53 bitb_9_53 gnd C_bl
Rb_9_54 bit_9_54 bit_9_55 R_bl
Rbb_9_54 bitb_9_54 bitb_9_55 R_bl
Cb_9_54 bit_9_54 gnd C_bl
Cbb_9_54 bitb_9_54 gnd C_bl
Rb_9_55 bit_9_55 bit_9_56 R_bl
Rbb_9_55 bitb_9_55 bitb_9_56 R_bl
Cb_9_55 bit_9_55 gnd C_bl
Cbb_9_55 bitb_9_55 gnd C_bl
Rb_9_56 bit_9_56 bit_9_57 R_bl
Rbb_9_56 bitb_9_56 bitb_9_57 R_bl
Cb_9_56 bit_9_56 gnd C_bl
Cbb_9_56 bitb_9_56 gnd C_bl
Rb_9_57 bit_9_57 bit_9_58 R_bl
Rbb_9_57 bitb_9_57 bitb_9_58 R_bl
Cb_9_57 bit_9_57 gnd C_bl
Cbb_9_57 bitb_9_57 gnd C_bl
Rb_9_58 bit_9_58 bit_9_59 R_bl
Rbb_9_58 bitb_9_58 bitb_9_59 R_bl
Cb_9_58 bit_9_58 gnd C_bl
Cbb_9_58 bitb_9_58 gnd C_bl
Rb_9_59 bit_9_59 bit_9_60 R_bl
Rbb_9_59 bitb_9_59 bitb_9_60 R_bl
Cb_9_59 bit_9_59 gnd C_bl
Cbb_9_59 bitb_9_59 gnd C_bl
Rb_9_60 bit_9_60 bit_9_61 R_bl
Rbb_9_60 bitb_9_60 bitb_9_61 R_bl
Cb_9_60 bit_9_60 gnd C_bl
Cbb_9_60 bitb_9_60 gnd C_bl
Rb_9_61 bit_9_61 bit_9_62 R_bl
Rbb_9_61 bitb_9_61 bitb_9_62 R_bl
Cb_9_61 bit_9_61 gnd C_bl
Cbb_9_61 bitb_9_61 gnd C_bl
Rb_9_62 bit_9_62 bit_9_63 R_bl
Rbb_9_62 bitb_9_62 bitb_9_63 R_bl
Cb_9_62 bit_9_62 gnd C_bl
Cbb_9_62 bitb_9_62 gnd C_bl
Rb_9_63 bit_9_63 bit_9_64 R_bl
Rbb_9_63 bitb_9_63 bitb_9_64 R_bl
Cb_9_63 bit_9_63 gnd C_bl
Cbb_9_63 bitb_9_63 gnd C_bl
Rb_9_64 bit_9_64 bit_9_65 R_bl
Rbb_9_64 bitb_9_64 bitb_9_65 R_bl
Cb_9_64 bit_9_64 gnd C_bl
Cbb_9_64 bitb_9_64 gnd C_bl
Rb_9_65 bit_9_65 bit_9_66 R_bl
Rbb_9_65 bitb_9_65 bitb_9_66 R_bl
Cb_9_65 bit_9_65 gnd C_bl
Cbb_9_65 bitb_9_65 gnd C_bl
Rb_9_66 bit_9_66 bit_9_67 R_bl
Rbb_9_66 bitb_9_66 bitb_9_67 R_bl
Cb_9_66 bit_9_66 gnd C_bl
Cbb_9_66 bitb_9_66 gnd C_bl
Rb_9_67 bit_9_67 bit_9_68 R_bl
Rbb_9_67 bitb_9_67 bitb_9_68 R_bl
Cb_9_67 bit_9_67 gnd C_bl
Cbb_9_67 bitb_9_67 gnd C_bl
Rb_9_68 bit_9_68 bit_9_69 R_bl
Rbb_9_68 bitb_9_68 bitb_9_69 R_bl
Cb_9_68 bit_9_68 gnd C_bl
Cbb_9_68 bitb_9_68 gnd C_bl
Rb_9_69 bit_9_69 bit_9_70 R_bl
Rbb_9_69 bitb_9_69 bitb_9_70 R_bl
Cb_9_69 bit_9_69 gnd C_bl
Cbb_9_69 bitb_9_69 gnd C_bl
Rb_9_70 bit_9_70 bit_9_71 R_bl
Rbb_9_70 bitb_9_70 bitb_9_71 R_bl
Cb_9_70 bit_9_70 gnd C_bl
Cbb_9_70 bitb_9_70 gnd C_bl
Rb_9_71 bit_9_71 bit_9_72 R_bl
Rbb_9_71 bitb_9_71 bitb_9_72 R_bl
Cb_9_71 bit_9_71 gnd C_bl
Cbb_9_71 bitb_9_71 gnd C_bl
Rb_9_72 bit_9_72 bit_9_73 R_bl
Rbb_9_72 bitb_9_72 bitb_9_73 R_bl
Cb_9_72 bit_9_72 gnd C_bl
Cbb_9_72 bitb_9_72 gnd C_bl
Rb_9_73 bit_9_73 bit_9_74 R_bl
Rbb_9_73 bitb_9_73 bitb_9_74 R_bl
Cb_9_73 bit_9_73 gnd C_bl
Cbb_9_73 bitb_9_73 gnd C_bl
Rb_9_74 bit_9_74 bit_9_75 R_bl
Rbb_9_74 bitb_9_74 bitb_9_75 R_bl
Cb_9_74 bit_9_74 gnd C_bl
Cbb_9_74 bitb_9_74 gnd C_bl
Rb_9_75 bit_9_75 bit_9_76 R_bl
Rbb_9_75 bitb_9_75 bitb_9_76 R_bl
Cb_9_75 bit_9_75 gnd C_bl
Cbb_9_75 bitb_9_75 gnd C_bl
Rb_9_76 bit_9_76 bit_9_77 R_bl
Rbb_9_76 bitb_9_76 bitb_9_77 R_bl
Cb_9_76 bit_9_76 gnd C_bl
Cbb_9_76 bitb_9_76 gnd C_bl
Rb_9_77 bit_9_77 bit_9_78 R_bl
Rbb_9_77 bitb_9_77 bitb_9_78 R_bl
Cb_9_77 bit_9_77 gnd C_bl
Cbb_9_77 bitb_9_77 gnd C_bl
Rb_9_78 bit_9_78 bit_9_79 R_bl
Rbb_9_78 bitb_9_78 bitb_9_79 R_bl
Cb_9_78 bit_9_78 gnd C_bl
Cbb_9_78 bitb_9_78 gnd C_bl
Rb_9_79 bit_9_79 bit_9_80 R_bl
Rbb_9_79 bitb_9_79 bitb_9_80 R_bl
Cb_9_79 bit_9_79 gnd C_bl
Cbb_9_79 bitb_9_79 gnd C_bl
Rb_9_80 bit_9_80 bit_9_81 R_bl
Rbb_9_80 bitb_9_80 bitb_9_81 R_bl
Cb_9_80 bit_9_80 gnd C_bl
Cbb_9_80 bitb_9_80 gnd C_bl
Rb_9_81 bit_9_81 bit_9_82 R_bl
Rbb_9_81 bitb_9_81 bitb_9_82 R_bl
Cb_9_81 bit_9_81 gnd C_bl
Cbb_9_81 bitb_9_81 gnd C_bl
Rb_9_82 bit_9_82 bit_9_83 R_bl
Rbb_9_82 bitb_9_82 bitb_9_83 R_bl
Cb_9_82 bit_9_82 gnd C_bl
Cbb_9_82 bitb_9_82 gnd C_bl
Rb_9_83 bit_9_83 bit_9_84 R_bl
Rbb_9_83 bitb_9_83 bitb_9_84 R_bl
Cb_9_83 bit_9_83 gnd C_bl
Cbb_9_83 bitb_9_83 gnd C_bl
Rb_9_84 bit_9_84 bit_9_85 R_bl
Rbb_9_84 bitb_9_84 bitb_9_85 R_bl
Cb_9_84 bit_9_84 gnd C_bl
Cbb_9_84 bitb_9_84 gnd C_bl
Rb_9_85 bit_9_85 bit_9_86 R_bl
Rbb_9_85 bitb_9_85 bitb_9_86 R_bl
Cb_9_85 bit_9_85 gnd C_bl
Cbb_9_85 bitb_9_85 gnd C_bl
Rb_9_86 bit_9_86 bit_9_87 R_bl
Rbb_9_86 bitb_9_86 bitb_9_87 R_bl
Cb_9_86 bit_9_86 gnd C_bl
Cbb_9_86 bitb_9_86 gnd C_bl
Rb_9_87 bit_9_87 bit_9_88 R_bl
Rbb_9_87 bitb_9_87 bitb_9_88 R_bl
Cb_9_87 bit_9_87 gnd C_bl
Cbb_9_87 bitb_9_87 gnd C_bl
Rb_9_88 bit_9_88 bit_9_89 R_bl
Rbb_9_88 bitb_9_88 bitb_9_89 R_bl
Cb_9_88 bit_9_88 gnd C_bl
Cbb_9_88 bitb_9_88 gnd C_bl
Rb_9_89 bit_9_89 bit_9_90 R_bl
Rbb_9_89 bitb_9_89 bitb_9_90 R_bl
Cb_9_89 bit_9_89 gnd C_bl
Cbb_9_89 bitb_9_89 gnd C_bl
Rb_9_90 bit_9_90 bit_9_91 R_bl
Rbb_9_90 bitb_9_90 bitb_9_91 R_bl
Cb_9_90 bit_9_90 gnd C_bl
Cbb_9_90 bitb_9_90 gnd C_bl
Rb_9_91 bit_9_91 bit_9_92 R_bl
Rbb_9_91 bitb_9_91 bitb_9_92 R_bl
Cb_9_91 bit_9_91 gnd C_bl
Cbb_9_91 bitb_9_91 gnd C_bl
Rb_9_92 bit_9_92 bit_9_93 R_bl
Rbb_9_92 bitb_9_92 bitb_9_93 R_bl
Cb_9_92 bit_9_92 gnd C_bl
Cbb_9_92 bitb_9_92 gnd C_bl
Rb_9_93 bit_9_93 bit_9_94 R_bl
Rbb_9_93 bitb_9_93 bitb_9_94 R_bl
Cb_9_93 bit_9_93 gnd C_bl
Cbb_9_93 bitb_9_93 gnd C_bl
Rb_9_94 bit_9_94 bit_9_95 R_bl
Rbb_9_94 bitb_9_94 bitb_9_95 R_bl
Cb_9_94 bit_9_94 gnd C_bl
Cbb_9_94 bitb_9_94 gnd C_bl
Rb_9_95 bit_9_95 bit_9_96 R_bl
Rbb_9_95 bitb_9_95 bitb_9_96 R_bl
Cb_9_95 bit_9_95 gnd C_bl
Cbb_9_95 bitb_9_95 gnd C_bl
Rb_9_96 bit_9_96 bit_9_97 R_bl
Rbb_9_96 bitb_9_96 bitb_9_97 R_bl
Cb_9_96 bit_9_96 gnd C_bl
Cbb_9_96 bitb_9_96 gnd C_bl
Rb_9_97 bit_9_97 bit_9_98 R_bl
Rbb_9_97 bitb_9_97 bitb_9_98 R_bl
Cb_9_97 bit_9_97 gnd C_bl
Cbb_9_97 bitb_9_97 gnd C_bl
Rb_9_98 bit_9_98 bit_9_99 R_bl
Rbb_9_98 bitb_9_98 bitb_9_99 R_bl
Cb_9_98 bit_9_98 gnd C_bl
Cbb_9_98 bitb_9_98 gnd C_bl
Rb_9_99 bit_9_99 bit_9_100 R_bl
Rbb_9_99 bitb_9_99 bitb_9_100 R_bl
Cb_9_99 bit_9_99 gnd C_bl
Cbb_9_99 bitb_9_99 gnd C_bl
Rb_10_0 bit_10_0 bit_10_1 R_bl
Rbb_10_0 bitb_10_0 bitb_10_1 R_bl
Cb_10_0 bit_10_0 gnd C_bl
Cbb_10_0 bitb_10_0 gnd C_bl
Rb_10_1 bit_10_1 bit_10_2 R_bl
Rbb_10_1 bitb_10_1 bitb_10_2 R_bl
Cb_10_1 bit_10_1 gnd C_bl
Cbb_10_1 bitb_10_1 gnd C_bl
Rb_10_2 bit_10_2 bit_10_3 R_bl
Rbb_10_2 bitb_10_2 bitb_10_3 R_bl
Cb_10_2 bit_10_2 gnd C_bl
Cbb_10_2 bitb_10_2 gnd C_bl
Rb_10_3 bit_10_3 bit_10_4 R_bl
Rbb_10_3 bitb_10_3 bitb_10_4 R_bl
Cb_10_3 bit_10_3 gnd C_bl
Cbb_10_3 bitb_10_3 gnd C_bl
Rb_10_4 bit_10_4 bit_10_5 R_bl
Rbb_10_4 bitb_10_4 bitb_10_5 R_bl
Cb_10_4 bit_10_4 gnd C_bl
Cbb_10_4 bitb_10_4 gnd C_bl
Rb_10_5 bit_10_5 bit_10_6 R_bl
Rbb_10_5 bitb_10_5 bitb_10_6 R_bl
Cb_10_5 bit_10_5 gnd C_bl
Cbb_10_5 bitb_10_5 gnd C_bl
Rb_10_6 bit_10_6 bit_10_7 R_bl
Rbb_10_6 bitb_10_6 bitb_10_7 R_bl
Cb_10_6 bit_10_6 gnd C_bl
Cbb_10_6 bitb_10_6 gnd C_bl
Rb_10_7 bit_10_7 bit_10_8 R_bl
Rbb_10_7 bitb_10_7 bitb_10_8 R_bl
Cb_10_7 bit_10_7 gnd C_bl
Cbb_10_7 bitb_10_7 gnd C_bl
Rb_10_8 bit_10_8 bit_10_9 R_bl
Rbb_10_8 bitb_10_8 bitb_10_9 R_bl
Cb_10_8 bit_10_8 gnd C_bl
Cbb_10_8 bitb_10_8 gnd C_bl
Rb_10_9 bit_10_9 bit_10_10 R_bl
Rbb_10_9 bitb_10_9 bitb_10_10 R_bl
Cb_10_9 bit_10_9 gnd C_bl
Cbb_10_9 bitb_10_9 gnd C_bl
Rb_10_10 bit_10_10 bit_10_11 R_bl
Rbb_10_10 bitb_10_10 bitb_10_11 R_bl
Cb_10_10 bit_10_10 gnd C_bl
Cbb_10_10 bitb_10_10 gnd C_bl
Rb_10_11 bit_10_11 bit_10_12 R_bl
Rbb_10_11 bitb_10_11 bitb_10_12 R_bl
Cb_10_11 bit_10_11 gnd C_bl
Cbb_10_11 bitb_10_11 gnd C_bl
Rb_10_12 bit_10_12 bit_10_13 R_bl
Rbb_10_12 bitb_10_12 bitb_10_13 R_bl
Cb_10_12 bit_10_12 gnd C_bl
Cbb_10_12 bitb_10_12 gnd C_bl
Rb_10_13 bit_10_13 bit_10_14 R_bl
Rbb_10_13 bitb_10_13 bitb_10_14 R_bl
Cb_10_13 bit_10_13 gnd C_bl
Cbb_10_13 bitb_10_13 gnd C_bl
Rb_10_14 bit_10_14 bit_10_15 R_bl
Rbb_10_14 bitb_10_14 bitb_10_15 R_bl
Cb_10_14 bit_10_14 gnd C_bl
Cbb_10_14 bitb_10_14 gnd C_bl
Rb_10_15 bit_10_15 bit_10_16 R_bl
Rbb_10_15 bitb_10_15 bitb_10_16 R_bl
Cb_10_15 bit_10_15 gnd C_bl
Cbb_10_15 bitb_10_15 gnd C_bl
Rb_10_16 bit_10_16 bit_10_17 R_bl
Rbb_10_16 bitb_10_16 bitb_10_17 R_bl
Cb_10_16 bit_10_16 gnd C_bl
Cbb_10_16 bitb_10_16 gnd C_bl
Rb_10_17 bit_10_17 bit_10_18 R_bl
Rbb_10_17 bitb_10_17 bitb_10_18 R_bl
Cb_10_17 bit_10_17 gnd C_bl
Cbb_10_17 bitb_10_17 gnd C_bl
Rb_10_18 bit_10_18 bit_10_19 R_bl
Rbb_10_18 bitb_10_18 bitb_10_19 R_bl
Cb_10_18 bit_10_18 gnd C_bl
Cbb_10_18 bitb_10_18 gnd C_bl
Rb_10_19 bit_10_19 bit_10_20 R_bl
Rbb_10_19 bitb_10_19 bitb_10_20 R_bl
Cb_10_19 bit_10_19 gnd C_bl
Cbb_10_19 bitb_10_19 gnd C_bl
Rb_10_20 bit_10_20 bit_10_21 R_bl
Rbb_10_20 bitb_10_20 bitb_10_21 R_bl
Cb_10_20 bit_10_20 gnd C_bl
Cbb_10_20 bitb_10_20 gnd C_bl
Rb_10_21 bit_10_21 bit_10_22 R_bl
Rbb_10_21 bitb_10_21 bitb_10_22 R_bl
Cb_10_21 bit_10_21 gnd C_bl
Cbb_10_21 bitb_10_21 gnd C_bl
Rb_10_22 bit_10_22 bit_10_23 R_bl
Rbb_10_22 bitb_10_22 bitb_10_23 R_bl
Cb_10_22 bit_10_22 gnd C_bl
Cbb_10_22 bitb_10_22 gnd C_bl
Rb_10_23 bit_10_23 bit_10_24 R_bl
Rbb_10_23 bitb_10_23 bitb_10_24 R_bl
Cb_10_23 bit_10_23 gnd C_bl
Cbb_10_23 bitb_10_23 gnd C_bl
Rb_10_24 bit_10_24 bit_10_25 R_bl
Rbb_10_24 bitb_10_24 bitb_10_25 R_bl
Cb_10_24 bit_10_24 gnd C_bl
Cbb_10_24 bitb_10_24 gnd C_bl
Rb_10_25 bit_10_25 bit_10_26 R_bl
Rbb_10_25 bitb_10_25 bitb_10_26 R_bl
Cb_10_25 bit_10_25 gnd C_bl
Cbb_10_25 bitb_10_25 gnd C_bl
Rb_10_26 bit_10_26 bit_10_27 R_bl
Rbb_10_26 bitb_10_26 bitb_10_27 R_bl
Cb_10_26 bit_10_26 gnd C_bl
Cbb_10_26 bitb_10_26 gnd C_bl
Rb_10_27 bit_10_27 bit_10_28 R_bl
Rbb_10_27 bitb_10_27 bitb_10_28 R_bl
Cb_10_27 bit_10_27 gnd C_bl
Cbb_10_27 bitb_10_27 gnd C_bl
Rb_10_28 bit_10_28 bit_10_29 R_bl
Rbb_10_28 bitb_10_28 bitb_10_29 R_bl
Cb_10_28 bit_10_28 gnd C_bl
Cbb_10_28 bitb_10_28 gnd C_bl
Rb_10_29 bit_10_29 bit_10_30 R_bl
Rbb_10_29 bitb_10_29 bitb_10_30 R_bl
Cb_10_29 bit_10_29 gnd C_bl
Cbb_10_29 bitb_10_29 gnd C_bl
Rb_10_30 bit_10_30 bit_10_31 R_bl
Rbb_10_30 bitb_10_30 bitb_10_31 R_bl
Cb_10_30 bit_10_30 gnd C_bl
Cbb_10_30 bitb_10_30 gnd C_bl
Rb_10_31 bit_10_31 bit_10_32 R_bl
Rbb_10_31 bitb_10_31 bitb_10_32 R_bl
Cb_10_31 bit_10_31 gnd C_bl
Cbb_10_31 bitb_10_31 gnd C_bl
Rb_10_32 bit_10_32 bit_10_33 R_bl
Rbb_10_32 bitb_10_32 bitb_10_33 R_bl
Cb_10_32 bit_10_32 gnd C_bl
Cbb_10_32 bitb_10_32 gnd C_bl
Rb_10_33 bit_10_33 bit_10_34 R_bl
Rbb_10_33 bitb_10_33 bitb_10_34 R_bl
Cb_10_33 bit_10_33 gnd C_bl
Cbb_10_33 bitb_10_33 gnd C_bl
Rb_10_34 bit_10_34 bit_10_35 R_bl
Rbb_10_34 bitb_10_34 bitb_10_35 R_bl
Cb_10_34 bit_10_34 gnd C_bl
Cbb_10_34 bitb_10_34 gnd C_bl
Rb_10_35 bit_10_35 bit_10_36 R_bl
Rbb_10_35 bitb_10_35 bitb_10_36 R_bl
Cb_10_35 bit_10_35 gnd C_bl
Cbb_10_35 bitb_10_35 gnd C_bl
Rb_10_36 bit_10_36 bit_10_37 R_bl
Rbb_10_36 bitb_10_36 bitb_10_37 R_bl
Cb_10_36 bit_10_36 gnd C_bl
Cbb_10_36 bitb_10_36 gnd C_bl
Rb_10_37 bit_10_37 bit_10_38 R_bl
Rbb_10_37 bitb_10_37 bitb_10_38 R_bl
Cb_10_37 bit_10_37 gnd C_bl
Cbb_10_37 bitb_10_37 gnd C_bl
Rb_10_38 bit_10_38 bit_10_39 R_bl
Rbb_10_38 bitb_10_38 bitb_10_39 R_bl
Cb_10_38 bit_10_38 gnd C_bl
Cbb_10_38 bitb_10_38 gnd C_bl
Rb_10_39 bit_10_39 bit_10_40 R_bl
Rbb_10_39 bitb_10_39 bitb_10_40 R_bl
Cb_10_39 bit_10_39 gnd C_bl
Cbb_10_39 bitb_10_39 gnd C_bl
Rb_10_40 bit_10_40 bit_10_41 R_bl
Rbb_10_40 bitb_10_40 bitb_10_41 R_bl
Cb_10_40 bit_10_40 gnd C_bl
Cbb_10_40 bitb_10_40 gnd C_bl
Rb_10_41 bit_10_41 bit_10_42 R_bl
Rbb_10_41 bitb_10_41 bitb_10_42 R_bl
Cb_10_41 bit_10_41 gnd C_bl
Cbb_10_41 bitb_10_41 gnd C_bl
Rb_10_42 bit_10_42 bit_10_43 R_bl
Rbb_10_42 bitb_10_42 bitb_10_43 R_bl
Cb_10_42 bit_10_42 gnd C_bl
Cbb_10_42 bitb_10_42 gnd C_bl
Rb_10_43 bit_10_43 bit_10_44 R_bl
Rbb_10_43 bitb_10_43 bitb_10_44 R_bl
Cb_10_43 bit_10_43 gnd C_bl
Cbb_10_43 bitb_10_43 gnd C_bl
Rb_10_44 bit_10_44 bit_10_45 R_bl
Rbb_10_44 bitb_10_44 bitb_10_45 R_bl
Cb_10_44 bit_10_44 gnd C_bl
Cbb_10_44 bitb_10_44 gnd C_bl
Rb_10_45 bit_10_45 bit_10_46 R_bl
Rbb_10_45 bitb_10_45 bitb_10_46 R_bl
Cb_10_45 bit_10_45 gnd C_bl
Cbb_10_45 bitb_10_45 gnd C_bl
Rb_10_46 bit_10_46 bit_10_47 R_bl
Rbb_10_46 bitb_10_46 bitb_10_47 R_bl
Cb_10_46 bit_10_46 gnd C_bl
Cbb_10_46 bitb_10_46 gnd C_bl
Rb_10_47 bit_10_47 bit_10_48 R_bl
Rbb_10_47 bitb_10_47 bitb_10_48 R_bl
Cb_10_47 bit_10_47 gnd C_bl
Cbb_10_47 bitb_10_47 gnd C_bl
Rb_10_48 bit_10_48 bit_10_49 R_bl
Rbb_10_48 bitb_10_48 bitb_10_49 R_bl
Cb_10_48 bit_10_48 gnd C_bl
Cbb_10_48 bitb_10_48 gnd C_bl
Rb_10_49 bit_10_49 bit_10_50 R_bl
Rbb_10_49 bitb_10_49 bitb_10_50 R_bl
Cb_10_49 bit_10_49 gnd C_bl
Cbb_10_49 bitb_10_49 gnd C_bl
Rb_10_50 bit_10_50 bit_10_51 R_bl
Rbb_10_50 bitb_10_50 bitb_10_51 R_bl
Cb_10_50 bit_10_50 gnd C_bl
Cbb_10_50 bitb_10_50 gnd C_bl
Rb_10_51 bit_10_51 bit_10_52 R_bl
Rbb_10_51 bitb_10_51 bitb_10_52 R_bl
Cb_10_51 bit_10_51 gnd C_bl
Cbb_10_51 bitb_10_51 gnd C_bl
Rb_10_52 bit_10_52 bit_10_53 R_bl
Rbb_10_52 bitb_10_52 bitb_10_53 R_bl
Cb_10_52 bit_10_52 gnd C_bl
Cbb_10_52 bitb_10_52 gnd C_bl
Rb_10_53 bit_10_53 bit_10_54 R_bl
Rbb_10_53 bitb_10_53 bitb_10_54 R_bl
Cb_10_53 bit_10_53 gnd C_bl
Cbb_10_53 bitb_10_53 gnd C_bl
Rb_10_54 bit_10_54 bit_10_55 R_bl
Rbb_10_54 bitb_10_54 bitb_10_55 R_bl
Cb_10_54 bit_10_54 gnd C_bl
Cbb_10_54 bitb_10_54 gnd C_bl
Rb_10_55 bit_10_55 bit_10_56 R_bl
Rbb_10_55 bitb_10_55 bitb_10_56 R_bl
Cb_10_55 bit_10_55 gnd C_bl
Cbb_10_55 bitb_10_55 gnd C_bl
Rb_10_56 bit_10_56 bit_10_57 R_bl
Rbb_10_56 bitb_10_56 bitb_10_57 R_bl
Cb_10_56 bit_10_56 gnd C_bl
Cbb_10_56 bitb_10_56 gnd C_bl
Rb_10_57 bit_10_57 bit_10_58 R_bl
Rbb_10_57 bitb_10_57 bitb_10_58 R_bl
Cb_10_57 bit_10_57 gnd C_bl
Cbb_10_57 bitb_10_57 gnd C_bl
Rb_10_58 bit_10_58 bit_10_59 R_bl
Rbb_10_58 bitb_10_58 bitb_10_59 R_bl
Cb_10_58 bit_10_58 gnd C_bl
Cbb_10_58 bitb_10_58 gnd C_bl
Rb_10_59 bit_10_59 bit_10_60 R_bl
Rbb_10_59 bitb_10_59 bitb_10_60 R_bl
Cb_10_59 bit_10_59 gnd C_bl
Cbb_10_59 bitb_10_59 gnd C_bl
Rb_10_60 bit_10_60 bit_10_61 R_bl
Rbb_10_60 bitb_10_60 bitb_10_61 R_bl
Cb_10_60 bit_10_60 gnd C_bl
Cbb_10_60 bitb_10_60 gnd C_bl
Rb_10_61 bit_10_61 bit_10_62 R_bl
Rbb_10_61 bitb_10_61 bitb_10_62 R_bl
Cb_10_61 bit_10_61 gnd C_bl
Cbb_10_61 bitb_10_61 gnd C_bl
Rb_10_62 bit_10_62 bit_10_63 R_bl
Rbb_10_62 bitb_10_62 bitb_10_63 R_bl
Cb_10_62 bit_10_62 gnd C_bl
Cbb_10_62 bitb_10_62 gnd C_bl
Rb_10_63 bit_10_63 bit_10_64 R_bl
Rbb_10_63 bitb_10_63 bitb_10_64 R_bl
Cb_10_63 bit_10_63 gnd C_bl
Cbb_10_63 bitb_10_63 gnd C_bl
Rb_10_64 bit_10_64 bit_10_65 R_bl
Rbb_10_64 bitb_10_64 bitb_10_65 R_bl
Cb_10_64 bit_10_64 gnd C_bl
Cbb_10_64 bitb_10_64 gnd C_bl
Rb_10_65 bit_10_65 bit_10_66 R_bl
Rbb_10_65 bitb_10_65 bitb_10_66 R_bl
Cb_10_65 bit_10_65 gnd C_bl
Cbb_10_65 bitb_10_65 gnd C_bl
Rb_10_66 bit_10_66 bit_10_67 R_bl
Rbb_10_66 bitb_10_66 bitb_10_67 R_bl
Cb_10_66 bit_10_66 gnd C_bl
Cbb_10_66 bitb_10_66 gnd C_bl
Rb_10_67 bit_10_67 bit_10_68 R_bl
Rbb_10_67 bitb_10_67 bitb_10_68 R_bl
Cb_10_67 bit_10_67 gnd C_bl
Cbb_10_67 bitb_10_67 gnd C_bl
Rb_10_68 bit_10_68 bit_10_69 R_bl
Rbb_10_68 bitb_10_68 bitb_10_69 R_bl
Cb_10_68 bit_10_68 gnd C_bl
Cbb_10_68 bitb_10_68 gnd C_bl
Rb_10_69 bit_10_69 bit_10_70 R_bl
Rbb_10_69 bitb_10_69 bitb_10_70 R_bl
Cb_10_69 bit_10_69 gnd C_bl
Cbb_10_69 bitb_10_69 gnd C_bl
Rb_10_70 bit_10_70 bit_10_71 R_bl
Rbb_10_70 bitb_10_70 bitb_10_71 R_bl
Cb_10_70 bit_10_70 gnd C_bl
Cbb_10_70 bitb_10_70 gnd C_bl
Rb_10_71 bit_10_71 bit_10_72 R_bl
Rbb_10_71 bitb_10_71 bitb_10_72 R_bl
Cb_10_71 bit_10_71 gnd C_bl
Cbb_10_71 bitb_10_71 gnd C_bl
Rb_10_72 bit_10_72 bit_10_73 R_bl
Rbb_10_72 bitb_10_72 bitb_10_73 R_bl
Cb_10_72 bit_10_72 gnd C_bl
Cbb_10_72 bitb_10_72 gnd C_bl
Rb_10_73 bit_10_73 bit_10_74 R_bl
Rbb_10_73 bitb_10_73 bitb_10_74 R_bl
Cb_10_73 bit_10_73 gnd C_bl
Cbb_10_73 bitb_10_73 gnd C_bl
Rb_10_74 bit_10_74 bit_10_75 R_bl
Rbb_10_74 bitb_10_74 bitb_10_75 R_bl
Cb_10_74 bit_10_74 gnd C_bl
Cbb_10_74 bitb_10_74 gnd C_bl
Rb_10_75 bit_10_75 bit_10_76 R_bl
Rbb_10_75 bitb_10_75 bitb_10_76 R_bl
Cb_10_75 bit_10_75 gnd C_bl
Cbb_10_75 bitb_10_75 gnd C_bl
Rb_10_76 bit_10_76 bit_10_77 R_bl
Rbb_10_76 bitb_10_76 bitb_10_77 R_bl
Cb_10_76 bit_10_76 gnd C_bl
Cbb_10_76 bitb_10_76 gnd C_bl
Rb_10_77 bit_10_77 bit_10_78 R_bl
Rbb_10_77 bitb_10_77 bitb_10_78 R_bl
Cb_10_77 bit_10_77 gnd C_bl
Cbb_10_77 bitb_10_77 gnd C_bl
Rb_10_78 bit_10_78 bit_10_79 R_bl
Rbb_10_78 bitb_10_78 bitb_10_79 R_bl
Cb_10_78 bit_10_78 gnd C_bl
Cbb_10_78 bitb_10_78 gnd C_bl
Rb_10_79 bit_10_79 bit_10_80 R_bl
Rbb_10_79 bitb_10_79 bitb_10_80 R_bl
Cb_10_79 bit_10_79 gnd C_bl
Cbb_10_79 bitb_10_79 gnd C_bl
Rb_10_80 bit_10_80 bit_10_81 R_bl
Rbb_10_80 bitb_10_80 bitb_10_81 R_bl
Cb_10_80 bit_10_80 gnd C_bl
Cbb_10_80 bitb_10_80 gnd C_bl
Rb_10_81 bit_10_81 bit_10_82 R_bl
Rbb_10_81 bitb_10_81 bitb_10_82 R_bl
Cb_10_81 bit_10_81 gnd C_bl
Cbb_10_81 bitb_10_81 gnd C_bl
Rb_10_82 bit_10_82 bit_10_83 R_bl
Rbb_10_82 bitb_10_82 bitb_10_83 R_bl
Cb_10_82 bit_10_82 gnd C_bl
Cbb_10_82 bitb_10_82 gnd C_bl
Rb_10_83 bit_10_83 bit_10_84 R_bl
Rbb_10_83 bitb_10_83 bitb_10_84 R_bl
Cb_10_83 bit_10_83 gnd C_bl
Cbb_10_83 bitb_10_83 gnd C_bl
Rb_10_84 bit_10_84 bit_10_85 R_bl
Rbb_10_84 bitb_10_84 bitb_10_85 R_bl
Cb_10_84 bit_10_84 gnd C_bl
Cbb_10_84 bitb_10_84 gnd C_bl
Rb_10_85 bit_10_85 bit_10_86 R_bl
Rbb_10_85 bitb_10_85 bitb_10_86 R_bl
Cb_10_85 bit_10_85 gnd C_bl
Cbb_10_85 bitb_10_85 gnd C_bl
Rb_10_86 bit_10_86 bit_10_87 R_bl
Rbb_10_86 bitb_10_86 bitb_10_87 R_bl
Cb_10_86 bit_10_86 gnd C_bl
Cbb_10_86 bitb_10_86 gnd C_bl
Rb_10_87 bit_10_87 bit_10_88 R_bl
Rbb_10_87 bitb_10_87 bitb_10_88 R_bl
Cb_10_87 bit_10_87 gnd C_bl
Cbb_10_87 bitb_10_87 gnd C_bl
Rb_10_88 bit_10_88 bit_10_89 R_bl
Rbb_10_88 bitb_10_88 bitb_10_89 R_bl
Cb_10_88 bit_10_88 gnd C_bl
Cbb_10_88 bitb_10_88 gnd C_bl
Rb_10_89 bit_10_89 bit_10_90 R_bl
Rbb_10_89 bitb_10_89 bitb_10_90 R_bl
Cb_10_89 bit_10_89 gnd C_bl
Cbb_10_89 bitb_10_89 gnd C_bl
Rb_10_90 bit_10_90 bit_10_91 R_bl
Rbb_10_90 bitb_10_90 bitb_10_91 R_bl
Cb_10_90 bit_10_90 gnd C_bl
Cbb_10_90 bitb_10_90 gnd C_bl
Rb_10_91 bit_10_91 bit_10_92 R_bl
Rbb_10_91 bitb_10_91 bitb_10_92 R_bl
Cb_10_91 bit_10_91 gnd C_bl
Cbb_10_91 bitb_10_91 gnd C_bl
Rb_10_92 bit_10_92 bit_10_93 R_bl
Rbb_10_92 bitb_10_92 bitb_10_93 R_bl
Cb_10_92 bit_10_92 gnd C_bl
Cbb_10_92 bitb_10_92 gnd C_bl
Rb_10_93 bit_10_93 bit_10_94 R_bl
Rbb_10_93 bitb_10_93 bitb_10_94 R_bl
Cb_10_93 bit_10_93 gnd C_bl
Cbb_10_93 bitb_10_93 gnd C_bl
Rb_10_94 bit_10_94 bit_10_95 R_bl
Rbb_10_94 bitb_10_94 bitb_10_95 R_bl
Cb_10_94 bit_10_94 gnd C_bl
Cbb_10_94 bitb_10_94 gnd C_bl
Rb_10_95 bit_10_95 bit_10_96 R_bl
Rbb_10_95 bitb_10_95 bitb_10_96 R_bl
Cb_10_95 bit_10_95 gnd C_bl
Cbb_10_95 bitb_10_95 gnd C_bl
Rb_10_96 bit_10_96 bit_10_97 R_bl
Rbb_10_96 bitb_10_96 bitb_10_97 R_bl
Cb_10_96 bit_10_96 gnd C_bl
Cbb_10_96 bitb_10_96 gnd C_bl
Rb_10_97 bit_10_97 bit_10_98 R_bl
Rbb_10_97 bitb_10_97 bitb_10_98 R_bl
Cb_10_97 bit_10_97 gnd C_bl
Cbb_10_97 bitb_10_97 gnd C_bl
Rb_10_98 bit_10_98 bit_10_99 R_bl
Rbb_10_98 bitb_10_98 bitb_10_99 R_bl
Cb_10_98 bit_10_98 gnd C_bl
Cbb_10_98 bitb_10_98 gnd C_bl
Rb_10_99 bit_10_99 bit_10_100 R_bl
Rbb_10_99 bitb_10_99 bitb_10_100 R_bl
Cb_10_99 bit_10_99 gnd C_bl
Cbb_10_99 bitb_10_99 gnd C_bl
Rb_11_0 bit_11_0 bit_11_1 R_bl
Rbb_11_0 bitb_11_0 bitb_11_1 R_bl
Cb_11_0 bit_11_0 gnd C_bl
Cbb_11_0 bitb_11_0 gnd C_bl
Rb_11_1 bit_11_1 bit_11_2 R_bl
Rbb_11_1 bitb_11_1 bitb_11_2 R_bl
Cb_11_1 bit_11_1 gnd C_bl
Cbb_11_1 bitb_11_1 gnd C_bl
Rb_11_2 bit_11_2 bit_11_3 R_bl
Rbb_11_2 bitb_11_2 bitb_11_3 R_bl
Cb_11_2 bit_11_2 gnd C_bl
Cbb_11_2 bitb_11_2 gnd C_bl
Rb_11_3 bit_11_3 bit_11_4 R_bl
Rbb_11_3 bitb_11_3 bitb_11_4 R_bl
Cb_11_3 bit_11_3 gnd C_bl
Cbb_11_3 bitb_11_3 gnd C_bl
Rb_11_4 bit_11_4 bit_11_5 R_bl
Rbb_11_4 bitb_11_4 bitb_11_5 R_bl
Cb_11_4 bit_11_4 gnd C_bl
Cbb_11_4 bitb_11_4 gnd C_bl
Rb_11_5 bit_11_5 bit_11_6 R_bl
Rbb_11_5 bitb_11_5 bitb_11_6 R_bl
Cb_11_5 bit_11_5 gnd C_bl
Cbb_11_5 bitb_11_5 gnd C_bl
Rb_11_6 bit_11_6 bit_11_7 R_bl
Rbb_11_6 bitb_11_6 bitb_11_7 R_bl
Cb_11_6 bit_11_6 gnd C_bl
Cbb_11_6 bitb_11_6 gnd C_bl
Rb_11_7 bit_11_7 bit_11_8 R_bl
Rbb_11_7 bitb_11_7 bitb_11_8 R_bl
Cb_11_7 bit_11_7 gnd C_bl
Cbb_11_7 bitb_11_7 gnd C_bl
Rb_11_8 bit_11_8 bit_11_9 R_bl
Rbb_11_8 bitb_11_8 bitb_11_9 R_bl
Cb_11_8 bit_11_8 gnd C_bl
Cbb_11_8 bitb_11_8 gnd C_bl
Rb_11_9 bit_11_9 bit_11_10 R_bl
Rbb_11_9 bitb_11_9 bitb_11_10 R_bl
Cb_11_9 bit_11_9 gnd C_bl
Cbb_11_9 bitb_11_9 gnd C_bl
Rb_11_10 bit_11_10 bit_11_11 R_bl
Rbb_11_10 bitb_11_10 bitb_11_11 R_bl
Cb_11_10 bit_11_10 gnd C_bl
Cbb_11_10 bitb_11_10 gnd C_bl
Rb_11_11 bit_11_11 bit_11_12 R_bl
Rbb_11_11 bitb_11_11 bitb_11_12 R_bl
Cb_11_11 bit_11_11 gnd C_bl
Cbb_11_11 bitb_11_11 gnd C_bl
Rb_11_12 bit_11_12 bit_11_13 R_bl
Rbb_11_12 bitb_11_12 bitb_11_13 R_bl
Cb_11_12 bit_11_12 gnd C_bl
Cbb_11_12 bitb_11_12 gnd C_bl
Rb_11_13 bit_11_13 bit_11_14 R_bl
Rbb_11_13 bitb_11_13 bitb_11_14 R_bl
Cb_11_13 bit_11_13 gnd C_bl
Cbb_11_13 bitb_11_13 gnd C_bl
Rb_11_14 bit_11_14 bit_11_15 R_bl
Rbb_11_14 bitb_11_14 bitb_11_15 R_bl
Cb_11_14 bit_11_14 gnd C_bl
Cbb_11_14 bitb_11_14 gnd C_bl
Rb_11_15 bit_11_15 bit_11_16 R_bl
Rbb_11_15 bitb_11_15 bitb_11_16 R_bl
Cb_11_15 bit_11_15 gnd C_bl
Cbb_11_15 bitb_11_15 gnd C_bl
Rb_11_16 bit_11_16 bit_11_17 R_bl
Rbb_11_16 bitb_11_16 bitb_11_17 R_bl
Cb_11_16 bit_11_16 gnd C_bl
Cbb_11_16 bitb_11_16 gnd C_bl
Rb_11_17 bit_11_17 bit_11_18 R_bl
Rbb_11_17 bitb_11_17 bitb_11_18 R_bl
Cb_11_17 bit_11_17 gnd C_bl
Cbb_11_17 bitb_11_17 gnd C_bl
Rb_11_18 bit_11_18 bit_11_19 R_bl
Rbb_11_18 bitb_11_18 bitb_11_19 R_bl
Cb_11_18 bit_11_18 gnd C_bl
Cbb_11_18 bitb_11_18 gnd C_bl
Rb_11_19 bit_11_19 bit_11_20 R_bl
Rbb_11_19 bitb_11_19 bitb_11_20 R_bl
Cb_11_19 bit_11_19 gnd C_bl
Cbb_11_19 bitb_11_19 gnd C_bl
Rb_11_20 bit_11_20 bit_11_21 R_bl
Rbb_11_20 bitb_11_20 bitb_11_21 R_bl
Cb_11_20 bit_11_20 gnd C_bl
Cbb_11_20 bitb_11_20 gnd C_bl
Rb_11_21 bit_11_21 bit_11_22 R_bl
Rbb_11_21 bitb_11_21 bitb_11_22 R_bl
Cb_11_21 bit_11_21 gnd C_bl
Cbb_11_21 bitb_11_21 gnd C_bl
Rb_11_22 bit_11_22 bit_11_23 R_bl
Rbb_11_22 bitb_11_22 bitb_11_23 R_bl
Cb_11_22 bit_11_22 gnd C_bl
Cbb_11_22 bitb_11_22 gnd C_bl
Rb_11_23 bit_11_23 bit_11_24 R_bl
Rbb_11_23 bitb_11_23 bitb_11_24 R_bl
Cb_11_23 bit_11_23 gnd C_bl
Cbb_11_23 bitb_11_23 gnd C_bl
Rb_11_24 bit_11_24 bit_11_25 R_bl
Rbb_11_24 bitb_11_24 bitb_11_25 R_bl
Cb_11_24 bit_11_24 gnd C_bl
Cbb_11_24 bitb_11_24 gnd C_bl
Rb_11_25 bit_11_25 bit_11_26 R_bl
Rbb_11_25 bitb_11_25 bitb_11_26 R_bl
Cb_11_25 bit_11_25 gnd C_bl
Cbb_11_25 bitb_11_25 gnd C_bl
Rb_11_26 bit_11_26 bit_11_27 R_bl
Rbb_11_26 bitb_11_26 bitb_11_27 R_bl
Cb_11_26 bit_11_26 gnd C_bl
Cbb_11_26 bitb_11_26 gnd C_bl
Rb_11_27 bit_11_27 bit_11_28 R_bl
Rbb_11_27 bitb_11_27 bitb_11_28 R_bl
Cb_11_27 bit_11_27 gnd C_bl
Cbb_11_27 bitb_11_27 gnd C_bl
Rb_11_28 bit_11_28 bit_11_29 R_bl
Rbb_11_28 bitb_11_28 bitb_11_29 R_bl
Cb_11_28 bit_11_28 gnd C_bl
Cbb_11_28 bitb_11_28 gnd C_bl
Rb_11_29 bit_11_29 bit_11_30 R_bl
Rbb_11_29 bitb_11_29 bitb_11_30 R_bl
Cb_11_29 bit_11_29 gnd C_bl
Cbb_11_29 bitb_11_29 gnd C_bl
Rb_11_30 bit_11_30 bit_11_31 R_bl
Rbb_11_30 bitb_11_30 bitb_11_31 R_bl
Cb_11_30 bit_11_30 gnd C_bl
Cbb_11_30 bitb_11_30 gnd C_bl
Rb_11_31 bit_11_31 bit_11_32 R_bl
Rbb_11_31 bitb_11_31 bitb_11_32 R_bl
Cb_11_31 bit_11_31 gnd C_bl
Cbb_11_31 bitb_11_31 gnd C_bl
Rb_11_32 bit_11_32 bit_11_33 R_bl
Rbb_11_32 bitb_11_32 bitb_11_33 R_bl
Cb_11_32 bit_11_32 gnd C_bl
Cbb_11_32 bitb_11_32 gnd C_bl
Rb_11_33 bit_11_33 bit_11_34 R_bl
Rbb_11_33 bitb_11_33 bitb_11_34 R_bl
Cb_11_33 bit_11_33 gnd C_bl
Cbb_11_33 bitb_11_33 gnd C_bl
Rb_11_34 bit_11_34 bit_11_35 R_bl
Rbb_11_34 bitb_11_34 bitb_11_35 R_bl
Cb_11_34 bit_11_34 gnd C_bl
Cbb_11_34 bitb_11_34 gnd C_bl
Rb_11_35 bit_11_35 bit_11_36 R_bl
Rbb_11_35 bitb_11_35 bitb_11_36 R_bl
Cb_11_35 bit_11_35 gnd C_bl
Cbb_11_35 bitb_11_35 gnd C_bl
Rb_11_36 bit_11_36 bit_11_37 R_bl
Rbb_11_36 bitb_11_36 bitb_11_37 R_bl
Cb_11_36 bit_11_36 gnd C_bl
Cbb_11_36 bitb_11_36 gnd C_bl
Rb_11_37 bit_11_37 bit_11_38 R_bl
Rbb_11_37 bitb_11_37 bitb_11_38 R_bl
Cb_11_37 bit_11_37 gnd C_bl
Cbb_11_37 bitb_11_37 gnd C_bl
Rb_11_38 bit_11_38 bit_11_39 R_bl
Rbb_11_38 bitb_11_38 bitb_11_39 R_bl
Cb_11_38 bit_11_38 gnd C_bl
Cbb_11_38 bitb_11_38 gnd C_bl
Rb_11_39 bit_11_39 bit_11_40 R_bl
Rbb_11_39 bitb_11_39 bitb_11_40 R_bl
Cb_11_39 bit_11_39 gnd C_bl
Cbb_11_39 bitb_11_39 gnd C_bl
Rb_11_40 bit_11_40 bit_11_41 R_bl
Rbb_11_40 bitb_11_40 bitb_11_41 R_bl
Cb_11_40 bit_11_40 gnd C_bl
Cbb_11_40 bitb_11_40 gnd C_bl
Rb_11_41 bit_11_41 bit_11_42 R_bl
Rbb_11_41 bitb_11_41 bitb_11_42 R_bl
Cb_11_41 bit_11_41 gnd C_bl
Cbb_11_41 bitb_11_41 gnd C_bl
Rb_11_42 bit_11_42 bit_11_43 R_bl
Rbb_11_42 bitb_11_42 bitb_11_43 R_bl
Cb_11_42 bit_11_42 gnd C_bl
Cbb_11_42 bitb_11_42 gnd C_bl
Rb_11_43 bit_11_43 bit_11_44 R_bl
Rbb_11_43 bitb_11_43 bitb_11_44 R_bl
Cb_11_43 bit_11_43 gnd C_bl
Cbb_11_43 bitb_11_43 gnd C_bl
Rb_11_44 bit_11_44 bit_11_45 R_bl
Rbb_11_44 bitb_11_44 bitb_11_45 R_bl
Cb_11_44 bit_11_44 gnd C_bl
Cbb_11_44 bitb_11_44 gnd C_bl
Rb_11_45 bit_11_45 bit_11_46 R_bl
Rbb_11_45 bitb_11_45 bitb_11_46 R_bl
Cb_11_45 bit_11_45 gnd C_bl
Cbb_11_45 bitb_11_45 gnd C_bl
Rb_11_46 bit_11_46 bit_11_47 R_bl
Rbb_11_46 bitb_11_46 bitb_11_47 R_bl
Cb_11_46 bit_11_46 gnd C_bl
Cbb_11_46 bitb_11_46 gnd C_bl
Rb_11_47 bit_11_47 bit_11_48 R_bl
Rbb_11_47 bitb_11_47 bitb_11_48 R_bl
Cb_11_47 bit_11_47 gnd C_bl
Cbb_11_47 bitb_11_47 gnd C_bl
Rb_11_48 bit_11_48 bit_11_49 R_bl
Rbb_11_48 bitb_11_48 bitb_11_49 R_bl
Cb_11_48 bit_11_48 gnd C_bl
Cbb_11_48 bitb_11_48 gnd C_bl
Rb_11_49 bit_11_49 bit_11_50 R_bl
Rbb_11_49 bitb_11_49 bitb_11_50 R_bl
Cb_11_49 bit_11_49 gnd C_bl
Cbb_11_49 bitb_11_49 gnd C_bl
Rb_11_50 bit_11_50 bit_11_51 R_bl
Rbb_11_50 bitb_11_50 bitb_11_51 R_bl
Cb_11_50 bit_11_50 gnd C_bl
Cbb_11_50 bitb_11_50 gnd C_bl
Rb_11_51 bit_11_51 bit_11_52 R_bl
Rbb_11_51 bitb_11_51 bitb_11_52 R_bl
Cb_11_51 bit_11_51 gnd C_bl
Cbb_11_51 bitb_11_51 gnd C_bl
Rb_11_52 bit_11_52 bit_11_53 R_bl
Rbb_11_52 bitb_11_52 bitb_11_53 R_bl
Cb_11_52 bit_11_52 gnd C_bl
Cbb_11_52 bitb_11_52 gnd C_bl
Rb_11_53 bit_11_53 bit_11_54 R_bl
Rbb_11_53 bitb_11_53 bitb_11_54 R_bl
Cb_11_53 bit_11_53 gnd C_bl
Cbb_11_53 bitb_11_53 gnd C_bl
Rb_11_54 bit_11_54 bit_11_55 R_bl
Rbb_11_54 bitb_11_54 bitb_11_55 R_bl
Cb_11_54 bit_11_54 gnd C_bl
Cbb_11_54 bitb_11_54 gnd C_bl
Rb_11_55 bit_11_55 bit_11_56 R_bl
Rbb_11_55 bitb_11_55 bitb_11_56 R_bl
Cb_11_55 bit_11_55 gnd C_bl
Cbb_11_55 bitb_11_55 gnd C_bl
Rb_11_56 bit_11_56 bit_11_57 R_bl
Rbb_11_56 bitb_11_56 bitb_11_57 R_bl
Cb_11_56 bit_11_56 gnd C_bl
Cbb_11_56 bitb_11_56 gnd C_bl
Rb_11_57 bit_11_57 bit_11_58 R_bl
Rbb_11_57 bitb_11_57 bitb_11_58 R_bl
Cb_11_57 bit_11_57 gnd C_bl
Cbb_11_57 bitb_11_57 gnd C_bl
Rb_11_58 bit_11_58 bit_11_59 R_bl
Rbb_11_58 bitb_11_58 bitb_11_59 R_bl
Cb_11_58 bit_11_58 gnd C_bl
Cbb_11_58 bitb_11_58 gnd C_bl
Rb_11_59 bit_11_59 bit_11_60 R_bl
Rbb_11_59 bitb_11_59 bitb_11_60 R_bl
Cb_11_59 bit_11_59 gnd C_bl
Cbb_11_59 bitb_11_59 gnd C_bl
Rb_11_60 bit_11_60 bit_11_61 R_bl
Rbb_11_60 bitb_11_60 bitb_11_61 R_bl
Cb_11_60 bit_11_60 gnd C_bl
Cbb_11_60 bitb_11_60 gnd C_bl
Rb_11_61 bit_11_61 bit_11_62 R_bl
Rbb_11_61 bitb_11_61 bitb_11_62 R_bl
Cb_11_61 bit_11_61 gnd C_bl
Cbb_11_61 bitb_11_61 gnd C_bl
Rb_11_62 bit_11_62 bit_11_63 R_bl
Rbb_11_62 bitb_11_62 bitb_11_63 R_bl
Cb_11_62 bit_11_62 gnd C_bl
Cbb_11_62 bitb_11_62 gnd C_bl
Rb_11_63 bit_11_63 bit_11_64 R_bl
Rbb_11_63 bitb_11_63 bitb_11_64 R_bl
Cb_11_63 bit_11_63 gnd C_bl
Cbb_11_63 bitb_11_63 gnd C_bl
Rb_11_64 bit_11_64 bit_11_65 R_bl
Rbb_11_64 bitb_11_64 bitb_11_65 R_bl
Cb_11_64 bit_11_64 gnd C_bl
Cbb_11_64 bitb_11_64 gnd C_bl
Rb_11_65 bit_11_65 bit_11_66 R_bl
Rbb_11_65 bitb_11_65 bitb_11_66 R_bl
Cb_11_65 bit_11_65 gnd C_bl
Cbb_11_65 bitb_11_65 gnd C_bl
Rb_11_66 bit_11_66 bit_11_67 R_bl
Rbb_11_66 bitb_11_66 bitb_11_67 R_bl
Cb_11_66 bit_11_66 gnd C_bl
Cbb_11_66 bitb_11_66 gnd C_bl
Rb_11_67 bit_11_67 bit_11_68 R_bl
Rbb_11_67 bitb_11_67 bitb_11_68 R_bl
Cb_11_67 bit_11_67 gnd C_bl
Cbb_11_67 bitb_11_67 gnd C_bl
Rb_11_68 bit_11_68 bit_11_69 R_bl
Rbb_11_68 bitb_11_68 bitb_11_69 R_bl
Cb_11_68 bit_11_68 gnd C_bl
Cbb_11_68 bitb_11_68 gnd C_bl
Rb_11_69 bit_11_69 bit_11_70 R_bl
Rbb_11_69 bitb_11_69 bitb_11_70 R_bl
Cb_11_69 bit_11_69 gnd C_bl
Cbb_11_69 bitb_11_69 gnd C_bl
Rb_11_70 bit_11_70 bit_11_71 R_bl
Rbb_11_70 bitb_11_70 bitb_11_71 R_bl
Cb_11_70 bit_11_70 gnd C_bl
Cbb_11_70 bitb_11_70 gnd C_bl
Rb_11_71 bit_11_71 bit_11_72 R_bl
Rbb_11_71 bitb_11_71 bitb_11_72 R_bl
Cb_11_71 bit_11_71 gnd C_bl
Cbb_11_71 bitb_11_71 gnd C_bl
Rb_11_72 bit_11_72 bit_11_73 R_bl
Rbb_11_72 bitb_11_72 bitb_11_73 R_bl
Cb_11_72 bit_11_72 gnd C_bl
Cbb_11_72 bitb_11_72 gnd C_bl
Rb_11_73 bit_11_73 bit_11_74 R_bl
Rbb_11_73 bitb_11_73 bitb_11_74 R_bl
Cb_11_73 bit_11_73 gnd C_bl
Cbb_11_73 bitb_11_73 gnd C_bl
Rb_11_74 bit_11_74 bit_11_75 R_bl
Rbb_11_74 bitb_11_74 bitb_11_75 R_bl
Cb_11_74 bit_11_74 gnd C_bl
Cbb_11_74 bitb_11_74 gnd C_bl
Rb_11_75 bit_11_75 bit_11_76 R_bl
Rbb_11_75 bitb_11_75 bitb_11_76 R_bl
Cb_11_75 bit_11_75 gnd C_bl
Cbb_11_75 bitb_11_75 gnd C_bl
Rb_11_76 bit_11_76 bit_11_77 R_bl
Rbb_11_76 bitb_11_76 bitb_11_77 R_bl
Cb_11_76 bit_11_76 gnd C_bl
Cbb_11_76 bitb_11_76 gnd C_bl
Rb_11_77 bit_11_77 bit_11_78 R_bl
Rbb_11_77 bitb_11_77 bitb_11_78 R_bl
Cb_11_77 bit_11_77 gnd C_bl
Cbb_11_77 bitb_11_77 gnd C_bl
Rb_11_78 bit_11_78 bit_11_79 R_bl
Rbb_11_78 bitb_11_78 bitb_11_79 R_bl
Cb_11_78 bit_11_78 gnd C_bl
Cbb_11_78 bitb_11_78 gnd C_bl
Rb_11_79 bit_11_79 bit_11_80 R_bl
Rbb_11_79 bitb_11_79 bitb_11_80 R_bl
Cb_11_79 bit_11_79 gnd C_bl
Cbb_11_79 bitb_11_79 gnd C_bl
Rb_11_80 bit_11_80 bit_11_81 R_bl
Rbb_11_80 bitb_11_80 bitb_11_81 R_bl
Cb_11_80 bit_11_80 gnd C_bl
Cbb_11_80 bitb_11_80 gnd C_bl
Rb_11_81 bit_11_81 bit_11_82 R_bl
Rbb_11_81 bitb_11_81 bitb_11_82 R_bl
Cb_11_81 bit_11_81 gnd C_bl
Cbb_11_81 bitb_11_81 gnd C_bl
Rb_11_82 bit_11_82 bit_11_83 R_bl
Rbb_11_82 bitb_11_82 bitb_11_83 R_bl
Cb_11_82 bit_11_82 gnd C_bl
Cbb_11_82 bitb_11_82 gnd C_bl
Rb_11_83 bit_11_83 bit_11_84 R_bl
Rbb_11_83 bitb_11_83 bitb_11_84 R_bl
Cb_11_83 bit_11_83 gnd C_bl
Cbb_11_83 bitb_11_83 gnd C_bl
Rb_11_84 bit_11_84 bit_11_85 R_bl
Rbb_11_84 bitb_11_84 bitb_11_85 R_bl
Cb_11_84 bit_11_84 gnd C_bl
Cbb_11_84 bitb_11_84 gnd C_bl
Rb_11_85 bit_11_85 bit_11_86 R_bl
Rbb_11_85 bitb_11_85 bitb_11_86 R_bl
Cb_11_85 bit_11_85 gnd C_bl
Cbb_11_85 bitb_11_85 gnd C_bl
Rb_11_86 bit_11_86 bit_11_87 R_bl
Rbb_11_86 bitb_11_86 bitb_11_87 R_bl
Cb_11_86 bit_11_86 gnd C_bl
Cbb_11_86 bitb_11_86 gnd C_bl
Rb_11_87 bit_11_87 bit_11_88 R_bl
Rbb_11_87 bitb_11_87 bitb_11_88 R_bl
Cb_11_87 bit_11_87 gnd C_bl
Cbb_11_87 bitb_11_87 gnd C_bl
Rb_11_88 bit_11_88 bit_11_89 R_bl
Rbb_11_88 bitb_11_88 bitb_11_89 R_bl
Cb_11_88 bit_11_88 gnd C_bl
Cbb_11_88 bitb_11_88 gnd C_bl
Rb_11_89 bit_11_89 bit_11_90 R_bl
Rbb_11_89 bitb_11_89 bitb_11_90 R_bl
Cb_11_89 bit_11_89 gnd C_bl
Cbb_11_89 bitb_11_89 gnd C_bl
Rb_11_90 bit_11_90 bit_11_91 R_bl
Rbb_11_90 bitb_11_90 bitb_11_91 R_bl
Cb_11_90 bit_11_90 gnd C_bl
Cbb_11_90 bitb_11_90 gnd C_bl
Rb_11_91 bit_11_91 bit_11_92 R_bl
Rbb_11_91 bitb_11_91 bitb_11_92 R_bl
Cb_11_91 bit_11_91 gnd C_bl
Cbb_11_91 bitb_11_91 gnd C_bl
Rb_11_92 bit_11_92 bit_11_93 R_bl
Rbb_11_92 bitb_11_92 bitb_11_93 R_bl
Cb_11_92 bit_11_92 gnd C_bl
Cbb_11_92 bitb_11_92 gnd C_bl
Rb_11_93 bit_11_93 bit_11_94 R_bl
Rbb_11_93 bitb_11_93 bitb_11_94 R_bl
Cb_11_93 bit_11_93 gnd C_bl
Cbb_11_93 bitb_11_93 gnd C_bl
Rb_11_94 bit_11_94 bit_11_95 R_bl
Rbb_11_94 bitb_11_94 bitb_11_95 R_bl
Cb_11_94 bit_11_94 gnd C_bl
Cbb_11_94 bitb_11_94 gnd C_bl
Rb_11_95 bit_11_95 bit_11_96 R_bl
Rbb_11_95 bitb_11_95 bitb_11_96 R_bl
Cb_11_95 bit_11_95 gnd C_bl
Cbb_11_95 bitb_11_95 gnd C_bl
Rb_11_96 bit_11_96 bit_11_97 R_bl
Rbb_11_96 bitb_11_96 bitb_11_97 R_bl
Cb_11_96 bit_11_96 gnd C_bl
Cbb_11_96 bitb_11_96 gnd C_bl
Rb_11_97 bit_11_97 bit_11_98 R_bl
Rbb_11_97 bitb_11_97 bitb_11_98 R_bl
Cb_11_97 bit_11_97 gnd C_bl
Cbb_11_97 bitb_11_97 gnd C_bl
Rb_11_98 bit_11_98 bit_11_99 R_bl
Rbb_11_98 bitb_11_98 bitb_11_99 R_bl
Cb_11_98 bit_11_98 gnd C_bl
Cbb_11_98 bitb_11_98 gnd C_bl
Rb_11_99 bit_11_99 bit_11_100 R_bl
Rbb_11_99 bitb_11_99 bitb_11_100 R_bl
Cb_11_99 bit_11_99 gnd C_bl
Cbb_11_99 bitb_11_99 gnd C_bl
Rb_12_0 bit_12_0 bit_12_1 R_bl
Rbb_12_0 bitb_12_0 bitb_12_1 R_bl
Cb_12_0 bit_12_0 gnd C_bl
Cbb_12_0 bitb_12_0 gnd C_bl
Rb_12_1 bit_12_1 bit_12_2 R_bl
Rbb_12_1 bitb_12_1 bitb_12_2 R_bl
Cb_12_1 bit_12_1 gnd C_bl
Cbb_12_1 bitb_12_1 gnd C_bl
Rb_12_2 bit_12_2 bit_12_3 R_bl
Rbb_12_2 bitb_12_2 bitb_12_3 R_bl
Cb_12_2 bit_12_2 gnd C_bl
Cbb_12_2 bitb_12_2 gnd C_bl
Rb_12_3 bit_12_3 bit_12_4 R_bl
Rbb_12_3 bitb_12_3 bitb_12_4 R_bl
Cb_12_3 bit_12_3 gnd C_bl
Cbb_12_3 bitb_12_3 gnd C_bl
Rb_12_4 bit_12_4 bit_12_5 R_bl
Rbb_12_4 bitb_12_4 bitb_12_5 R_bl
Cb_12_4 bit_12_4 gnd C_bl
Cbb_12_4 bitb_12_4 gnd C_bl
Rb_12_5 bit_12_5 bit_12_6 R_bl
Rbb_12_5 bitb_12_5 bitb_12_6 R_bl
Cb_12_5 bit_12_5 gnd C_bl
Cbb_12_5 bitb_12_5 gnd C_bl
Rb_12_6 bit_12_6 bit_12_7 R_bl
Rbb_12_6 bitb_12_6 bitb_12_7 R_bl
Cb_12_6 bit_12_6 gnd C_bl
Cbb_12_6 bitb_12_6 gnd C_bl
Rb_12_7 bit_12_7 bit_12_8 R_bl
Rbb_12_7 bitb_12_7 bitb_12_8 R_bl
Cb_12_7 bit_12_7 gnd C_bl
Cbb_12_7 bitb_12_7 gnd C_bl
Rb_12_8 bit_12_8 bit_12_9 R_bl
Rbb_12_8 bitb_12_8 bitb_12_9 R_bl
Cb_12_8 bit_12_8 gnd C_bl
Cbb_12_8 bitb_12_8 gnd C_bl
Rb_12_9 bit_12_9 bit_12_10 R_bl
Rbb_12_9 bitb_12_9 bitb_12_10 R_bl
Cb_12_9 bit_12_9 gnd C_bl
Cbb_12_9 bitb_12_9 gnd C_bl
Rb_12_10 bit_12_10 bit_12_11 R_bl
Rbb_12_10 bitb_12_10 bitb_12_11 R_bl
Cb_12_10 bit_12_10 gnd C_bl
Cbb_12_10 bitb_12_10 gnd C_bl
Rb_12_11 bit_12_11 bit_12_12 R_bl
Rbb_12_11 bitb_12_11 bitb_12_12 R_bl
Cb_12_11 bit_12_11 gnd C_bl
Cbb_12_11 bitb_12_11 gnd C_bl
Rb_12_12 bit_12_12 bit_12_13 R_bl
Rbb_12_12 bitb_12_12 bitb_12_13 R_bl
Cb_12_12 bit_12_12 gnd C_bl
Cbb_12_12 bitb_12_12 gnd C_bl
Rb_12_13 bit_12_13 bit_12_14 R_bl
Rbb_12_13 bitb_12_13 bitb_12_14 R_bl
Cb_12_13 bit_12_13 gnd C_bl
Cbb_12_13 bitb_12_13 gnd C_bl
Rb_12_14 bit_12_14 bit_12_15 R_bl
Rbb_12_14 bitb_12_14 bitb_12_15 R_bl
Cb_12_14 bit_12_14 gnd C_bl
Cbb_12_14 bitb_12_14 gnd C_bl
Rb_12_15 bit_12_15 bit_12_16 R_bl
Rbb_12_15 bitb_12_15 bitb_12_16 R_bl
Cb_12_15 bit_12_15 gnd C_bl
Cbb_12_15 bitb_12_15 gnd C_bl
Rb_12_16 bit_12_16 bit_12_17 R_bl
Rbb_12_16 bitb_12_16 bitb_12_17 R_bl
Cb_12_16 bit_12_16 gnd C_bl
Cbb_12_16 bitb_12_16 gnd C_bl
Rb_12_17 bit_12_17 bit_12_18 R_bl
Rbb_12_17 bitb_12_17 bitb_12_18 R_bl
Cb_12_17 bit_12_17 gnd C_bl
Cbb_12_17 bitb_12_17 gnd C_bl
Rb_12_18 bit_12_18 bit_12_19 R_bl
Rbb_12_18 bitb_12_18 bitb_12_19 R_bl
Cb_12_18 bit_12_18 gnd C_bl
Cbb_12_18 bitb_12_18 gnd C_bl
Rb_12_19 bit_12_19 bit_12_20 R_bl
Rbb_12_19 bitb_12_19 bitb_12_20 R_bl
Cb_12_19 bit_12_19 gnd C_bl
Cbb_12_19 bitb_12_19 gnd C_bl
Rb_12_20 bit_12_20 bit_12_21 R_bl
Rbb_12_20 bitb_12_20 bitb_12_21 R_bl
Cb_12_20 bit_12_20 gnd C_bl
Cbb_12_20 bitb_12_20 gnd C_bl
Rb_12_21 bit_12_21 bit_12_22 R_bl
Rbb_12_21 bitb_12_21 bitb_12_22 R_bl
Cb_12_21 bit_12_21 gnd C_bl
Cbb_12_21 bitb_12_21 gnd C_bl
Rb_12_22 bit_12_22 bit_12_23 R_bl
Rbb_12_22 bitb_12_22 bitb_12_23 R_bl
Cb_12_22 bit_12_22 gnd C_bl
Cbb_12_22 bitb_12_22 gnd C_bl
Rb_12_23 bit_12_23 bit_12_24 R_bl
Rbb_12_23 bitb_12_23 bitb_12_24 R_bl
Cb_12_23 bit_12_23 gnd C_bl
Cbb_12_23 bitb_12_23 gnd C_bl
Rb_12_24 bit_12_24 bit_12_25 R_bl
Rbb_12_24 bitb_12_24 bitb_12_25 R_bl
Cb_12_24 bit_12_24 gnd C_bl
Cbb_12_24 bitb_12_24 gnd C_bl
Rb_12_25 bit_12_25 bit_12_26 R_bl
Rbb_12_25 bitb_12_25 bitb_12_26 R_bl
Cb_12_25 bit_12_25 gnd C_bl
Cbb_12_25 bitb_12_25 gnd C_bl
Rb_12_26 bit_12_26 bit_12_27 R_bl
Rbb_12_26 bitb_12_26 bitb_12_27 R_bl
Cb_12_26 bit_12_26 gnd C_bl
Cbb_12_26 bitb_12_26 gnd C_bl
Rb_12_27 bit_12_27 bit_12_28 R_bl
Rbb_12_27 bitb_12_27 bitb_12_28 R_bl
Cb_12_27 bit_12_27 gnd C_bl
Cbb_12_27 bitb_12_27 gnd C_bl
Rb_12_28 bit_12_28 bit_12_29 R_bl
Rbb_12_28 bitb_12_28 bitb_12_29 R_bl
Cb_12_28 bit_12_28 gnd C_bl
Cbb_12_28 bitb_12_28 gnd C_bl
Rb_12_29 bit_12_29 bit_12_30 R_bl
Rbb_12_29 bitb_12_29 bitb_12_30 R_bl
Cb_12_29 bit_12_29 gnd C_bl
Cbb_12_29 bitb_12_29 gnd C_bl
Rb_12_30 bit_12_30 bit_12_31 R_bl
Rbb_12_30 bitb_12_30 bitb_12_31 R_bl
Cb_12_30 bit_12_30 gnd C_bl
Cbb_12_30 bitb_12_30 gnd C_bl
Rb_12_31 bit_12_31 bit_12_32 R_bl
Rbb_12_31 bitb_12_31 bitb_12_32 R_bl
Cb_12_31 bit_12_31 gnd C_bl
Cbb_12_31 bitb_12_31 gnd C_bl
Rb_12_32 bit_12_32 bit_12_33 R_bl
Rbb_12_32 bitb_12_32 bitb_12_33 R_bl
Cb_12_32 bit_12_32 gnd C_bl
Cbb_12_32 bitb_12_32 gnd C_bl
Rb_12_33 bit_12_33 bit_12_34 R_bl
Rbb_12_33 bitb_12_33 bitb_12_34 R_bl
Cb_12_33 bit_12_33 gnd C_bl
Cbb_12_33 bitb_12_33 gnd C_bl
Rb_12_34 bit_12_34 bit_12_35 R_bl
Rbb_12_34 bitb_12_34 bitb_12_35 R_bl
Cb_12_34 bit_12_34 gnd C_bl
Cbb_12_34 bitb_12_34 gnd C_bl
Rb_12_35 bit_12_35 bit_12_36 R_bl
Rbb_12_35 bitb_12_35 bitb_12_36 R_bl
Cb_12_35 bit_12_35 gnd C_bl
Cbb_12_35 bitb_12_35 gnd C_bl
Rb_12_36 bit_12_36 bit_12_37 R_bl
Rbb_12_36 bitb_12_36 bitb_12_37 R_bl
Cb_12_36 bit_12_36 gnd C_bl
Cbb_12_36 bitb_12_36 gnd C_bl
Rb_12_37 bit_12_37 bit_12_38 R_bl
Rbb_12_37 bitb_12_37 bitb_12_38 R_bl
Cb_12_37 bit_12_37 gnd C_bl
Cbb_12_37 bitb_12_37 gnd C_bl
Rb_12_38 bit_12_38 bit_12_39 R_bl
Rbb_12_38 bitb_12_38 bitb_12_39 R_bl
Cb_12_38 bit_12_38 gnd C_bl
Cbb_12_38 bitb_12_38 gnd C_bl
Rb_12_39 bit_12_39 bit_12_40 R_bl
Rbb_12_39 bitb_12_39 bitb_12_40 R_bl
Cb_12_39 bit_12_39 gnd C_bl
Cbb_12_39 bitb_12_39 gnd C_bl
Rb_12_40 bit_12_40 bit_12_41 R_bl
Rbb_12_40 bitb_12_40 bitb_12_41 R_bl
Cb_12_40 bit_12_40 gnd C_bl
Cbb_12_40 bitb_12_40 gnd C_bl
Rb_12_41 bit_12_41 bit_12_42 R_bl
Rbb_12_41 bitb_12_41 bitb_12_42 R_bl
Cb_12_41 bit_12_41 gnd C_bl
Cbb_12_41 bitb_12_41 gnd C_bl
Rb_12_42 bit_12_42 bit_12_43 R_bl
Rbb_12_42 bitb_12_42 bitb_12_43 R_bl
Cb_12_42 bit_12_42 gnd C_bl
Cbb_12_42 bitb_12_42 gnd C_bl
Rb_12_43 bit_12_43 bit_12_44 R_bl
Rbb_12_43 bitb_12_43 bitb_12_44 R_bl
Cb_12_43 bit_12_43 gnd C_bl
Cbb_12_43 bitb_12_43 gnd C_bl
Rb_12_44 bit_12_44 bit_12_45 R_bl
Rbb_12_44 bitb_12_44 bitb_12_45 R_bl
Cb_12_44 bit_12_44 gnd C_bl
Cbb_12_44 bitb_12_44 gnd C_bl
Rb_12_45 bit_12_45 bit_12_46 R_bl
Rbb_12_45 bitb_12_45 bitb_12_46 R_bl
Cb_12_45 bit_12_45 gnd C_bl
Cbb_12_45 bitb_12_45 gnd C_bl
Rb_12_46 bit_12_46 bit_12_47 R_bl
Rbb_12_46 bitb_12_46 bitb_12_47 R_bl
Cb_12_46 bit_12_46 gnd C_bl
Cbb_12_46 bitb_12_46 gnd C_bl
Rb_12_47 bit_12_47 bit_12_48 R_bl
Rbb_12_47 bitb_12_47 bitb_12_48 R_bl
Cb_12_47 bit_12_47 gnd C_bl
Cbb_12_47 bitb_12_47 gnd C_bl
Rb_12_48 bit_12_48 bit_12_49 R_bl
Rbb_12_48 bitb_12_48 bitb_12_49 R_bl
Cb_12_48 bit_12_48 gnd C_bl
Cbb_12_48 bitb_12_48 gnd C_bl
Rb_12_49 bit_12_49 bit_12_50 R_bl
Rbb_12_49 bitb_12_49 bitb_12_50 R_bl
Cb_12_49 bit_12_49 gnd C_bl
Cbb_12_49 bitb_12_49 gnd C_bl
Rb_12_50 bit_12_50 bit_12_51 R_bl
Rbb_12_50 bitb_12_50 bitb_12_51 R_bl
Cb_12_50 bit_12_50 gnd C_bl
Cbb_12_50 bitb_12_50 gnd C_bl
Rb_12_51 bit_12_51 bit_12_52 R_bl
Rbb_12_51 bitb_12_51 bitb_12_52 R_bl
Cb_12_51 bit_12_51 gnd C_bl
Cbb_12_51 bitb_12_51 gnd C_bl
Rb_12_52 bit_12_52 bit_12_53 R_bl
Rbb_12_52 bitb_12_52 bitb_12_53 R_bl
Cb_12_52 bit_12_52 gnd C_bl
Cbb_12_52 bitb_12_52 gnd C_bl
Rb_12_53 bit_12_53 bit_12_54 R_bl
Rbb_12_53 bitb_12_53 bitb_12_54 R_bl
Cb_12_53 bit_12_53 gnd C_bl
Cbb_12_53 bitb_12_53 gnd C_bl
Rb_12_54 bit_12_54 bit_12_55 R_bl
Rbb_12_54 bitb_12_54 bitb_12_55 R_bl
Cb_12_54 bit_12_54 gnd C_bl
Cbb_12_54 bitb_12_54 gnd C_bl
Rb_12_55 bit_12_55 bit_12_56 R_bl
Rbb_12_55 bitb_12_55 bitb_12_56 R_bl
Cb_12_55 bit_12_55 gnd C_bl
Cbb_12_55 bitb_12_55 gnd C_bl
Rb_12_56 bit_12_56 bit_12_57 R_bl
Rbb_12_56 bitb_12_56 bitb_12_57 R_bl
Cb_12_56 bit_12_56 gnd C_bl
Cbb_12_56 bitb_12_56 gnd C_bl
Rb_12_57 bit_12_57 bit_12_58 R_bl
Rbb_12_57 bitb_12_57 bitb_12_58 R_bl
Cb_12_57 bit_12_57 gnd C_bl
Cbb_12_57 bitb_12_57 gnd C_bl
Rb_12_58 bit_12_58 bit_12_59 R_bl
Rbb_12_58 bitb_12_58 bitb_12_59 R_bl
Cb_12_58 bit_12_58 gnd C_bl
Cbb_12_58 bitb_12_58 gnd C_bl
Rb_12_59 bit_12_59 bit_12_60 R_bl
Rbb_12_59 bitb_12_59 bitb_12_60 R_bl
Cb_12_59 bit_12_59 gnd C_bl
Cbb_12_59 bitb_12_59 gnd C_bl
Rb_12_60 bit_12_60 bit_12_61 R_bl
Rbb_12_60 bitb_12_60 bitb_12_61 R_bl
Cb_12_60 bit_12_60 gnd C_bl
Cbb_12_60 bitb_12_60 gnd C_bl
Rb_12_61 bit_12_61 bit_12_62 R_bl
Rbb_12_61 bitb_12_61 bitb_12_62 R_bl
Cb_12_61 bit_12_61 gnd C_bl
Cbb_12_61 bitb_12_61 gnd C_bl
Rb_12_62 bit_12_62 bit_12_63 R_bl
Rbb_12_62 bitb_12_62 bitb_12_63 R_bl
Cb_12_62 bit_12_62 gnd C_bl
Cbb_12_62 bitb_12_62 gnd C_bl
Rb_12_63 bit_12_63 bit_12_64 R_bl
Rbb_12_63 bitb_12_63 bitb_12_64 R_bl
Cb_12_63 bit_12_63 gnd C_bl
Cbb_12_63 bitb_12_63 gnd C_bl
Rb_12_64 bit_12_64 bit_12_65 R_bl
Rbb_12_64 bitb_12_64 bitb_12_65 R_bl
Cb_12_64 bit_12_64 gnd C_bl
Cbb_12_64 bitb_12_64 gnd C_bl
Rb_12_65 bit_12_65 bit_12_66 R_bl
Rbb_12_65 bitb_12_65 bitb_12_66 R_bl
Cb_12_65 bit_12_65 gnd C_bl
Cbb_12_65 bitb_12_65 gnd C_bl
Rb_12_66 bit_12_66 bit_12_67 R_bl
Rbb_12_66 bitb_12_66 bitb_12_67 R_bl
Cb_12_66 bit_12_66 gnd C_bl
Cbb_12_66 bitb_12_66 gnd C_bl
Rb_12_67 bit_12_67 bit_12_68 R_bl
Rbb_12_67 bitb_12_67 bitb_12_68 R_bl
Cb_12_67 bit_12_67 gnd C_bl
Cbb_12_67 bitb_12_67 gnd C_bl
Rb_12_68 bit_12_68 bit_12_69 R_bl
Rbb_12_68 bitb_12_68 bitb_12_69 R_bl
Cb_12_68 bit_12_68 gnd C_bl
Cbb_12_68 bitb_12_68 gnd C_bl
Rb_12_69 bit_12_69 bit_12_70 R_bl
Rbb_12_69 bitb_12_69 bitb_12_70 R_bl
Cb_12_69 bit_12_69 gnd C_bl
Cbb_12_69 bitb_12_69 gnd C_bl
Rb_12_70 bit_12_70 bit_12_71 R_bl
Rbb_12_70 bitb_12_70 bitb_12_71 R_bl
Cb_12_70 bit_12_70 gnd C_bl
Cbb_12_70 bitb_12_70 gnd C_bl
Rb_12_71 bit_12_71 bit_12_72 R_bl
Rbb_12_71 bitb_12_71 bitb_12_72 R_bl
Cb_12_71 bit_12_71 gnd C_bl
Cbb_12_71 bitb_12_71 gnd C_bl
Rb_12_72 bit_12_72 bit_12_73 R_bl
Rbb_12_72 bitb_12_72 bitb_12_73 R_bl
Cb_12_72 bit_12_72 gnd C_bl
Cbb_12_72 bitb_12_72 gnd C_bl
Rb_12_73 bit_12_73 bit_12_74 R_bl
Rbb_12_73 bitb_12_73 bitb_12_74 R_bl
Cb_12_73 bit_12_73 gnd C_bl
Cbb_12_73 bitb_12_73 gnd C_bl
Rb_12_74 bit_12_74 bit_12_75 R_bl
Rbb_12_74 bitb_12_74 bitb_12_75 R_bl
Cb_12_74 bit_12_74 gnd C_bl
Cbb_12_74 bitb_12_74 gnd C_bl
Rb_12_75 bit_12_75 bit_12_76 R_bl
Rbb_12_75 bitb_12_75 bitb_12_76 R_bl
Cb_12_75 bit_12_75 gnd C_bl
Cbb_12_75 bitb_12_75 gnd C_bl
Rb_12_76 bit_12_76 bit_12_77 R_bl
Rbb_12_76 bitb_12_76 bitb_12_77 R_bl
Cb_12_76 bit_12_76 gnd C_bl
Cbb_12_76 bitb_12_76 gnd C_bl
Rb_12_77 bit_12_77 bit_12_78 R_bl
Rbb_12_77 bitb_12_77 bitb_12_78 R_bl
Cb_12_77 bit_12_77 gnd C_bl
Cbb_12_77 bitb_12_77 gnd C_bl
Rb_12_78 bit_12_78 bit_12_79 R_bl
Rbb_12_78 bitb_12_78 bitb_12_79 R_bl
Cb_12_78 bit_12_78 gnd C_bl
Cbb_12_78 bitb_12_78 gnd C_bl
Rb_12_79 bit_12_79 bit_12_80 R_bl
Rbb_12_79 bitb_12_79 bitb_12_80 R_bl
Cb_12_79 bit_12_79 gnd C_bl
Cbb_12_79 bitb_12_79 gnd C_bl
Rb_12_80 bit_12_80 bit_12_81 R_bl
Rbb_12_80 bitb_12_80 bitb_12_81 R_bl
Cb_12_80 bit_12_80 gnd C_bl
Cbb_12_80 bitb_12_80 gnd C_bl
Rb_12_81 bit_12_81 bit_12_82 R_bl
Rbb_12_81 bitb_12_81 bitb_12_82 R_bl
Cb_12_81 bit_12_81 gnd C_bl
Cbb_12_81 bitb_12_81 gnd C_bl
Rb_12_82 bit_12_82 bit_12_83 R_bl
Rbb_12_82 bitb_12_82 bitb_12_83 R_bl
Cb_12_82 bit_12_82 gnd C_bl
Cbb_12_82 bitb_12_82 gnd C_bl
Rb_12_83 bit_12_83 bit_12_84 R_bl
Rbb_12_83 bitb_12_83 bitb_12_84 R_bl
Cb_12_83 bit_12_83 gnd C_bl
Cbb_12_83 bitb_12_83 gnd C_bl
Rb_12_84 bit_12_84 bit_12_85 R_bl
Rbb_12_84 bitb_12_84 bitb_12_85 R_bl
Cb_12_84 bit_12_84 gnd C_bl
Cbb_12_84 bitb_12_84 gnd C_bl
Rb_12_85 bit_12_85 bit_12_86 R_bl
Rbb_12_85 bitb_12_85 bitb_12_86 R_bl
Cb_12_85 bit_12_85 gnd C_bl
Cbb_12_85 bitb_12_85 gnd C_bl
Rb_12_86 bit_12_86 bit_12_87 R_bl
Rbb_12_86 bitb_12_86 bitb_12_87 R_bl
Cb_12_86 bit_12_86 gnd C_bl
Cbb_12_86 bitb_12_86 gnd C_bl
Rb_12_87 bit_12_87 bit_12_88 R_bl
Rbb_12_87 bitb_12_87 bitb_12_88 R_bl
Cb_12_87 bit_12_87 gnd C_bl
Cbb_12_87 bitb_12_87 gnd C_bl
Rb_12_88 bit_12_88 bit_12_89 R_bl
Rbb_12_88 bitb_12_88 bitb_12_89 R_bl
Cb_12_88 bit_12_88 gnd C_bl
Cbb_12_88 bitb_12_88 gnd C_bl
Rb_12_89 bit_12_89 bit_12_90 R_bl
Rbb_12_89 bitb_12_89 bitb_12_90 R_bl
Cb_12_89 bit_12_89 gnd C_bl
Cbb_12_89 bitb_12_89 gnd C_bl
Rb_12_90 bit_12_90 bit_12_91 R_bl
Rbb_12_90 bitb_12_90 bitb_12_91 R_bl
Cb_12_90 bit_12_90 gnd C_bl
Cbb_12_90 bitb_12_90 gnd C_bl
Rb_12_91 bit_12_91 bit_12_92 R_bl
Rbb_12_91 bitb_12_91 bitb_12_92 R_bl
Cb_12_91 bit_12_91 gnd C_bl
Cbb_12_91 bitb_12_91 gnd C_bl
Rb_12_92 bit_12_92 bit_12_93 R_bl
Rbb_12_92 bitb_12_92 bitb_12_93 R_bl
Cb_12_92 bit_12_92 gnd C_bl
Cbb_12_92 bitb_12_92 gnd C_bl
Rb_12_93 bit_12_93 bit_12_94 R_bl
Rbb_12_93 bitb_12_93 bitb_12_94 R_bl
Cb_12_93 bit_12_93 gnd C_bl
Cbb_12_93 bitb_12_93 gnd C_bl
Rb_12_94 bit_12_94 bit_12_95 R_bl
Rbb_12_94 bitb_12_94 bitb_12_95 R_bl
Cb_12_94 bit_12_94 gnd C_bl
Cbb_12_94 bitb_12_94 gnd C_bl
Rb_12_95 bit_12_95 bit_12_96 R_bl
Rbb_12_95 bitb_12_95 bitb_12_96 R_bl
Cb_12_95 bit_12_95 gnd C_bl
Cbb_12_95 bitb_12_95 gnd C_bl
Rb_12_96 bit_12_96 bit_12_97 R_bl
Rbb_12_96 bitb_12_96 bitb_12_97 R_bl
Cb_12_96 bit_12_96 gnd C_bl
Cbb_12_96 bitb_12_96 gnd C_bl
Rb_12_97 bit_12_97 bit_12_98 R_bl
Rbb_12_97 bitb_12_97 bitb_12_98 R_bl
Cb_12_97 bit_12_97 gnd C_bl
Cbb_12_97 bitb_12_97 gnd C_bl
Rb_12_98 bit_12_98 bit_12_99 R_bl
Rbb_12_98 bitb_12_98 bitb_12_99 R_bl
Cb_12_98 bit_12_98 gnd C_bl
Cbb_12_98 bitb_12_98 gnd C_bl
Rb_12_99 bit_12_99 bit_12_100 R_bl
Rbb_12_99 bitb_12_99 bitb_12_100 R_bl
Cb_12_99 bit_12_99 gnd C_bl
Cbb_12_99 bitb_12_99 gnd C_bl
Rb_13_0 bit_13_0 bit_13_1 R_bl
Rbb_13_0 bitb_13_0 bitb_13_1 R_bl
Cb_13_0 bit_13_0 gnd C_bl
Cbb_13_0 bitb_13_0 gnd C_bl
Rb_13_1 bit_13_1 bit_13_2 R_bl
Rbb_13_1 bitb_13_1 bitb_13_2 R_bl
Cb_13_1 bit_13_1 gnd C_bl
Cbb_13_1 bitb_13_1 gnd C_bl
Rb_13_2 bit_13_2 bit_13_3 R_bl
Rbb_13_2 bitb_13_2 bitb_13_3 R_bl
Cb_13_2 bit_13_2 gnd C_bl
Cbb_13_2 bitb_13_2 gnd C_bl
Rb_13_3 bit_13_3 bit_13_4 R_bl
Rbb_13_3 bitb_13_3 bitb_13_4 R_bl
Cb_13_3 bit_13_3 gnd C_bl
Cbb_13_3 bitb_13_3 gnd C_bl
Rb_13_4 bit_13_4 bit_13_5 R_bl
Rbb_13_4 bitb_13_4 bitb_13_5 R_bl
Cb_13_4 bit_13_4 gnd C_bl
Cbb_13_4 bitb_13_4 gnd C_bl
Rb_13_5 bit_13_5 bit_13_6 R_bl
Rbb_13_5 bitb_13_5 bitb_13_6 R_bl
Cb_13_5 bit_13_5 gnd C_bl
Cbb_13_5 bitb_13_5 gnd C_bl
Rb_13_6 bit_13_6 bit_13_7 R_bl
Rbb_13_6 bitb_13_6 bitb_13_7 R_bl
Cb_13_6 bit_13_6 gnd C_bl
Cbb_13_6 bitb_13_6 gnd C_bl
Rb_13_7 bit_13_7 bit_13_8 R_bl
Rbb_13_7 bitb_13_7 bitb_13_8 R_bl
Cb_13_7 bit_13_7 gnd C_bl
Cbb_13_7 bitb_13_7 gnd C_bl
Rb_13_8 bit_13_8 bit_13_9 R_bl
Rbb_13_8 bitb_13_8 bitb_13_9 R_bl
Cb_13_8 bit_13_8 gnd C_bl
Cbb_13_8 bitb_13_8 gnd C_bl
Rb_13_9 bit_13_9 bit_13_10 R_bl
Rbb_13_9 bitb_13_9 bitb_13_10 R_bl
Cb_13_9 bit_13_9 gnd C_bl
Cbb_13_9 bitb_13_9 gnd C_bl
Rb_13_10 bit_13_10 bit_13_11 R_bl
Rbb_13_10 bitb_13_10 bitb_13_11 R_bl
Cb_13_10 bit_13_10 gnd C_bl
Cbb_13_10 bitb_13_10 gnd C_bl
Rb_13_11 bit_13_11 bit_13_12 R_bl
Rbb_13_11 bitb_13_11 bitb_13_12 R_bl
Cb_13_11 bit_13_11 gnd C_bl
Cbb_13_11 bitb_13_11 gnd C_bl
Rb_13_12 bit_13_12 bit_13_13 R_bl
Rbb_13_12 bitb_13_12 bitb_13_13 R_bl
Cb_13_12 bit_13_12 gnd C_bl
Cbb_13_12 bitb_13_12 gnd C_bl
Rb_13_13 bit_13_13 bit_13_14 R_bl
Rbb_13_13 bitb_13_13 bitb_13_14 R_bl
Cb_13_13 bit_13_13 gnd C_bl
Cbb_13_13 bitb_13_13 gnd C_bl
Rb_13_14 bit_13_14 bit_13_15 R_bl
Rbb_13_14 bitb_13_14 bitb_13_15 R_bl
Cb_13_14 bit_13_14 gnd C_bl
Cbb_13_14 bitb_13_14 gnd C_bl
Rb_13_15 bit_13_15 bit_13_16 R_bl
Rbb_13_15 bitb_13_15 bitb_13_16 R_bl
Cb_13_15 bit_13_15 gnd C_bl
Cbb_13_15 bitb_13_15 gnd C_bl
Rb_13_16 bit_13_16 bit_13_17 R_bl
Rbb_13_16 bitb_13_16 bitb_13_17 R_bl
Cb_13_16 bit_13_16 gnd C_bl
Cbb_13_16 bitb_13_16 gnd C_bl
Rb_13_17 bit_13_17 bit_13_18 R_bl
Rbb_13_17 bitb_13_17 bitb_13_18 R_bl
Cb_13_17 bit_13_17 gnd C_bl
Cbb_13_17 bitb_13_17 gnd C_bl
Rb_13_18 bit_13_18 bit_13_19 R_bl
Rbb_13_18 bitb_13_18 bitb_13_19 R_bl
Cb_13_18 bit_13_18 gnd C_bl
Cbb_13_18 bitb_13_18 gnd C_bl
Rb_13_19 bit_13_19 bit_13_20 R_bl
Rbb_13_19 bitb_13_19 bitb_13_20 R_bl
Cb_13_19 bit_13_19 gnd C_bl
Cbb_13_19 bitb_13_19 gnd C_bl
Rb_13_20 bit_13_20 bit_13_21 R_bl
Rbb_13_20 bitb_13_20 bitb_13_21 R_bl
Cb_13_20 bit_13_20 gnd C_bl
Cbb_13_20 bitb_13_20 gnd C_bl
Rb_13_21 bit_13_21 bit_13_22 R_bl
Rbb_13_21 bitb_13_21 bitb_13_22 R_bl
Cb_13_21 bit_13_21 gnd C_bl
Cbb_13_21 bitb_13_21 gnd C_bl
Rb_13_22 bit_13_22 bit_13_23 R_bl
Rbb_13_22 bitb_13_22 bitb_13_23 R_bl
Cb_13_22 bit_13_22 gnd C_bl
Cbb_13_22 bitb_13_22 gnd C_bl
Rb_13_23 bit_13_23 bit_13_24 R_bl
Rbb_13_23 bitb_13_23 bitb_13_24 R_bl
Cb_13_23 bit_13_23 gnd C_bl
Cbb_13_23 bitb_13_23 gnd C_bl
Rb_13_24 bit_13_24 bit_13_25 R_bl
Rbb_13_24 bitb_13_24 bitb_13_25 R_bl
Cb_13_24 bit_13_24 gnd C_bl
Cbb_13_24 bitb_13_24 gnd C_bl
Rb_13_25 bit_13_25 bit_13_26 R_bl
Rbb_13_25 bitb_13_25 bitb_13_26 R_bl
Cb_13_25 bit_13_25 gnd C_bl
Cbb_13_25 bitb_13_25 gnd C_bl
Rb_13_26 bit_13_26 bit_13_27 R_bl
Rbb_13_26 bitb_13_26 bitb_13_27 R_bl
Cb_13_26 bit_13_26 gnd C_bl
Cbb_13_26 bitb_13_26 gnd C_bl
Rb_13_27 bit_13_27 bit_13_28 R_bl
Rbb_13_27 bitb_13_27 bitb_13_28 R_bl
Cb_13_27 bit_13_27 gnd C_bl
Cbb_13_27 bitb_13_27 gnd C_bl
Rb_13_28 bit_13_28 bit_13_29 R_bl
Rbb_13_28 bitb_13_28 bitb_13_29 R_bl
Cb_13_28 bit_13_28 gnd C_bl
Cbb_13_28 bitb_13_28 gnd C_bl
Rb_13_29 bit_13_29 bit_13_30 R_bl
Rbb_13_29 bitb_13_29 bitb_13_30 R_bl
Cb_13_29 bit_13_29 gnd C_bl
Cbb_13_29 bitb_13_29 gnd C_bl
Rb_13_30 bit_13_30 bit_13_31 R_bl
Rbb_13_30 bitb_13_30 bitb_13_31 R_bl
Cb_13_30 bit_13_30 gnd C_bl
Cbb_13_30 bitb_13_30 gnd C_bl
Rb_13_31 bit_13_31 bit_13_32 R_bl
Rbb_13_31 bitb_13_31 bitb_13_32 R_bl
Cb_13_31 bit_13_31 gnd C_bl
Cbb_13_31 bitb_13_31 gnd C_bl
Rb_13_32 bit_13_32 bit_13_33 R_bl
Rbb_13_32 bitb_13_32 bitb_13_33 R_bl
Cb_13_32 bit_13_32 gnd C_bl
Cbb_13_32 bitb_13_32 gnd C_bl
Rb_13_33 bit_13_33 bit_13_34 R_bl
Rbb_13_33 bitb_13_33 bitb_13_34 R_bl
Cb_13_33 bit_13_33 gnd C_bl
Cbb_13_33 bitb_13_33 gnd C_bl
Rb_13_34 bit_13_34 bit_13_35 R_bl
Rbb_13_34 bitb_13_34 bitb_13_35 R_bl
Cb_13_34 bit_13_34 gnd C_bl
Cbb_13_34 bitb_13_34 gnd C_bl
Rb_13_35 bit_13_35 bit_13_36 R_bl
Rbb_13_35 bitb_13_35 bitb_13_36 R_bl
Cb_13_35 bit_13_35 gnd C_bl
Cbb_13_35 bitb_13_35 gnd C_bl
Rb_13_36 bit_13_36 bit_13_37 R_bl
Rbb_13_36 bitb_13_36 bitb_13_37 R_bl
Cb_13_36 bit_13_36 gnd C_bl
Cbb_13_36 bitb_13_36 gnd C_bl
Rb_13_37 bit_13_37 bit_13_38 R_bl
Rbb_13_37 bitb_13_37 bitb_13_38 R_bl
Cb_13_37 bit_13_37 gnd C_bl
Cbb_13_37 bitb_13_37 gnd C_bl
Rb_13_38 bit_13_38 bit_13_39 R_bl
Rbb_13_38 bitb_13_38 bitb_13_39 R_bl
Cb_13_38 bit_13_38 gnd C_bl
Cbb_13_38 bitb_13_38 gnd C_bl
Rb_13_39 bit_13_39 bit_13_40 R_bl
Rbb_13_39 bitb_13_39 bitb_13_40 R_bl
Cb_13_39 bit_13_39 gnd C_bl
Cbb_13_39 bitb_13_39 gnd C_bl
Rb_13_40 bit_13_40 bit_13_41 R_bl
Rbb_13_40 bitb_13_40 bitb_13_41 R_bl
Cb_13_40 bit_13_40 gnd C_bl
Cbb_13_40 bitb_13_40 gnd C_bl
Rb_13_41 bit_13_41 bit_13_42 R_bl
Rbb_13_41 bitb_13_41 bitb_13_42 R_bl
Cb_13_41 bit_13_41 gnd C_bl
Cbb_13_41 bitb_13_41 gnd C_bl
Rb_13_42 bit_13_42 bit_13_43 R_bl
Rbb_13_42 bitb_13_42 bitb_13_43 R_bl
Cb_13_42 bit_13_42 gnd C_bl
Cbb_13_42 bitb_13_42 gnd C_bl
Rb_13_43 bit_13_43 bit_13_44 R_bl
Rbb_13_43 bitb_13_43 bitb_13_44 R_bl
Cb_13_43 bit_13_43 gnd C_bl
Cbb_13_43 bitb_13_43 gnd C_bl
Rb_13_44 bit_13_44 bit_13_45 R_bl
Rbb_13_44 bitb_13_44 bitb_13_45 R_bl
Cb_13_44 bit_13_44 gnd C_bl
Cbb_13_44 bitb_13_44 gnd C_bl
Rb_13_45 bit_13_45 bit_13_46 R_bl
Rbb_13_45 bitb_13_45 bitb_13_46 R_bl
Cb_13_45 bit_13_45 gnd C_bl
Cbb_13_45 bitb_13_45 gnd C_bl
Rb_13_46 bit_13_46 bit_13_47 R_bl
Rbb_13_46 bitb_13_46 bitb_13_47 R_bl
Cb_13_46 bit_13_46 gnd C_bl
Cbb_13_46 bitb_13_46 gnd C_bl
Rb_13_47 bit_13_47 bit_13_48 R_bl
Rbb_13_47 bitb_13_47 bitb_13_48 R_bl
Cb_13_47 bit_13_47 gnd C_bl
Cbb_13_47 bitb_13_47 gnd C_bl
Rb_13_48 bit_13_48 bit_13_49 R_bl
Rbb_13_48 bitb_13_48 bitb_13_49 R_bl
Cb_13_48 bit_13_48 gnd C_bl
Cbb_13_48 bitb_13_48 gnd C_bl
Rb_13_49 bit_13_49 bit_13_50 R_bl
Rbb_13_49 bitb_13_49 bitb_13_50 R_bl
Cb_13_49 bit_13_49 gnd C_bl
Cbb_13_49 bitb_13_49 gnd C_bl
Rb_13_50 bit_13_50 bit_13_51 R_bl
Rbb_13_50 bitb_13_50 bitb_13_51 R_bl
Cb_13_50 bit_13_50 gnd C_bl
Cbb_13_50 bitb_13_50 gnd C_bl
Rb_13_51 bit_13_51 bit_13_52 R_bl
Rbb_13_51 bitb_13_51 bitb_13_52 R_bl
Cb_13_51 bit_13_51 gnd C_bl
Cbb_13_51 bitb_13_51 gnd C_bl
Rb_13_52 bit_13_52 bit_13_53 R_bl
Rbb_13_52 bitb_13_52 bitb_13_53 R_bl
Cb_13_52 bit_13_52 gnd C_bl
Cbb_13_52 bitb_13_52 gnd C_bl
Rb_13_53 bit_13_53 bit_13_54 R_bl
Rbb_13_53 bitb_13_53 bitb_13_54 R_bl
Cb_13_53 bit_13_53 gnd C_bl
Cbb_13_53 bitb_13_53 gnd C_bl
Rb_13_54 bit_13_54 bit_13_55 R_bl
Rbb_13_54 bitb_13_54 bitb_13_55 R_bl
Cb_13_54 bit_13_54 gnd C_bl
Cbb_13_54 bitb_13_54 gnd C_bl
Rb_13_55 bit_13_55 bit_13_56 R_bl
Rbb_13_55 bitb_13_55 bitb_13_56 R_bl
Cb_13_55 bit_13_55 gnd C_bl
Cbb_13_55 bitb_13_55 gnd C_bl
Rb_13_56 bit_13_56 bit_13_57 R_bl
Rbb_13_56 bitb_13_56 bitb_13_57 R_bl
Cb_13_56 bit_13_56 gnd C_bl
Cbb_13_56 bitb_13_56 gnd C_bl
Rb_13_57 bit_13_57 bit_13_58 R_bl
Rbb_13_57 bitb_13_57 bitb_13_58 R_bl
Cb_13_57 bit_13_57 gnd C_bl
Cbb_13_57 bitb_13_57 gnd C_bl
Rb_13_58 bit_13_58 bit_13_59 R_bl
Rbb_13_58 bitb_13_58 bitb_13_59 R_bl
Cb_13_58 bit_13_58 gnd C_bl
Cbb_13_58 bitb_13_58 gnd C_bl
Rb_13_59 bit_13_59 bit_13_60 R_bl
Rbb_13_59 bitb_13_59 bitb_13_60 R_bl
Cb_13_59 bit_13_59 gnd C_bl
Cbb_13_59 bitb_13_59 gnd C_bl
Rb_13_60 bit_13_60 bit_13_61 R_bl
Rbb_13_60 bitb_13_60 bitb_13_61 R_bl
Cb_13_60 bit_13_60 gnd C_bl
Cbb_13_60 bitb_13_60 gnd C_bl
Rb_13_61 bit_13_61 bit_13_62 R_bl
Rbb_13_61 bitb_13_61 bitb_13_62 R_bl
Cb_13_61 bit_13_61 gnd C_bl
Cbb_13_61 bitb_13_61 gnd C_bl
Rb_13_62 bit_13_62 bit_13_63 R_bl
Rbb_13_62 bitb_13_62 bitb_13_63 R_bl
Cb_13_62 bit_13_62 gnd C_bl
Cbb_13_62 bitb_13_62 gnd C_bl
Rb_13_63 bit_13_63 bit_13_64 R_bl
Rbb_13_63 bitb_13_63 bitb_13_64 R_bl
Cb_13_63 bit_13_63 gnd C_bl
Cbb_13_63 bitb_13_63 gnd C_bl
Rb_13_64 bit_13_64 bit_13_65 R_bl
Rbb_13_64 bitb_13_64 bitb_13_65 R_bl
Cb_13_64 bit_13_64 gnd C_bl
Cbb_13_64 bitb_13_64 gnd C_bl
Rb_13_65 bit_13_65 bit_13_66 R_bl
Rbb_13_65 bitb_13_65 bitb_13_66 R_bl
Cb_13_65 bit_13_65 gnd C_bl
Cbb_13_65 bitb_13_65 gnd C_bl
Rb_13_66 bit_13_66 bit_13_67 R_bl
Rbb_13_66 bitb_13_66 bitb_13_67 R_bl
Cb_13_66 bit_13_66 gnd C_bl
Cbb_13_66 bitb_13_66 gnd C_bl
Rb_13_67 bit_13_67 bit_13_68 R_bl
Rbb_13_67 bitb_13_67 bitb_13_68 R_bl
Cb_13_67 bit_13_67 gnd C_bl
Cbb_13_67 bitb_13_67 gnd C_bl
Rb_13_68 bit_13_68 bit_13_69 R_bl
Rbb_13_68 bitb_13_68 bitb_13_69 R_bl
Cb_13_68 bit_13_68 gnd C_bl
Cbb_13_68 bitb_13_68 gnd C_bl
Rb_13_69 bit_13_69 bit_13_70 R_bl
Rbb_13_69 bitb_13_69 bitb_13_70 R_bl
Cb_13_69 bit_13_69 gnd C_bl
Cbb_13_69 bitb_13_69 gnd C_bl
Rb_13_70 bit_13_70 bit_13_71 R_bl
Rbb_13_70 bitb_13_70 bitb_13_71 R_bl
Cb_13_70 bit_13_70 gnd C_bl
Cbb_13_70 bitb_13_70 gnd C_bl
Rb_13_71 bit_13_71 bit_13_72 R_bl
Rbb_13_71 bitb_13_71 bitb_13_72 R_bl
Cb_13_71 bit_13_71 gnd C_bl
Cbb_13_71 bitb_13_71 gnd C_bl
Rb_13_72 bit_13_72 bit_13_73 R_bl
Rbb_13_72 bitb_13_72 bitb_13_73 R_bl
Cb_13_72 bit_13_72 gnd C_bl
Cbb_13_72 bitb_13_72 gnd C_bl
Rb_13_73 bit_13_73 bit_13_74 R_bl
Rbb_13_73 bitb_13_73 bitb_13_74 R_bl
Cb_13_73 bit_13_73 gnd C_bl
Cbb_13_73 bitb_13_73 gnd C_bl
Rb_13_74 bit_13_74 bit_13_75 R_bl
Rbb_13_74 bitb_13_74 bitb_13_75 R_bl
Cb_13_74 bit_13_74 gnd C_bl
Cbb_13_74 bitb_13_74 gnd C_bl
Rb_13_75 bit_13_75 bit_13_76 R_bl
Rbb_13_75 bitb_13_75 bitb_13_76 R_bl
Cb_13_75 bit_13_75 gnd C_bl
Cbb_13_75 bitb_13_75 gnd C_bl
Rb_13_76 bit_13_76 bit_13_77 R_bl
Rbb_13_76 bitb_13_76 bitb_13_77 R_bl
Cb_13_76 bit_13_76 gnd C_bl
Cbb_13_76 bitb_13_76 gnd C_bl
Rb_13_77 bit_13_77 bit_13_78 R_bl
Rbb_13_77 bitb_13_77 bitb_13_78 R_bl
Cb_13_77 bit_13_77 gnd C_bl
Cbb_13_77 bitb_13_77 gnd C_bl
Rb_13_78 bit_13_78 bit_13_79 R_bl
Rbb_13_78 bitb_13_78 bitb_13_79 R_bl
Cb_13_78 bit_13_78 gnd C_bl
Cbb_13_78 bitb_13_78 gnd C_bl
Rb_13_79 bit_13_79 bit_13_80 R_bl
Rbb_13_79 bitb_13_79 bitb_13_80 R_bl
Cb_13_79 bit_13_79 gnd C_bl
Cbb_13_79 bitb_13_79 gnd C_bl
Rb_13_80 bit_13_80 bit_13_81 R_bl
Rbb_13_80 bitb_13_80 bitb_13_81 R_bl
Cb_13_80 bit_13_80 gnd C_bl
Cbb_13_80 bitb_13_80 gnd C_bl
Rb_13_81 bit_13_81 bit_13_82 R_bl
Rbb_13_81 bitb_13_81 bitb_13_82 R_bl
Cb_13_81 bit_13_81 gnd C_bl
Cbb_13_81 bitb_13_81 gnd C_bl
Rb_13_82 bit_13_82 bit_13_83 R_bl
Rbb_13_82 bitb_13_82 bitb_13_83 R_bl
Cb_13_82 bit_13_82 gnd C_bl
Cbb_13_82 bitb_13_82 gnd C_bl
Rb_13_83 bit_13_83 bit_13_84 R_bl
Rbb_13_83 bitb_13_83 bitb_13_84 R_bl
Cb_13_83 bit_13_83 gnd C_bl
Cbb_13_83 bitb_13_83 gnd C_bl
Rb_13_84 bit_13_84 bit_13_85 R_bl
Rbb_13_84 bitb_13_84 bitb_13_85 R_bl
Cb_13_84 bit_13_84 gnd C_bl
Cbb_13_84 bitb_13_84 gnd C_bl
Rb_13_85 bit_13_85 bit_13_86 R_bl
Rbb_13_85 bitb_13_85 bitb_13_86 R_bl
Cb_13_85 bit_13_85 gnd C_bl
Cbb_13_85 bitb_13_85 gnd C_bl
Rb_13_86 bit_13_86 bit_13_87 R_bl
Rbb_13_86 bitb_13_86 bitb_13_87 R_bl
Cb_13_86 bit_13_86 gnd C_bl
Cbb_13_86 bitb_13_86 gnd C_bl
Rb_13_87 bit_13_87 bit_13_88 R_bl
Rbb_13_87 bitb_13_87 bitb_13_88 R_bl
Cb_13_87 bit_13_87 gnd C_bl
Cbb_13_87 bitb_13_87 gnd C_bl
Rb_13_88 bit_13_88 bit_13_89 R_bl
Rbb_13_88 bitb_13_88 bitb_13_89 R_bl
Cb_13_88 bit_13_88 gnd C_bl
Cbb_13_88 bitb_13_88 gnd C_bl
Rb_13_89 bit_13_89 bit_13_90 R_bl
Rbb_13_89 bitb_13_89 bitb_13_90 R_bl
Cb_13_89 bit_13_89 gnd C_bl
Cbb_13_89 bitb_13_89 gnd C_bl
Rb_13_90 bit_13_90 bit_13_91 R_bl
Rbb_13_90 bitb_13_90 bitb_13_91 R_bl
Cb_13_90 bit_13_90 gnd C_bl
Cbb_13_90 bitb_13_90 gnd C_bl
Rb_13_91 bit_13_91 bit_13_92 R_bl
Rbb_13_91 bitb_13_91 bitb_13_92 R_bl
Cb_13_91 bit_13_91 gnd C_bl
Cbb_13_91 bitb_13_91 gnd C_bl
Rb_13_92 bit_13_92 bit_13_93 R_bl
Rbb_13_92 bitb_13_92 bitb_13_93 R_bl
Cb_13_92 bit_13_92 gnd C_bl
Cbb_13_92 bitb_13_92 gnd C_bl
Rb_13_93 bit_13_93 bit_13_94 R_bl
Rbb_13_93 bitb_13_93 bitb_13_94 R_bl
Cb_13_93 bit_13_93 gnd C_bl
Cbb_13_93 bitb_13_93 gnd C_bl
Rb_13_94 bit_13_94 bit_13_95 R_bl
Rbb_13_94 bitb_13_94 bitb_13_95 R_bl
Cb_13_94 bit_13_94 gnd C_bl
Cbb_13_94 bitb_13_94 gnd C_bl
Rb_13_95 bit_13_95 bit_13_96 R_bl
Rbb_13_95 bitb_13_95 bitb_13_96 R_bl
Cb_13_95 bit_13_95 gnd C_bl
Cbb_13_95 bitb_13_95 gnd C_bl
Rb_13_96 bit_13_96 bit_13_97 R_bl
Rbb_13_96 bitb_13_96 bitb_13_97 R_bl
Cb_13_96 bit_13_96 gnd C_bl
Cbb_13_96 bitb_13_96 gnd C_bl
Rb_13_97 bit_13_97 bit_13_98 R_bl
Rbb_13_97 bitb_13_97 bitb_13_98 R_bl
Cb_13_97 bit_13_97 gnd C_bl
Cbb_13_97 bitb_13_97 gnd C_bl
Rb_13_98 bit_13_98 bit_13_99 R_bl
Rbb_13_98 bitb_13_98 bitb_13_99 R_bl
Cb_13_98 bit_13_98 gnd C_bl
Cbb_13_98 bitb_13_98 gnd C_bl
Rb_13_99 bit_13_99 bit_13_100 R_bl
Rbb_13_99 bitb_13_99 bitb_13_100 R_bl
Cb_13_99 bit_13_99 gnd C_bl
Cbb_13_99 bitb_13_99 gnd C_bl
Rb_14_0 bit_14_0 bit_14_1 R_bl
Rbb_14_0 bitb_14_0 bitb_14_1 R_bl
Cb_14_0 bit_14_0 gnd C_bl
Cbb_14_0 bitb_14_0 gnd C_bl
Rb_14_1 bit_14_1 bit_14_2 R_bl
Rbb_14_1 bitb_14_1 bitb_14_2 R_bl
Cb_14_1 bit_14_1 gnd C_bl
Cbb_14_1 bitb_14_1 gnd C_bl
Rb_14_2 bit_14_2 bit_14_3 R_bl
Rbb_14_2 bitb_14_2 bitb_14_3 R_bl
Cb_14_2 bit_14_2 gnd C_bl
Cbb_14_2 bitb_14_2 gnd C_bl
Rb_14_3 bit_14_3 bit_14_4 R_bl
Rbb_14_3 bitb_14_3 bitb_14_4 R_bl
Cb_14_3 bit_14_3 gnd C_bl
Cbb_14_3 bitb_14_3 gnd C_bl
Rb_14_4 bit_14_4 bit_14_5 R_bl
Rbb_14_4 bitb_14_4 bitb_14_5 R_bl
Cb_14_4 bit_14_4 gnd C_bl
Cbb_14_4 bitb_14_4 gnd C_bl
Rb_14_5 bit_14_5 bit_14_6 R_bl
Rbb_14_5 bitb_14_5 bitb_14_6 R_bl
Cb_14_5 bit_14_5 gnd C_bl
Cbb_14_5 bitb_14_5 gnd C_bl
Rb_14_6 bit_14_6 bit_14_7 R_bl
Rbb_14_6 bitb_14_6 bitb_14_7 R_bl
Cb_14_6 bit_14_6 gnd C_bl
Cbb_14_6 bitb_14_6 gnd C_bl
Rb_14_7 bit_14_7 bit_14_8 R_bl
Rbb_14_7 bitb_14_7 bitb_14_8 R_bl
Cb_14_7 bit_14_7 gnd C_bl
Cbb_14_7 bitb_14_7 gnd C_bl
Rb_14_8 bit_14_8 bit_14_9 R_bl
Rbb_14_8 bitb_14_8 bitb_14_9 R_bl
Cb_14_8 bit_14_8 gnd C_bl
Cbb_14_8 bitb_14_8 gnd C_bl
Rb_14_9 bit_14_9 bit_14_10 R_bl
Rbb_14_9 bitb_14_9 bitb_14_10 R_bl
Cb_14_9 bit_14_9 gnd C_bl
Cbb_14_9 bitb_14_9 gnd C_bl
Rb_14_10 bit_14_10 bit_14_11 R_bl
Rbb_14_10 bitb_14_10 bitb_14_11 R_bl
Cb_14_10 bit_14_10 gnd C_bl
Cbb_14_10 bitb_14_10 gnd C_bl
Rb_14_11 bit_14_11 bit_14_12 R_bl
Rbb_14_11 bitb_14_11 bitb_14_12 R_bl
Cb_14_11 bit_14_11 gnd C_bl
Cbb_14_11 bitb_14_11 gnd C_bl
Rb_14_12 bit_14_12 bit_14_13 R_bl
Rbb_14_12 bitb_14_12 bitb_14_13 R_bl
Cb_14_12 bit_14_12 gnd C_bl
Cbb_14_12 bitb_14_12 gnd C_bl
Rb_14_13 bit_14_13 bit_14_14 R_bl
Rbb_14_13 bitb_14_13 bitb_14_14 R_bl
Cb_14_13 bit_14_13 gnd C_bl
Cbb_14_13 bitb_14_13 gnd C_bl
Rb_14_14 bit_14_14 bit_14_15 R_bl
Rbb_14_14 bitb_14_14 bitb_14_15 R_bl
Cb_14_14 bit_14_14 gnd C_bl
Cbb_14_14 bitb_14_14 gnd C_bl
Rb_14_15 bit_14_15 bit_14_16 R_bl
Rbb_14_15 bitb_14_15 bitb_14_16 R_bl
Cb_14_15 bit_14_15 gnd C_bl
Cbb_14_15 bitb_14_15 gnd C_bl
Rb_14_16 bit_14_16 bit_14_17 R_bl
Rbb_14_16 bitb_14_16 bitb_14_17 R_bl
Cb_14_16 bit_14_16 gnd C_bl
Cbb_14_16 bitb_14_16 gnd C_bl
Rb_14_17 bit_14_17 bit_14_18 R_bl
Rbb_14_17 bitb_14_17 bitb_14_18 R_bl
Cb_14_17 bit_14_17 gnd C_bl
Cbb_14_17 bitb_14_17 gnd C_bl
Rb_14_18 bit_14_18 bit_14_19 R_bl
Rbb_14_18 bitb_14_18 bitb_14_19 R_bl
Cb_14_18 bit_14_18 gnd C_bl
Cbb_14_18 bitb_14_18 gnd C_bl
Rb_14_19 bit_14_19 bit_14_20 R_bl
Rbb_14_19 bitb_14_19 bitb_14_20 R_bl
Cb_14_19 bit_14_19 gnd C_bl
Cbb_14_19 bitb_14_19 gnd C_bl
Rb_14_20 bit_14_20 bit_14_21 R_bl
Rbb_14_20 bitb_14_20 bitb_14_21 R_bl
Cb_14_20 bit_14_20 gnd C_bl
Cbb_14_20 bitb_14_20 gnd C_bl
Rb_14_21 bit_14_21 bit_14_22 R_bl
Rbb_14_21 bitb_14_21 bitb_14_22 R_bl
Cb_14_21 bit_14_21 gnd C_bl
Cbb_14_21 bitb_14_21 gnd C_bl
Rb_14_22 bit_14_22 bit_14_23 R_bl
Rbb_14_22 bitb_14_22 bitb_14_23 R_bl
Cb_14_22 bit_14_22 gnd C_bl
Cbb_14_22 bitb_14_22 gnd C_bl
Rb_14_23 bit_14_23 bit_14_24 R_bl
Rbb_14_23 bitb_14_23 bitb_14_24 R_bl
Cb_14_23 bit_14_23 gnd C_bl
Cbb_14_23 bitb_14_23 gnd C_bl
Rb_14_24 bit_14_24 bit_14_25 R_bl
Rbb_14_24 bitb_14_24 bitb_14_25 R_bl
Cb_14_24 bit_14_24 gnd C_bl
Cbb_14_24 bitb_14_24 gnd C_bl
Rb_14_25 bit_14_25 bit_14_26 R_bl
Rbb_14_25 bitb_14_25 bitb_14_26 R_bl
Cb_14_25 bit_14_25 gnd C_bl
Cbb_14_25 bitb_14_25 gnd C_bl
Rb_14_26 bit_14_26 bit_14_27 R_bl
Rbb_14_26 bitb_14_26 bitb_14_27 R_bl
Cb_14_26 bit_14_26 gnd C_bl
Cbb_14_26 bitb_14_26 gnd C_bl
Rb_14_27 bit_14_27 bit_14_28 R_bl
Rbb_14_27 bitb_14_27 bitb_14_28 R_bl
Cb_14_27 bit_14_27 gnd C_bl
Cbb_14_27 bitb_14_27 gnd C_bl
Rb_14_28 bit_14_28 bit_14_29 R_bl
Rbb_14_28 bitb_14_28 bitb_14_29 R_bl
Cb_14_28 bit_14_28 gnd C_bl
Cbb_14_28 bitb_14_28 gnd C_bl
Rb_14_29 bit_14_29 bit_14_30 R_bl
Rbb_14_29 bitb_14_29 bitb_14_30 R_bl
Cb_14_29 bit_14_29 gnd C_bl
Cbb_14_29 bitb_14_29 gnd C_bl
Rb_14_30 bit_14_30 bit_14_31 R_bl
Rbb_14_30 bitb_14_30 bitb_14_31 R_bl
Cb_14_30 bit_14_30 gnd C_bl
Cbb_14_30 bitb_14_30 gnd C_bl
Rb_14_31 bit_14_31 bit_14_32 R_bl
Rbb_14_31 bitb_14_31 bitb_14_32 R_bl
Cb_14_31 bit_14_31 gnd C_bl
Cbb_14_31 bitb_14_31 gnd C_bl
Rb_14_32 bit_14_32 bit_14_33 R_bl
Rbb_14_32 bitb_14_32 bitb_14_33 R_bl
Cb_14_32 bit_14_32 gnd C_bl
Cbb_14_32 bitb_14_32 gnd C_bl
Rb_14_33 bit_14_33 bit_14_34 R_bl
Rbb_14_33 bitb_14_33 bitb_14_34 R_bl
Cb_14_33 bit_14_33 gnd C_bl
Cbb_14_33 bitb_14_33 gnd C_bl
Rb_14_34 bit_14_34 bit_14_35 R_bl
Rbb_14_34 bitb_14_34 bitb_14_35 R_bl
Cb_14_34 bit_14_34 gnd C_bl
Cbb_14_34 bitb_14_34 gnd C_bl
Rb_14_35 bit_14_35 bit_14_36 R_bl
Rbb_14_35 bitb_14_35 bitb_14_36 R_bl
Cb_14_35 bit_14_35 gnd C_bl
Cbb_14_35 bitb_14_35 gnd C_bl
Rb_14_36 bit_14_36 bit_14_37 R_bl
Rbb_14_36 bitb_14_36 bitb_14_37 R_bl
Cb_14_36 bit_14_36 gnd C_bl
Cbb_14_36 bitb_14_36 gnd C_bl
Rb_14_37 bit_14_37 bit_14_38 R_bl
Rbb_14_37 bitb_14_37 bitb_14_38 R_bl
Cb_14_37 bit_14_37 gnd C_bl
Cbb_14_37 bitb_14_37 gnd C_bl
Rb_14_38 bit_14_38 bit_14_39 R_bl
Rbb_14_38 bitb_14_38 bitb_14_39 R_bl
Cb_14_38 bit_14_38 gnd C_bl
Cbb_14_38 bitb_14_38 gnd C_bl
Rb_14_39 bit_14_39 bit_14_40 R_bl
Rbb_14_39 bitb_14_39 bitb_14_40 R_bl
Cb_14_39 bit_14_39 gnd C_bl
Cbb_14_39 bitb_14_39 gnd C_bl
Rb_14_40 bit_14_40 bit_14_41 R_bl
Rbb_14_40 bitb_14_40 bitb_14_41 R_bl
Cb_14_40 bit_14_40 gnd C_bl
Cbb_14_40 bitb_14_40 gnd C_bl
Rb_14_41 bit_14_41 bit_14_42 R_bl
Rbb_14_41 bitb_14_41 bitb_14_42 R_bl
Cb_14_41 bit_14_41 gnd C_bl
Cbb_14_41 bitb_14_41 gnd C_bl
Rb_14_42 bit_14_42 bit_14_43 R_bl
Rbb_14_42 bitb_14_42 bitb_14_43 R_bl
Cb_14_42 bit_14_42 gnd C_bl
Cbb_14_42 bitb_14_42 gnd C_bl
Rb_14_43 bit_14_43 bit_14_44 R_bl
Rbb_14_43 bitb_14_43 bitb_14_44 R_bl
Cb_14_43 bit_14_43 gnd C_bl
Cbb_14_43 bitb_14_43 gnd C_bl
Rb_14_44 bit_14_44 bit_14_45 R_bl
Rbb_14_44 bitb_14_44 bitb_14_45 R_bl
Cb_14_44 bit_14_44 gnd C_bl
Cbb_14_44 bitb_14_44 gnd C_bl
Rb_14_45 bit_14_45 bit_14_46 R_bl
Rbb_14_45 bitb_14_45 bitb_14_46 R_bl
Cb_14_45 bit_14_45 gnd C_bl
Cbb_14_45 bitb_14_45 gnd C_bl
Rb_14_46 bit_14_46 bit_14_47 R_bl
Rbb_14_46 bitb_14_46 bitb_14_47 R_bl
Cb_14_46 bit_14_46 gnd C_bl
Cbb_14_46 bitb_14_46 gnd C_bl
Rb_14_47 bit_14_47 bit_14_48 R_bl
Rbb_14_47 bitb_14_47 bitb_14_48 R_bl
Cb_14_47 bit_14_47 gnd C_bl
Cbb_14_47 bitb_14_47 gnd C_bl
Rb_14_48 bit_14_48 bit_14_49 R_bl
Rbb_14_48 bitb_14_48 bitb_14_49 R_bl
Cb_14_48 bit_14_48 gnd C_bl
Cbb_14_48 bitb_14_48 gnd C_bl
Rb_14_49 bit_14_49 bit_14_50 R_bl
Rbb_14_49 bitb_14_49 bitb_14_50 R_bl
Cb_14_49 bit_14_49 gnd C_bl
Cbb_14_49 bitb_14_49 gnd C_bl
Rb_14_50 bit_14_50 bit_14_51 R_bl
Rbb_14_50 bitb_14_50 bitb_14_51 R_bl
Cb_14_50 bit_14_50 gnd C_bl
Cbb_14_50 bitb_14_50 gnd C_bl
Rb_14_51 bit_14_51 bit_14_52 R_bl
Rbb_14_51 bitb_14_51 bitb_14_52 R_bl
Cb_14_51 bit_14_51 gnd C_bl
Cbb_14_51 bitb_14_51 gnd C_bl
Rb_14_52 bit_14_52 bit_14_53 R_bl
Rbb_14_52 bitb_14_52 bitb_14_53 R_bl
Cb_14_52 bit_14_52 gnd C_bl
Cbb_14_52 bitb_14_52 gnd C_bl
Rb_14_53 bit_14_53 bit_14_54 R_bl
Rbb_14_53 bitb_14_53 bitb_14_54 R_bl
Cb_14_53 bit_14_53 gnd C_bl
Cbb_14_53 bitb_14_53 gnd C_bl
Rb_14_54 bit_14_54 bit_14_55 R_bl
Rbb_14_54 bitb_14_54 bitb_14_55 R_bl
Cb_14_54 bit_14_54 gnd C_bl
Cbb_14_54 bitb_14_54 gnd C_bl
Rb_14_55 bit_14_55 bit_14_56 R_bl
Rbb_14_55 bitb_14_55 bitb_14_56 R_bl
Cb_14_55 bit_14_55 gnd C_bl
Cbb_14_55 bitb_14_55 gnd C_bl
Rb_14_56 bit_14_56 bit_14_57 R_bl
Rbb_14_56 bitb_14_56 bitb_14_57 R_bl
Cb_14_56 bit_14_56 gnd C_bl
Cbb_14_56 bitb_14_56 gnd C_bl
Rb_14_57 bit_14_57 bit_14_58 R_bl
Rbb_14_57 bitb_14_57 bitb_14_58 R_bl
Cb_14_57 bit_14_57 gnd C_bl
Cbb_14_57 bitb_14_57 gnd C_bl
Rb_14_58 bit_14_58 bit_14_59 R_bl
Rbb_14_58 bitb_14_58 bitb_14_59 R_bl
Cb_14_58 bit_14_58 gnd C_bl
Cbb_14_58 bitb_14_58 gnd C_bl
Rb_14_59 bit_14_59 bit_14_60 R_bl
Rbb_14_59 bitb_14_59 bitb_14_60 R_bl
Cb_14_59 bit_14_59 gnd C_bl
Cbb_14_59 bitb_14_59 gnd C_bl
Rb_14_60 bit_14_60 bit_14_61 R_bl
Rbb_14_60 bitb_14_60 bitb_14_61 R_bl
Cb_14_60 bit_14_60 gnd C_bl
Cbb_14_60 bitb_14_60 gnd C_bl
Rb_14_61 bit_14_61 bit_14_62 R_bl
Rbb_14_61 bitb_14_61 bitb_14_62 R_bl
Cb_14_61 bit_14_61 gnd C_bl
Cbb_14_61 bitb_14_61 gnd C_bl
Rb_14_62 bit_14_62 bit_14_63 R_bl
Rbb_14_62 bitb_14_62 bitb_14_63 R_bl
Cb_14_62 bit_14_62 gnd C_bl
Cbb_14_62 bitb_14_62 gnd C_bl
Rb_14_63 bit_14_63 bit_14_64 R_bl
Rbb_14_63 bitb_14_63 bitb_14_64 R_bl
Cb_14_63 bit_14_63 gnd C_bl
Cbb_14_63 bitb_14_63 gnd C_bl
Rb_14_64 bit_14_64 bit_14_65 R_bl
Rbb_14_64 bitb_14_64 bitb_14_65 R_bl
Cb_14_64 bit_14_64 gnd C_bl
Cbb_14_64 bitb_14_64 gnd C_bl
Rb_14_65 bit_14_65 bit_14_66 R_bl
Rbb_14_65 bitb_14_65 bitb_14_66 R_bl
Cb_14_65 bit_14_65 gnd C_bl
Cbb_14_65 bitb_14_65 gnd C_bl
Rb_14_66 bit_14_66 bit_14_67 R_bl
Rbb_14_66 bitb_14_66 bitb_14_67 R_bl
Cb_14_66 bit_14_66 gnd C_bl
Cbb_14_66 bitb_14_66 gnd C_bl
Rb_14_67 bit_14_67 bit_14_68 R_bl
Rbb_14_67 bitb_14_67 bitb_14_68 R_bl
Cb_14_67 bit_14_67 gnd C_bl
Cbb_14_67 bitb_14_67 gnd C_bl
Rb_14_68 bit_14_68 bit_14_69 R_bl
Rbb_14_68 bitb_14_68 bitb_14_69 R_bl
Cb_14_68 bit_14_68 gnd C_bl
Cbb_14_68 bitb_14_68 gnd C_bl
Rb_14_69 bit_14_69 bit_14_70 R_bl
Rbb_14_69 bitb_14_69 bitb_14_70 R_bl
Cb_14_69 bit_14_69 gnd C_bl
Cbb_14_69 bitb_14_69 gnd C_bl
Rb_14_70 bit_14_70 bit_14_71 R_bl
Rbb_14_70 bitb_14_70 bitb_14_71 R_bl
Cb_14_70 bit_14_70 gnd C_bl
Cbb_14_70 bitb_14_70 gnd C_bl
Rb_14_71 bit_14_71 bit_14_72 R_bl
Rbb_14_71 bitb_14_71 bitb_14_72 R_bl
Cb_14_71 bit_14_71 gnd C_bl
Cbb_14_71 bitb_14_71 gnd C_bl
Rb_14_72 bit_14_72 bit_14_73 R_bl
Rbb_14_72 bitb_14_72 bitb_14_73 R_bl
Cb_14_72 bit_14_72 gnd C_bl
Cbb_14_72 bitb_14_72 gnd C_bl
Rb_14_73 bit_14_73 bit_14_74 R_bl
Rbb_14_73 bitb_14_73 bitb_14_74 R_bl
Cb_14_73 bit_14_73 gnd C_bl
Cbb_14_73 bitb_14_73 gnd C_bl
Rb_14_74 bit_14_74 bit_14_75 R_bl
Rbb_14_74 bitb_14_74 bitb_14_75 R_bl
Cb_14_74 bit_14_74 gnd C_bl
Cbb_14_74 bitb_14_74 gnd C_bl
Rb_14_75 bit_14_75 bit_14_76 R_bl
Rbb_14_75 bitb_14_75 bitb_14_76 R_bl
Cb_14_75 bit_14_75 gnd C_bl
Cbb_14_75 bitb_14_75 gnd C_bl
Rb_14_76 bit_14_76 bit_14_77 R_bl
Rbb_14_76 bitb_14_76 bitb_14_77 R_bl
Cb_14_76 bit_14_76 gnd C_bl
Cbb_14_76 bitb_14_76 gnd C_bl
Rb_14_77 bit_14_77 bit_14_78 R_bl
Rbb_14_77 bitb_14_77 bitb_14_78 R_bl
Cb_14_77 bit_14_77 gnd C_bl
Cbb_14_77 bitb_14_77 gnd C_bl
Rb_14_78 bit_14_78 bit_14_79 R_bl
Rbb_14_78 bitb_14_78 bitb_14_79 R_bl
Cb_14_78 bit_14_78 gnd C_bl
Cbb_14_78 bitb_14_78 gnd C_bl
Rb_14_79 bit_14_79 bit_14_80 R_bl
Rbb_14_79 bitb_14_79 bitb_14_80 R_bl
Cb_14_79 bit_14_79 gnd C_bl
Cbb_14_79 bitb_14_79 gnd C_bl
Rb_14_80 bit_14_80 bit_14_81 R_bl
Rbb_14_80 bitb_14_80 bitb_14_81 R_bl
Cb_14_80 bit_14_80 gnd C_bl
Cbb_14_80 bitb_14_80 gnd C_bl
Rb_14_81 bit_14_81 bit_14_82 R_bl
Rbb_14_81 bitb_14_81 bitb_14_82 R_bl
Cb_14_81 bit_14_81 gnd C_bl
Cbb_14_81 bitb_14_81 gnd C_bl
Rb_14_82 bit_14_82 bit_14_83 R_bl
Rbb_14_82 bitb_14_82 bitb_14_83 R_bl
Cb_14_82 bit_14_82 gnd C_bl
Cbb_14_82 bitb_14_82 gnd C_bl
Rb_14_83 bit_14_83 bit_14_84 R_bl
Rbb_14_83 bitb_14_83 bitb_14_84 R_bl
Cb_14_83 bit_14_83 gnd C_bl
Cbb_14_83 bitb_14_83 gnd C_bl
Rb_14_84 bit_14_84 bit_14_85 R_bl
Rbb_14_84 bitb_14_84 bitb_14_85 R_bl
Cb_14_84 bit_14_84 gnd C_bl
Cbb_14_84 bitb_14_84 gnd C_bl
Rb_14_85 bit_14_85 bit_14_86 R_bl
Rbb_14_85 bitb_14_85 bitb_14_86 R_bl
Cb_14_85 bit_14_85 gnd C_bl
Cbb_14_85 bitb_14_85 gnd C_bl
Rb_14_86 bit_14_86 bit_14_87 R_bl
Rbb_14_86 bitb_14_86 bitb_14_87 R_bl
Cb_14_86 bit_14_86 gnd C_bl
Cbb_14_86 bitb_14_86 gnd C_bl
Rb_14_87 bit_14_87 bit_14_88 R_bl
Rbb_14_87 bitb_14_87 bitb_14_88 R_bl
Cb_14_87 bit_14_87 gnd C_bl
Cbb_14_87 bitb_14_87 gnd C_bl
Rb_14_88 bit_14_88 bit_14_89 R_bl
Rbb_14_88 bitb_14_88 bitb_14_89 R_bl
Cb_14_88 bit_14_88 gnd C_bl
Cbb_14_88 bitb_14_88 gnd C_bl
Rb_14_89 bit_14_89 bit_14_90 R_bl
Rbb_14_89 bitb_14_89 bitb_14_90 R_bl
Cb_14_89 bit_14_89 gnd C_bl
Cbb_14_89 bitb_14_89 gnd C_bl
Rb_14_90 bit_14_90 bit_14_91 R_bl
Rbb_14_90 bitb_14_90 bitb_14_91 R_bl
Cb_14_90 bit_14_90 gnd C_bl
Cbb_14_90 bitb_14_90 gnd C_bl
Rb_14_91 bit_14_91 bit_14_92 R_bl
Rbb_14_91 bitb_14_91 bitb_14_92 R_bl
Cb_14_91 bit_14_91 gnd C_bl
Cbb_14_91 bitb_14_91 gnd C_bl
Rb_14_92 bit_14_92 bit_14_93 R_bl
Rbb_14_92 bitb_14_92 bitb_14_93 R_bl
Cb_14_92 bit_14_92 gnd C_bl
Cbb_14_92 bitb_14_92 gnd C_bl
Rb_14_93 bit_14_93 bit_14_94 R_bl
Rbb_14_93 bitb_14_93 bitb_14_94 R_bl
Cb_14_93 bit_14_93 gnd C_bl
Cbb_14_93 bitb_14_93 gnd C_bl
Rb_14_94 bit_14_94 bit_14_95 R_bl
Rbb_14_94 bitb_14_94 bitb_14_95 R_bl
Cb_14_94 bit_14_94 gnd C_bl
Cbb_14_94 bitb_14_94 gnd C_bl
Rb_14_95 bit_14_95 bit_14_96 R_bl
Rbb_14_95 bitb_14_95 bitb_14_96 R_bl
Cb_14_95 bit_14_95 gnd C_bl
Cbb_14_95 bitb_14_95 gnd C_bl
Rb_14_96 bit_14_96 bit_14_97 R_bl
Rbb_14_96 bitb_14_96 bitb_14_97 R_bl
Cb_14_96 bit_14_96 gnd C_bl
Cbb_14_96 bitb_14_96 gnd C_bl
Rb_14_97 bit_14_97 bit_14_98 R_bl
Rbb_14_97 bitb_14_97 bitb_14_98 R_bl
Cb_14_97 bit_14_97 gnd C_bl
Cbb_14_97 bitb_14_97 gnd C_bl
Rb_14_98 bit_14_98 bit_14_99 R_bl
Rbb_14_98 bitb_14_98 bitb_14_99 R_bl
Cb_14_98 bit_14_98 gnd C_bl
Cbb_14_98 bitb_14_98 gnd C_bl
Rb_14_99 bit_14_99 bit_14_100 R_bl
Rbb_14_99 bitb_14_99 bitb_14_100 R_bl
Cb_14_99 bit_14_99 gnd C_bl
Cbb_14_99 bitb_14_99 gnd C_bl
Rb_15_0 bit_15_0 bit_15_1 R_bl
Rbb_15_0 bitb_15_0 bitb_15_1 R_bl
Cb_15_0 bit_15_0 gnd C_bl
Cbb_15_0 bitb_15_0 gnd C_bl
Rb_15_1 bit_15_1 bit_15_2 R_bl
Rbb_15_1 bitb_15_1 bitb_15_2 R_bl
Cb_15_1 bit_15_1 gnd C_bl
Cbb_15_1 bitb_15_1 gnd C_bl
Rb_15_2 bit_15_2 bit_15_3 R_bl
Rbb_15_2 bitb_15_2 bitb_15_3 R_bl
Cb_15_2 bit_15_2 gnd C_bl
Cbb_15_2 bitb_15_2 gnd C_bl
Rb_15_3 bit_15_3 bit_15_4 R_bl
Rbb_15_3 bitb_15_3 bitb_15_4 R_bl
Cb_15_3 bit_15_3 gnd C_bl
Cbb_15_3 bitb_15_3 gnd C_bl
Rb_15_4 bit_15_4 bit_15_5 R_bl
Rbb_15_4 bitb_15_4 bitb_15_5 R_bl
Cb_15_4 bit_15_4 gnd C_bl
Cbb_15_4 bitb_15_4 gnd C_bl
Rb_15_5 bit_15_5 bit_15_6 R_bl
Rbb_15_5 bitb_15_5 bitb_15_6 R_bl
Cb_15_5 bit_15_5 gnd C_bl
Cbb_15_5 bitb_15_5 gnd C_bl
Rb_15_6 bit_15_6 bit_15_7 R_bl
Rbb_15_6 bitb_15_6 bitb_15_7 R_bl
Cb_15_6 bit_15_6 gnd C_bl
Cbb_15_6 bitb_15_6 gnd C_bl
Rb_15_7 bit_15_7 bit_15_8 R_bl
Rbb_15_7 bitb_15_7 bitb_15_8 R_bl
Cb_15_7 bit_15_7 gnd C_bl
Cbb_15_7 bitb_15_7 gnd C_bl
Rb_15_8 bit_15_8 bit_15_9 R_bl
Rbb_15_8 bitb_15_8 bitb_15_9 R_bl
Cb_15_8 bit_15_8 gnd C_bl
Cbb_15_8 bitb_15_8 gnd C_bl
Rb_15_9 bit_15_9 bit_15_10 R_bl
Rbb_15_9 bitb_15_9 bitb_15_10 R_bl
Cb_15_9 bit_15_9 gnd C_bl
Cbb_15_9 bitb_15_9 gnd C_bl
Rb_15_10 bit_15_10 bit_15_11 R_bl
Rbb_15_10 bitb_15_10 bitb_15_11 R_bl
Cb_15_10 bit_15_10 gnd C_bl
Cbb_15_10 bitb_15_10 gnd C_bl
Rb_15_11 bit_15_11 bit_15_12 R_bl
Rbb_15_11 bitb_15_11 bitb_15_12 R_bl
Cb_15_11 bit_15_11 gnd C_bl
Cbb_15_11 bitb_15_11 gnd C_bl
Rb_15_12 bit_15_12 bit_15_13 R_bl
Rbb_15_12 bitb_15_12 bitb_15_13 R_bl
Cb_15_12 bit_15_12 gnd C_bl
Cbb_15_12 bitb_15_12 gnd C_bl
Rb_15_13 bit_15_13 bit_15_14 R_bl
Rbb_15_13 bitb_15_13 bitb_15_14 R_bl
Cb_15_13 bit_15_13 gnd C_bl
Cbb_15_13 bitb_15_13 gnd C_bl
Rb_15_14 bit_15_14 bit_15_15 R_bl
Rbb_15_14 bitb_15_14 bitb_15_15 R_bl
Cb_15_14 bit_15_14 gnd C_bl
Cbb_15_14 bitb_15_14 gnd C_bl
Rb_15_15 bit_15_15 bit_15_16 R_bl
Rbb_15_15 bitb_15_15 bitb_15_16 R_bl
Cb_15_15 bit_15_15 gnd C_bl
Cbb_15_15 bitb_15_15 gnd C_bl
Rb_15_16 bit_15_16 bit_15_17 R_bl
Rbb_15_16 bitb_15_16 bitb_15_17 R_bl
Cb_15_16 bit_15_16 gnd C_bl
Cbb_15_16 bitb_15_16 gnd C_bl
Rb_15_17 bit_15_17 bit_15_18 R_bl
Rbb_15_17 bitb_15_17 bitb_15_18 R_bl
Cb_15_17 bit_15_17 gnd C_bl
Cbb_15_17 bitb_15_17 gnd C_bl
Rb_15_18 bit_15_18 bit_15_19 R_bl
Rbb_15_18 bitb_15_18 bitb_15_19 R_bl
Cb_15_18 bit_15_18 gnd C_bl
Cbb_15_18 bitb_15_18 gnd C_bl
Rb_15_19 bit_15_19 bit_15_20 R_bl
Rbb_15_19 bitb_15_19 bitb_15_20 R_bl
Cb_15_19 bit_15_19 gnd C_bl
Cbb_15_19 bitb_15_19 gnd C_bl
Rb_15_20 bit_15_20 bit_15_21 R_bl
Rbb_15_20 bitb_15_20 bitb_15_21 R_bl
Cb_15_20 bit_15_20 gnd C_bl
Cbb_15_20 bitb_15_20 gnd C_bl
Rb_15_21 bit_15_21 bit_15_22 R_bl
Rbb_15_21 bitb_15_21 bitb_15_22 R_bl
Cb_15_21 bit_15_21 gnd C_bl
Cbb_15_21 bitb_15_21 gnd C_bl
Rb_15_22 bit_15_22 bit_15_23 R_bl
Rbb_15_22 bitb_15_22 bitb_15_23 R_bl
Cb_15_22 bit_15_22 gnd C_bl
Cbb_15_22 bitb_15_22 gnd C_bl
Rb_15_23 bit_15_23 bit_15_24 R_bl
Rbb_15_23 bitb_15_23 bitb_15_24 R_bl
Cb_15_23 bit_15_23 gnd C_bl
Cbb_15_23 bitb_15_23 gnd C_bl
Rb_15_24 bit_15_24 bit_15_25 R_bl
Rbb_15_24 bitb_15_24 bitb_15_25 R_bl
Cb_15_24 bit_15_24 gnd C_bl
Cbb_15_24 bitb_15_24 gnd C_bl
Rb_15_25 bit_15_25 bit_15_26 R_bl
Rbb_15_25 bitb_15_25 bitb_15_26 R_bl
Cb_15_25 bit_15_25 gnd C_bl
Cbb_15_25 bitb_15_25 gnd C_bl
Rb_15_26 bit_15_26 bit_15_27 R_bl
Rbb_15_26 bitb_15_26 bitb_15_27 R_bl
Cb_15_26 bit_15_26 gnd C_bl
Cbb_15_26 bitb_15_26 gnd C_bl
Rb_15_27 bit_15_27 bit_15_28 R_bl
Rbb_15_27 bitb_15_27 bitb_15_28 R_bl
Cb_15_27 bit_15_27 gnd C_bl
Cbb_15_27 bitb_15_27 gnd C_bl
Rb_15_28 bit_15_28 bit_15_29 R_bl
Rbb_15_28 bitb_15_28 bitb_15_29 R_bl
Cb_15_28 bit_15_28 gnd C_bl
Cbb_15_28 bitb_15_28 gnd C_bl
Rb_15_29 bit_15_29 bit_15_30 R_bl
Rbb_15_29 bitb_15_29 bitb_15_30 R_bl
Cb_15_29 bit_15_29 gnd C_bl
Cbb_15_29 bitb_15_29 gnd C_bl
Rb_15_30 bit_15_30 bit_15_31 R_bl
Rbb_15_30 bitb_15_30 bitb_15_31 R_bl
Cb_15_30 bit_15_30 gnd C_bl
Cbb_15_30 bitb_15_30 gnd C_bl
Rb_15_31 bit_15_31 bit_15_32 R_bl
Rbb_15_31 bitb_15_31 bitb_15_32 R_bl
Cb_15_31 bit_15_31 gnd C_bl
Cbb_15_31 bitb_15_31 gnd C_bl
Rb_15_32 bit_15_32 bit_15_33 R_bl
Rbb_15_32 bitb_15_32 bitb_15_33 R_bl
Cb_15_32 bit_15_32 gnd C_bl
Cbb_15_32 bitb_15_32 gnd C_bl
Rb_15_33 bit_15_33 bit_15_34 R_bl
Rbb_15_33 bitb_15_33 bitb_15_34 R_bl
Cb_15_33 bit_15_33 gnd C_bl
Cbb_15_33 bitb_15_33 gnd C_bl
Rb_15_34 bit_15_34 bit_15_35 R_bl
Rbb_15_34 bitb_15_34 bitb_15_35 R_bl
Cb_15_34 bit_15_34 gnd C_bl
Cbb_15_34 bitb_15_34 gnd C_bl
Rb_15_35 bit_15_35 bit_15_36 R_bl
Rbb_15_35 bitb_15_35 bitb_15_36 R_bl
Cb_15_35 bit_15_35 gnd C_bl
Cbb_15_35 bitb_15_35 gnd C_bl
Rb_15_36 bit_15_36 bit_15_37 R_bl
Rbb_15_36 bitb_15_36 bitb_15_37 R_bl
Cb_15_36 bit_15_36 gnd C_bl
Cbb_15_36 bitb_15_36 gnd C_bl
Rb_15_37 bit_15_37 bit_15_38 R_bl
Rbb_15_37 bitb_15_37 bitb_15_38 R_bl
Cb_15_37 bit_15_37 gnd C_bl
Cbb_15_37 bitb_15_37 gnd C_bl
Rb_15_38 bit_15_38 bit_15_39 R_bl
Rbb_15_38 bitb_15_38 bitb_15_39 R_bl
Cb_15_38 bit_15_38 gnd C_bl
Cbb_15_38 bitb_15_38 gnd C_bl
Rb_15_39 bit_15_39 bit_15_40 R_bl
Rbb_15_39 bitb_15_39 bitb_15_40 R_bl
Cb_15_39 bit_15_39 gnd C_bl
Cbb_15_39 bitb_15_39 gnd C_bl
Rb_15_40 bit_15_40 bit_15_41 R_bl
Rbb_15_40 bitb_15_40 bitb_15_41 R_bl
Cb_15_40 bit_15_40 gnd C_bl
Cbb_15_40 bitb_15_40 gnd C_bl
Rb_15_41 bit_15_41 bit_15_42 R_bl
Rbb_15_41 bitb_15_41 bitb_15_42 R_bl
Cb_15_41 bit_15_41 gnd C_bl
Cbb_15_41 bitb_15_41 gnd C_bl
Rb_15_42 bit_15_42 bit_15_43 R_bl
Rbb_15_42 bitb_15_42 bitb_15_43 R_bl
Cb_15_42 bit_15_42 gnd C_bl
Cbb_15_42 bitb_15_42 gnd C_bl
Rb_15_43 bit_15_43 bit_15_44 R_bl
Rbb_15_43 bitb_15_43 bitb_15_44 R_bl
Cb_15_43 bit_15_43 gnd C_bl
Cbb_15_43 bitb_15_43 gnd C_bl
Rb_15_44 bit_15_44 bit_15_45 R_bl
Rbb_15_44 bitb_15_44 bitb_15_45 R_bl
Cb_15_44 bit_15_44 gnd C_bl
Cbb_15_44 bitb_15_44 gnd C_bl
Rb_15_45 bit_15_45 bit_15_46 R_bl
Rbb_15_45 bitb_15_45 bitb_15_46 R_bl
Cb_15_45 bit_15_45 gnd C_bl
Cbb_15_45 bitb_15_45 gnd C_bl
Rb_15_46 bit_15_46 bit_15_47 R_bl
Rbb_15_46 bitb_15_46 bitb_15_47 R_bl
Cb_15_46 bit_15_46 gnd C_bl
Cbb_15_46 bitb_15_46 gnd C_bl
Rb_15_47 bit_15_47 bit_15_48 R_bl
Rbb_15_47 bitb_15_47 bitb_15_48 R_bl
Cb_15_47 bit_15_47 gnd C_bl
Cbb_15_47 bitb_15_47 gnd C_bl
Rb_15_48 bit_15_48 bit_15_49 R_bl
Rbb_15_48 bitb_15_48 bitb_15_49 R_bl
Cb_15_48 bit_15_48 gnd C_bl
Cbb_15_48 bitb_15_48 gnd C_bl
Rb_15_49 bit_15_49 bit_15_50 R_bl
Rbb_15_49 bitb_15_49 bitb_15_50 R_bl
Cb_15_49 bit_15_49 gnd C_bl
Cbb_15_49 bitb_15_49 gnd C_bl
Rb_15_50 bit_15_50 bit_15_51 R_bl
Rbb_15_50 bitb_15_50 bitb_15_51 R_bl
Cb_15_50 bit_15_50 gnd C_bl
Cbb_15_50 bitb_15_50 gnd C_bl
Rb_15_51 bit_15_51 bit_15_52 R_bl
Rbb_15_51 bitb_15_51 bitb_15_52 R_bl
Cb_15_51 bit_15_51 gnd C_bl
Cbb_15_51 bitb_15_51 gnd C_bl
Rb_15_52 bit_15_52 bit_15_53 R_bl
Rbb_15_52 bitb_15_52 bitb_15_53 R_bl
Cb_15_52 bit_15_52 gnd C_bl
Cbb_15_52 bitb_15_52 gnd C_bl
Rb_15_53 bit_15_53 bit_15_54 R_bl
Rbb_15_53 bitb_15_53 bitb_15_54 R_bl
Cb_15_53 bit_15_53 gnd C_bl
Cbb_15_53 bitb_15_53 gnd C_bl
Rb_15_54 bit_15_54 bit_15_55 R_bl
Rbb_15_54 bitb_15_54 bitb_15_55 R_bl
Cb_15_54 bit_15_54 gnd C_bl
Cbb_15_54 bitb_15_54 gnd C_bl
Rb_15_55 bit_15_55 bit_15_56 R_bl
Rbb_15_55 bitb_15_55 bitb_15_56 R_bl
Cb_15_55 bit_15_55 gnd C_bl
Cbb_15_55 bitb_15_55 gnd C_bl
Rb_15_56 bit_15_56 bit_15_57 R_bl
Rbb_15_56 bitb_15_56 bitb_15_57 R_bl
Cb_15_56 bit_15_56 gnd C_bl
Cbb_15_56 bitb_15_56 gnd C_bl
Rb_15_57 bit_15_57 bit_15_58 R_bl
Rbb_15_57 bitb_15_57 bitb_15_58 R_bl
Cb_15_57 bit_15_57 gnd C_bl
Cbb_15_57 bitb_15_57 gnd C_bl
Rb_15_58 bit_15_58 bit_15_59 R_bl
Rbb_15_58 bitb_15_58 bitb_15_59 R_bl
Cb_15_58 bit_15_58 gnd C_bl
Cbb_15_58 bitb_15_58 gnd C_bl
Rb_15_59 bit_15_59 bit_15_60 R_bl
Rbb_15_59 bitb_15_59 bitb_15_60 R_bl
Cb_15_59 bit_15_59 gnd C_bl
Cbb_15_59 bitb_15_59 gnd C_bl
Rb_15_60 bit_15_60 bit_15_61 R_bl
Rbb_15_60 bitb_15_60 bitb_15_61 R_bl
Cb_15_60 bit_15_60 gnd C_bl
Cbb_15_60 bitb_15_60 gnd C_bl
Rb_15_61 bit_15_61 bit_15_62 R_bl
Rbb_15_61 bitb_15_61 bitb_15_62 R_bl
Cb_15_61 bit_15_61 gnd C_bl
Cbb_15_61 bitb_15_61 gnd C_bl
Rb_15_62 bit_15_62 bit_15_63 R_bl
Rbb_15_62 bitb_15_62 bitb_15_63 R_bl
Cb_15_62 bit_15_62 gnd C_bl
Cbb_15_62 bitb_15_62 gnd C_bl
Rb_15_63 bit_15_63 bit_15_64 R_bl
Rbb_15_63 bitb_15_63 bitb_15_64 R_bl
Cb_15_63 bit_15_63 gnd C_bl
Cbb_15_63 bitb_15_63 gnd C_bl
Rb_15_64 bit_15_64 bit_15_65 R_bl
Rbb_15_64 bitb_15_64 bitb_15_65 R_bl
Cb_15_64 bit_15_64 gnd C_bl
Cbb_15_64 bitb_15_64 gnd C_bl
Rb_15_65 bit_15_65 bit_15_66 R_bl
Rbb_15_65 bitb_15_65 bitb_15_66 R_bl
Cb_15_65 bit_15_65 gnd C_bl
Cbb_15_65 bitb_15_65 gnd C_bl
Rb_15_66 bit_15_66 bit_15_67 R_bl
Rbb_15_66 bitb_15_66 bitb_15_67 R_bl
Cb_15_66 bit_15_66 gnd C_bl
Cbb_15_66 bitb_15_66 gnd C_bl
Rb_15_67 bit_15_67 bit_15_68 R_bl
Rbb_15_67 bitb_15_67 bitb_15_68 R_bl
Cb_15_67 bit_15_67 gnd C_bl
Cbb_15_67 bitb_15_67 gnd C_bl
Rb_15_68 bit_15_68 bit_15_69 R_bl
Rbb_15_68 bitb_15_68 bitb_15_69 R_bl
Cb_15_68 bit_15_68 gnd C_bl
Cbb_15_68 bitb_15_68 gnd C_bl
Rb_15_69 bit_15_69 bit_15_70 R_bl
Rbb_15_69 bitb_15_69 bitb_15_70 R_bl
Cb_15_69 bit_15_69 gnd C_bl
Cbb_15_69 bitb_15_69 gnd C_bl
Rb_15_70 bit_15_70 bit_15_71 R_bl
Rbb_15_70 bitb_15_70 bitb_15_71 R_bl
Cb_15_70 bit_15_70 gnd C_bl
Cbb_15_70 bitb_15_70 gnd C_bl
Rb_15_71 bit_15_71 bit_15_72 R_bl
Rbb_15_71 bitb_15_71 bitb_15_72 R_bl
Cb_15_71 bit_15_71 gnd C_bl
Cbb_15_71 bitb_15_71 gnd C_bl
Rb_15_72 bit_15_72 bit_15_73 R_bl
Rbb_15_72 bitb_15_72 bitb_15_73 R_bl
Cb_15_72 bit_15_72 gnd C_bl
Cbb_15_72 bitb_15_72 gnd C_bl
Rb_15_73 bit_15_73 bit_15_74 R_bl
Rbb_15_73 bitb_15_73 bitb_15_74 R_bl
Cb_15_73 bit_15_73 gnd C_bl
Cbb_15_73 bitb_15_73 gnd C_bl
Rb_15_74 bit_15_74 bit_15_75 R_bl
Rbb_15_74 bitb_15_74 bitb_15_75 R_bl
Cb_15_74 bit_15_74 gnd C_bl
Cbb_15_74 bitb_15_74 gnd C_bl
Rb_15_75 bit_15_75 bit_15_76 R_bl
Rbb_15_75 bitb_15_75 bitb_15_76 R_bl
Cb_15_75 bit_15_75 gnd C_bl
Cbb_15_75 bitb_15_75 gnd C_bl
Rb_15_76 bit_15_76 bit_15_77 R_bl
Rbb_15_76 bitb_15_76 bitb_15_77 R_bl
Cb_15_76 bit_15_76 gnd C_bl
Cbb_15_76 bitb_15_76 gnd C_bl
Rb_15_77 bit_15_77 bit_15_78 R_bl
Rbb_15_77 bitb_15_77 bitb_15_78 R_bl
Cb_15_77 bit_15_77 gnd C_bl
Cbb_15_77 bitb_15_77 gnd C_bl
Rb_15_78 bit_15_78 bit_15_79 R_bl
Rbb_15_78 bitb_15_78 bitb_15_79 R_bl
Cb_15_78 bit_15_78 gnd C_bl
Cbb_15_78 bitb_15_78 gnd C_bl
Rb_15_79 bit_15_79 bit_15_80 R_bl
Rbb_15_79 bitb_15_79 bitb_15_80 R_bl
Cb_15_79 bit_15_79 gnd C_bl
Cbb_15_79 bitb_15_79 gnd C_bl
Rb_15_80 bit_15_80 bit_15_81 R_bl
Rbb_15_80 bitb_15_80 bitb_15_81 R_bl
Cb_15_80 bit_15_80 gnd C_bl
Cbb_15_80 bitb_15_80 gnd C_bl
Rb_15_81 bit_15_81 bit_15_82 R_bl
Rbb_15_81 bitb_15_81 bitb_15_82 R_bl
Cb_15_81 bit_15_81 gnd C_bl
Cbb_15_81 bitb_15_81 gnd C_bl
Rb_15_82 bit_15_82 bit_15_83 R_bl
Rbb_15_82 bitb_15_82 bitb_15_83 R_bl
Cb_15_82 bit_15_82 gnd C_bl
Cbb_15_82 bitb_15_82 gnd C_bl
Rb_15_83 bit_15_83 bit_15_84 R_bl
Rbb_15_83 bitb_15_83 bitb_15_84 R_bl
Cb_15_83 bit_15_83 gnd C_bl
Cbb_15_83 bitb_15_83 gnd C_bl
Rb_15_84 bit_15_84 bit_15_85 R_bl
Rbb_15_84 bitb_15_84 bitb_15_85 R_bl
Cb_15_84 bit_15_84 gnd C_bl
Cbb_15_84 bitb_15_84 gnd C_bl
Rb_15_85 bit_15_85 bit_15_86 R_bl
Rbb_15_85 bitb_15_85 bitb_15_86 R_bl
Cb_15_85 bit_15_85 gnd C_bl
Cbb_15_85 bitb_15_85 gnd C_bl
Rb_15_86 bit_15_86 bit_15_87 R_bl
Rbb_15_86 bitb_15_86 bitb_15_87 R_bl
Cb_15_86 bit_15_86 gnd C_bl
Cbb_15_86 bitb_15_86 gnd C_bl
Rb_15_87 bit_15_87 bit_15_88 R_bl
Rbb_15_87 bitb_15_87 bitb_15_88 R_bl
Cb_15_87 bit_15_87 gnd C_bl
Cbb_15_87 bitb_15_87 gnd C_bl
Rb_15_88 bit_15_88 bit_15_89 R_bl
Rbb_15_88 bitb_15_88 bitb_15_89 R_bl
Cb_15_88 bit_15_88 gnd C_bl
Cbb_15_88 bitb_15_88 gnd C_bl
Rb_15_89 bit_15_89 bit_15_90 R_bl
Rbb_15_89 bitb_15_89 bitb_15_90 R_bl
Cb_15_89 bit_15_89 gnd C_bl
Cbb_15_89 bitb_15_89 gnd C_bl
Rb_15_90 bit_15_90 bit_15_91 R_bl
Rbb_15_90 bitb_15_90 bitb_15_91 R_bl
Cb_15_90 bit_15_90 gnd C_bl
Cbb_15_90 bitb_15_90 gnd C_bl
Rb_15_91 bit_15_91 bit_15_92 R_bl
Rbb_15_91 bitb_15_91 bitb_15_92 R_bl
Cb_15_91 bit_15_91 gnd C_bl
Cbb_15_91 bitb_15_91 gnd C_bl
Rb_15_92 bit_15_92 bit_15_93 R_bl
Rbb_15_92 bitb_15_92 bitb_15_93 R_bl
Cb_15_92 bit_15_92 gnd C_bl
Cbb_15_92 bitb_15_92 gnd C_bl
Rb_15_93 bit_15_93 bit_15_94 R_bl
Rbb_15_93 bitb_15_93 bitb_15_94 R_bl
Cb_15_93 bit_15_93 gnd C_bl
Cbb_15_93 bitb_15_93 gnd C_bl
Rb_15_94 bit_15_94 bit_15_95 R_bl
Rbb_15_94 bitb_15_94 bitb_15_95 R_bl
Cb_15_94 bit_15_94 gnd C_bl
Cbb_15_94 bitb_15_94 gnd C_bl
Rb_15_95 bit_15_95 bit_15_96 R_bl
Rbb_15_95 bitb_15_95 bitb_15_96 R_bl
Cb_15_95 bit_15_95 gnd C_bl
Cbb_15_95 bitb_15_95 gnd C_bl
Rb_15_96 bit_15_96 bit_15_97 R_bl
Rbb_15_96 bitb_15_96 bitb_15_97 R_bl
Cb_15_96 bit_15_96 gnd C_bl
Cbb_15_96 bitb_15_96 gnd C_bl
Rb_15_97 bit_15_97 bit_15_98 R_bl
Rbb_15_97 bitb_15_97 bitb_15_98 R_bl
Cb_15_97 bit_15_97 gnd C_bl
Cbb_15_97 bitb_15_97 gnd C_bl
Rb_15_98 bit_15_98 bit_15_99 R_bl
Rbb_15_98 bitb_15_98 bitb_15_99 R_bl
Cb_15_98 bit_15_98 gnd C_bl
Cbb_15_98 bitb_15_98 gnd C_bl
Rb_15_99 bit_15_99 bit_15_100 R_bl
Rbb_15_99 bitb_15_99 bitb_15_100 R_bl
Cb_15_99 bit_15_99 gnd C_bl
Cbb_15_99 bitb_15_99 gnd C_bl
Rb_16_0 bit_16_0 bit_16_1 R_bl
Rbb_16_0 bitb_16_0 bitb_16_1 R_bl
Cb_16_0 bit_16_0 gnd C_bl
Cbb_16_0 bitb_16_0 gnd C_bl
Rb_16_1 bit_16_1 bit_16_2 R_bl
Rbb_16_1 bitb_16_1 bitb_16_2 R_bl
Cb_16_1 bit_16_1 gnd C_bl
Cbb_16_1 bitb_16_1 gnd C_bl
Rb_16_2 bit_16_2 bit_16_3 R_bl
Rbb_16_2 bitb_16_2 bitb_16_3 R_bl
Cb_16_2 bit_16_2 gnd C_bl
Cbb_16_2 bitb_16_2 gnd C_bl
Rb_16_3 bit_16_3 bit_16_4 R_bl
Rbb_16_3 bitb_16_3 bitb_16_4 R_bl
Cb_16_3 bit_16_3 gnd C_bl
Cbb_16_3 bitb_16_3 gnd C_bl
Rb_16_4 bit_16_4 bit_16_5 R_bl
Rbb_16_4 bitb_16_4 bitb_16_5 R_bl
Cb_16_4 bit_16_4 gnd C_bl
Cbb_16_4 bitb_16_4 gnd C_bl
Rb_16_5 bit_16_5 bit_16_6 R_bl
Rbb_16_5 bitb_16_5 bitb_16_6 R_bl
Cb_16_5 bit_16_5 gnd C_bl
Cbb_16_5 bitb_16_5 gnd C_bl
Rb_16_6 bit_16_6 bit_16_7 R_bl
Rbb_16_6 bitb_16_6 bitb_16_7 R_bl
Cb_16_6 bit_16_6 gnd C_bl
Cbb_16_6 bitb_16_6 gnd C_bl
Rb_16_7 bit_16_7 bit_16_8 R_bl
Rbb_16_7 bitb_16_7 bitb_16_8 R_bl
Cb_16_7 bit_16_7 gnd C_bl
Cbb_16_7 bitb_16_7 gnd C_bl
Rb_16_8 bit_16_8 bit_16_9 R_bl
Rbb_16_8 bitb_16_8 bitb_16_9 R_bl
Cb_16_8 bit_16_8 gnd C_bl
Cbb_16_8 bitb_16_8 gnd C_bl
Rb_16_9 bit_16_9 bit_16_10 R_bl
Rbb_16_9 bitb_16_9 bitb_16_10 R_bl
Cb_16_9 bit_16_9 gnd C_bl
Cbb_16_9 bitb_16_9 gnd C_bl
Rb_16_10 bit_16_10 bit_16_11 R_bl
Rbb_16_10 bitb_16_10 bitb_16_11 R_bl
Cb_16_10 bit_16_10 gnd C_bl
Cbb_16_10 bitb_16_10 gnd C_bl
Rb_16_11 bit_16_11 bit_16_12 R_bl
Rbb_16_11 bitb_16_11 bitb_16_12 R_bl
Cb_16_11 bit_16_11 gnd C_bl
Cbb_16_11 bitb_16_11 gnd C_bl
Rb_16_12 bit_16_12 bit_16_13 R_bl
Rbb_16_12 bitb_16_12 bitb_16_13 R_bl
Cb_16_12 bit_16_12 gnd C_bl
Cbb_16_12 bitb_16_12 gnd C_bl
Rb_16_13 bit_16_13 bit_16_14 R_bl
Rbb_16_13 bitb_16_13 bitb_16_14 R_bl
Cb_16_13 bit_16_13 gnd C_bl
Cbb_16_13 bitb_16_13 gnd C_bl
Rb_16_14 bit_16_14 bit_16_15 R_bl
Rbb_16_14 bitb_16_14 bitb_16_15 R_bl
Cb_16_14 bit_16_14 gnd C_bl
Cbb_16_14 bitb_16_14 gnd C_bl
Rb_16_15 bit_16_15 bit_16_16 R_bl
Rbb_16_15 bitb_16_15 bitb_16_16 R_bl
Cb_16_15 bit_16_15 gnd C_bl
Cbb_16_15 bitb_16_15 gnd C_bl
Rb_16_16 bit_16_16 bit_16_17 R_bl
Rbb_16_16 bitb_16_16 bitb_16_17 R_bl
Cb_16_16 bit_16_16 gnd C_bl
Cbb_16_16 bitb_16_16 gnd C_bl
Rb_16_17 bit_16_17 bit_16_18 R_bl
Rbb_16_17 bitb_16_17 bitb_16_18 R_bl
Cb_16_17 bit_16_17 gnd C_bl
Cbb_16_17 bitb_16_17 gnd C_bl
Rb_16_18 bit_16_18 bit_16_19 R_bl
Rbb_16_18 bitb_16_18 bitb_16_19 R_bl
Cb_16_18 bit_16_18 gnd C_bl
Cbb_16_18 bitb_16_18 gnd C_bl
Rb_16_19 bit_16_19 bit_16_20 R_bl
Rbb_16_19 bitb_16_19 bitb_16_20 R_bl
Cb_16_19 bit_16_19 gnd C_bl
Cbb_16_19 bitb_16_19 gnd C_bl
Rb_16_20 bit_16_20 bit_16_21 R_bl
Rbb_16_20 bitb_16_20 bitb_16_21 R_bl
Cb_16_20 bit_16_20 gnd C_bl
Cbb_16_20 bitb_16_20 gnd C_bl
Rb_16_21 bit_16_21 bit_16_22 R_bl
Rbb_16_21 bitb_16_21 bitb_16_22 R_bl
Cb_16_21 bit_16_21 gnd C_bl
Cbb_16_21 bitb_16_21 gnd C_bl
Rb_16_22 bit_16_22 bit_16_23 R_bl
Rbb_16_22 bitb_16_22 bitb_16_23 R_bl
Cb_16_22 bit_16_22 gnd C_bl
Cbb_16_22 bitb_16_22 gnd C_bl
Rb_16_23 bit_16_23 bit_16_24 R_bl
Rbb_16_23 bitb_16_23 bitb_16_24 R_bl
Cb_16_23 bit_16_23 gnd C_bl
Cbb_16_23 bitb_16_23 gnd C_bl
Rb_16_24 bit_16_24 bit_16_25 R_bl
Rbb_16_24 bitb_16_24 bitb_16_25 R_bl
Cb_16_24 bit_16_24 gnd C_bl
Cbb_16_24 bitb_16_24 gnd C_bl
Rb_16_25 bit_16_25 bit_16_26 R_bl
Rbb_16_25 bitb_16_25 bitb_16_26 R_bl
Cb_16_25 bit_16_25 gnd C_bl
Cbb_16_25 bitb_16_25 gnd C_bl
Rb_16_26 bit_16_26 bit_16_27 R_bl
Rbb_16_26 bitb_16_26 bitb_16_27 R_bl
Cb_16_26 bit_16_26 gnd C_bl
Cbb_16_26 bitb_16_26 gnd C_bl
Rb_16_27 bit_16_27 bit_16_28 R_bl
Rbb_16_27 bitb_16_27 bitb_16_28 R_bl
Cb_16_27 bit_16_27 gnd C_bl
Cbb_16_27 bitb_16_27 gnd C_bl
Rb_16_28 bit_16_28 bit_16_29 R_bl
Rbb_16_28 bitb_16_28 bitb_16_29 R_bl
Cb_16_28 bit_16_28 gnd C_bl
Cbb_16_28 bitb_16_28 gnd C_bl
Rb_16_29 bit_16_29 bit_16_30 R_bl
Rbb_16_29 bitb_16_29 bitb_16_30 R_bl
Cb_16_29 bit_16_29 gnd C_bl
Cbb_16_29 bitb_16_29 gnd C_bl
Rb_16_30 bit_16_30 bit_16_31 R_bl
Rbb_16_30 bitb_16_30 bitb_16_31 R_bl
Cb_16_30 bit_16_30 gnd C_bl
Cbb_16_30 bitb_16_30 gnd C_bl
Rb_16_31 bit_16_31 bit_16_32 R_bl
Rbb_16_31 bitb_16_31 bitb_16_32 R_bl
Cb_16_31 bit_16_31 gnd C_bl
Cbb_16_31 bitb_16_31 gnd C_bl
Rb_16_32 bit_16_32 bit_16_33 R_bl
Rbb_16_32 bitb_16_32 bitb_16_33 R_bl
Cb_16_32 bit_16_32 gnd C_bl
Cbb_16_32 bitb_16_32 gnd C_bl
Rb_16_33 bit_16_33 bit_16_34 R_bl
Rbb_16_33 bitb_16_33 bitb_16_34 R_bl
Cb_16_33 bit_16_33 gnd C_bl
Cbb_16_33 bitb_16_33 gnd C_bl
Rb_16_34 bit_16_34 bit_16_35 R_bl
Rbb_16_34 bitb_16_34 bitb_16_35 R_bl
Cb_16_34 bit_16_34 gnd C_bl
Cbb_16_34 bitb_16_34 gnd C_bl
Rb_16_35 bit_16_35 bit_16_36 R_bl
Rbb_16_35 bitb_16_35 bitb_16_36 R_bl
Cb_16_35 bit_16_35 gnd C_bl
Cbb_16_35 bitb_16_35 gnd C_bl
Rb_16_36 bit_16_36 bit_16_37 R_bl
Rbb_16_36 bitb_16_36 bitb_16_37 R_bl
Cb_16_36 bit_16_36 gnd C_bl
Cbb_16_36 bitb_16_36 gnd C_bl
Rb_16_37 bit_16_37 bit_16_38 R_bl
Rbb_16_37 bitb_16_37 bitb_16_38 R_bl
Cb_16_37 bit_16_37 gnd C_bl
Cbb_16_37 bitb_16_37 gnd C_bl
Rb_16_38 bit_16_38 bit_16_39 R_bl
Rbb_16_38 bitb_16_38 bitb_16_39 R_bl
Cb_16_38 bit_16_38 gnd C_bl
Cbb_16_38 bitb_16_38 gnd C_bl
Rb_16_39 bit_16_39 bit_16_40 R_bl
Rbb_16_39 bitb_16_39 bitb_16_40 R_bl
Cb_16_39 bit_16_39 gnd C_bl
Cbb_16_39 bitb_16_39 gnd C_bl
Rb_16_40 bit_16_40 bit_16_41 R_bl
Rbb_16_40 bitb_16_40 bitb_16_41 R_bl
Cb_16_40 bit_16_40 gnd C_bl
Cbb_16_40 bitb_16_40 gnd C_bl
Rb_16_41 bit_16_41 bit_16_42 R_bl
Rbb_16_41 bitb_16_41 bitb_16_42 R_bl
Cb_16_41 bit_16_41 gnd C_bl
Cbb_16_41 bitb_16_41 gnd C_bl
Rb_16_42 bit_16_42 bit_16_43 R_bl
Rbb_16_42 bitb_16_42 bitb_16_43 R_bl
Cb_16_42 bit_16_42 gnd C_bl
Cbb_16_42 bitb_16_42 gnd C_bl
Rb_16_43 bit_16_43 bit_16_44 R_bl
Rbb_16_43 bitb_16_43 bitb_16_44 R_bl
Cb_16_43 bit_16_43 gnd C_bl
Cbb_16_43 bitb_16_43 gnd C_bl
Rb_16_44 bit_16_44 bit_16_45 R_bl
Rbb_16_44 bitb_16_44 bitb_16_45 R_bl
Cb_16_44 bit_16_44 gnd C_bl
Cbb_16_44 bitb_16_44 gnd C_bl
Rb_16_45 bit_16_45 bit_16_46 R_bl
Rbb_16_45 bitb_16_45 bitb_16_46 R_bl
Cb_16_45 bit_16_45 gnd C_bl
Cbb_16_45 bitb_16_45 gnd C_bl
Rb_16_46 bit_16_46 bit_16_47 R_bl
Rbb_16_46 bitb_16_46 bitb_16_47 R_bl
Cb_16_46 bit_16_46 gnd C_bl
Cbb_16_46 bitb_16_46 gnd C_bl
Rb_16_47 bit_16_47 bit_16_48 R_bl
Rbb_16_47 bitb_16_47 bitb_16_48 R_bl
Cb_16_47 bit_16_47 gnd C_bl
Cbb_16_47 bitb_16_47 gnd C_bl
Rb_16_48 bit_16_48 bit_16_49 R_bl
Rbb_16_48 bitb_16_48 bitb_16_49 R_bl
Cb_16_48 bit_16_48 gnd C_bl
Cbb_16_48 bitb_16_48 gnd C_bl
Rb_16_49 bit_16_49 bit_16_50 R_bl
Rbb_16_49 bitb_16_49 bitb_16_50 R_bl
Cb_16_49 bit_16_49 gnd C_bl
Cbb_16_49 bitb_16_49 gnd C_bl
Rb_16_50 bit_16_50 bit_16_51 R_bl
Rbb_16_50 bitb_16_50 bitb_16_51 R_bl
Cb_16_50 bit_16_50 gnd C_bl
Cbb_16_50 bitb_16_50 gnd C_bl
Rb_16_51 bit_16_51 bit_16_52 R_bl
Rbb_16_51 bitb_16_51 bitb_16_52 R_bl
Cb_16_51 bit_16_51 gnd C_bl
Cbb_16_51 bitb_16_51 gnd C_bl
Rb_16_52 bit_16_52 bit_16_53 R_bl
Rbb_16_52 bitb_16_52 bitb_16_53 R_bl
Cb_16_52 bit_16_52 gnd C_bl
Cbb_16_52 bitb_16_52 gnd C_bl
Rb_16_53 bit_16_53 bit_16_54 R_bl
Rbb_16_53 bitb_16_53 bitb_16_54 R_bl
Cb_16_53 bit_16_53 gnd C_bl
Cbb_16_53 bitb_16_53 gnd C_bl
Rb_16_54 bit_16_54 bit_16_55 R_bl
Rbb_16_54 bitb_16_54 bitb_16_55 R_bl
Cb_16_54 bit_16_54 gnd C_bl
Cbb_16_54 bitb_16_54 gnd C_bl
Rb_16_55 bit_16_55 bit_16_56 R_bl
Rbb_16_55 bitb_16_55 bitb_16_56 R_bl
Cb_16_55 bit_16_55 gnd C_bl
Cbb_16_55 bitb_16_55 gnd C_bl
Rb_16_56 bit_16_56 bit_16_57 R_bl
Rbb_16_56 bitb_16_56 bitb_16_57 R_bl
Cb_16_56 bit_16_56 gnd C_bl
Cbb_16_56 bitb_16_56 gnd C_bl
Rb_16_57 bit_16_57 bit_16_58 R_bl
Rbb_16_57 bitb_16_57 bitb_16_58 R_bl
Cb_16_57 bit_16_57 gnd C_bl
Cbb_16_57 bitb_16_57 gnd C_bl
Rb_16_58 bit_16_58 bit_16_59 R_bl
Rbb_16_58 bitb_16_58 bitb_16_59 R_bl
Cb_16_58 bit_16_58 gnd C_bl
Cbb_16_58 bitb_16_58 gnd C_bl
Rb_16_59 bit_16_59 bit_16_60 R_bl
Rbb_16_59 bitb_16_59 bitb_16_60 R_bl
Cb_16_59 bit_16_59 gnd C_bl
Cbb_16_59 bitb_16_59 gnd C_bl
Rb_16_60 bit_16_60 bit_16_61 R_bl
Rbb_16_60 bitb_16_60 bitb_16_61 R_bl
Cb_16_60 bit_16_60 gnd C_bl
Cbb_16_60 bitb_16_60 gnd C_bl
Rb_16_61 bit_16_61 bit_16_62 R_bl
Rbb_16_61 bitb_16_61 bitb_16_62 R_bl
Cb_16_61 bit_16_61 gnd C_bl
Cbb_16_61 bitb_16_61 gnd C_bl
Rb_16_62 bit_16_62 bit_16_63 R_bl
Rbb_16_62 bitb_16_62 bitb_16_63 R_bl
Cb_16_62 bit_16_62 gnd C_bl
Cbb_16_62 bitb_16_62 gnd C_bl
Rb_16_63 bit_16_63 bit_16_64 R_bl
Rbb_16_63 bitb_16_63 bitb_16_64 R_bl
Cb_16_63 bit_16_63 gnd C_bl
Cbb_16_63 bitb_16_63 gnd C_bl
Rb_16_64 bit_16_64 bit_16_65 R_bl
Rbb_16_64 bitb_16_64 bitb_16_65 R_bl
Cb_16_64 bit_16_64 gnd C_bl
Cbb_16_64 bitb_16_64 gnd C_bl
Rb_16_65 bit_16_65 bit_16_66 R_bl
Rbb_16_65 bitb_16_65 bitb_16_66 R_bl
Cb_16_65 bit_16_65 gnd C_bl
Cbb_16_65 bitb_16_65 gnd C_bl
Rb_16_66 bit_16_66 bit_16_67 R_bl
Rbb_16_66 bitb_16_66 bitb_16_67 R_bl
Cb_16_66 bit_16_66 gnd C_bl
Cbb_16_66 bitb_16_66 gnd C_bl
Rb_16_67 bit_16_67 bit_16_68 R_bl
Rbb_16_67 bitb_16_67 bitb_16_68 R_bl
Cb_16_67 bit_16_67 gnd C_bl
Cbb_16_67 bitb_16_67 gnd C_bl
Rb_16_68 bit_16_68 bit_16_69 R_bl
Rbb_16_68 bitb_16_68 bitb_16_69 R_bl
Cb_16_68 bit_16_68 gnd C_bl
Cbb_16_68 bitb_16_68 gnd C_bl
Rb_16_69 bit_16_69 bit_16_70 R_bl
Rbb_16_69 bitb_16_69 bitb_16_70 R_bl
Cb_16_69 bit_16_69 gnd C_bl
Cbb_16_69 bitb_16_69 gnd C_bl
Rb_16_70 bit_16_70 bit_16_71 R_bl
Rbb_16_70 bitb_16_70 bitb_16_71 R_bl
Cb_16_70 bit_16_70 gnd C_bl
Cbb_16_70 bitb_16_70 gnd C_bl
Rb_16_71 bit_16_71 bit_16_72 R_bl
Rbb_16_71 bitb_16_71 bitb_16_72 R_bl
Cb_16_71 bit_16_71 gnd C_bl
Cbb_16_71 bitb_16_71 gnd C_bl
Rb_16_72 bit_16_72 bit_16_73 R_bl
Rbb_16_72 bitb_16_72 bitb_16_73 R_bl
Cb_16_72 bit_16_72 gnd C_bl
Cbb_16_72 bitb_16_72 gnd C_bl
Rb_16_73 bit_16_73 bit_16_74 R_bl
Rbb_16_73 bitb_16_73 bitb_16_74 R_bl
Cb_16_73 bit_16_73 gnd C_bl
Cbb_16_73 bitb_16_73 gnd C_bl
Rb_16_74 bit_16_74 bit_16_75 R_bl
Rbb_16_74 bitb_16_74 bitb_16_75 R_bl
Cb_16_74 bit_16_74 gnd C_bl
Cbb_16_74 bitb_16_74 gnd C_bl
Rb_16_75 bit_16_75 bit_16_76 R_bl
Rbb_16_75 bitb_16_75 bitb_16_76 R_bl
Cb_16_75 bit_16_75 gnd C_bl
Cbb_16_75 bitb_16_75 gnd C_bl
Rb_16_76 bit_16_76 bit_16_77 R_bl
Rbb_16_76 bitb_16_76 bitb_16_77 R_bl
Cb_16_76 bit_16_76 gnd C_bl
Cbb_16_76 bitb_16_76 gnd C_bl
Rb_16_77 bit_16_77 bit_16_78 R_bl
Rbb_16_77 bitb_16_77 bitb_16_78 R_bl
Cb_16_77 bit_16_77 gnd C_bl
Cbb_16_77 bitb_16_77 gnd C_bl
Rb_16_78 bit_16_78 bit_16_79 R_bl
Rbb_16_78 bitb_16_78 bitb_16_79 R_bl
Cb_16_78 bit_16_78 gnd C_bl
Cbb_16_78 bitb_16_78 gnd C_bl
Rb_16_79 bit_16_79 bit_16_80 R_bl
Rbb_16_79 bitb_16_79 bitb_16_80 R_bl
Cb_16_79 bit_16_79 gnd C_bl
Cbb_16_79 bitb_16_79 gnd C_bl
Rb_16_80 bit_16_80 bit_16_81 R_bl
Rbb_16_80 bitb_16_80 bitb_16_81 R_bl
Cb_16_80 bit_16_80 gnd C_bl
Cbb_16_80 bitb_16_80 gnd C_bl
Rb_16_81 bit_16_81 bit_16_82 R_bl
Rbb_16_81 bitb_16_81 bitb_16_82 R_bl
Cb_16_81 bit_16_81 gnd C_bl
Cbb_16_81 bitb_16_81 gnd C_bl
Rb_16_82 bit_16_82 bit_16_83 R_bl
Rbb_16_82 bitb_16_82 bitb_16_83 R_bl
Cb_16_82 bit_16_82 gnd C_bl
Cbb_16_82 bitb_16_82 gnd C_bl
Rb_16_83 bit_16_83 bit_16_84 R_bl
Rbb_16_83 bitb_16_83 bitb_16_84 R_bl
Cb_16_83 bit_16_83 gnd C_bl
Cbb_16_83 bitb_16_83 gnd C_bl
Rb_16_84 bit_16_84 bit_16_85 R_bl
Rbb_16_84 bitb_16_84 bitb_16_85 R_bl
Cb_16_84 bit_16_84 gnd C_bl
Cbb_16_84 bitb_16_84 gnd C_bl
Rb_16_85 bit_16_85 bit_16_86 R_bl
Rbb_16_85 bitb_16_85 bitb_16_86 R_bl
Cb_16_85 bit_16_85 gnd C_bl
Cbb_16_85 bitb_16_85 gnd C_bl
Rb_16_86 bit_16_86 bit_16_87 R_bl
Rbb_16_86 bitb_16_86 bitb_16_87 R_bl
Cb_16_86 bit_16_86 gnd C_bl
Cbb_16_86 bitb_16_86 gnd C_bl
Rb_16_87 bit_16_87 bit_16_88 R_bl
Rbb_16_87 bitb_16_87 bitb_16_88 R_bl
Cb_16_87 bit_16_87 gnd C_bl
Cbb_16_87 bitb_16_87 gnd C_bl
Rb_16_88 bit_16_88 bit_16_89 R_bl
Rbb_16_88 bitb_16_88 bitb_16_89 R_bl
Cb_16_88 bit_16_88 gnd C_bl
Cbb_16_88 bitb_16_88 gnd C_bl
Rb_16_89 bit_16_89 bit_16_90 R_bl
Rbb_16_89 bitb_16_89 bitb_16_90 R_bl
Cb_16_89 bit_16_89 gnd C_bl
Cbb_16_89 bitb_16_89 gnd C_bl
Rb_16_90 bit_16_90 bit_16_91 R_bl
Rbb_16_90 bitb_16_90 bitb_16_91 R_bl
Cb_16_90 bit_16_90 gnd C_bl
Cbb_16_90 bitb_16_90 gnd C_bl
Rb_16_91 bit_16_91 bit_16_92 R_bl
Rbb_16_91 bitb_16_91 bitb_16_92 R_bl
Cb_16_91 bit_16_91 gnd C_bl
Cbb_16_91 bitb_16_91 gnd C_bl
Rb_16_92 bit_16_92 bit_16_93 R_bl
Rbb_16_92 bitb_16_92 bitb_16_93 R_bl
Cb_16_92 bit_16_92 gnd C_bl
Cbb_16_92 bitb_16_92 gnd C_bl
Rb_16_93 bit_16_93 bit_16_94 R_bl
Rbb_16_93 bitb_16_93 bitb_16_94 R_bl
Cb_16_93 bit_16_93 gnd C_bl
Cbb_16_93 bitb_16_93 gnd C_bl
Rb_16_94 bit_16_94 bit_16_95 R_bl
Rbb_16_94 bitb_16_94 bitb_16_95 R_bl
Cb_16_94 bit_16_94 gnd C_bl
Cbb_16_94 bitb_16_94 gnd C_bl
Rb_16_95 bit_16_95 bit_16_96 R_bl
Rbb_16_95 bitb_16_95 bitb_16_96 R_bl
Cb_16_95 bit_16_95 gnd C_bl
Cbb_16_95 bitb_16_95 gnd C_bl
Rb_16_96 bit_16_96 bit_16_97 R_bl
Rbb_16_96 bitb_16_96 bitb_16_97 R_bl
Cb_16_96 bit_16_96 gnd C_bl
Cbb_16_96 bitb_16_96 gnd C_bl
Rb_16_97 bit_16_97 bit_16_98 R_bl
Rbb_16_97 bitb_16_97 bitb_16_98 R_bl
Cb_16_97 bit_16_97 gnd C_bl
Cbb_16_97 bitb_16_97 gnd C_bl
Rb_16_98 bit_16_98 bit_16_99 R_bl
Rbb_16_98 bitb_16_98 bitb_16_99 R_bl
Cb_16_98 bit_16_98 gnd C_bl
Cbb_16_98 bitb_16_98 gnd C_bl
Rb_16_99 bit_16_99 bit_16_100 R_bl
Rbb_16_99 bitb_16_99 bitb_16_100 R_bl
Cb_16_99 bit_16_99 gnd C_bl
Cbb_16_99 bitb_16_99 gnd C_bl
Rb_17_0 bit_17_0 bit_17_1 R_bl
Rbb_17_0 bitb_17_0 bitb_17_1 R_bl
Cb_17_0 bit_17_0 gnd C_bl
Cbb_17_0 bitb_17_0 gnd C_bl
Rb_17_1 bit_17_1 bit_17_2 R_bl
Rbb_17_1 bitb_17_1 bitb_17_2 R_bl
Cb_17_1 bit_17_1 gnd C_bl
Cbb_17_1 bitb_17_1 gnd C_bl
Rb_17_2 bit_17_2 bit_17_3 R_bl
Rbb_17_2 bitb_17_2 bitb_17_3 R_bl
Cb_17_2 bit_17_2 gnd C_bl
Cbb_17_2 bitb_17_2 gnd C_bl
Rb_17_3 bit_17_3 bit_17_4 R_bl
Rbb_17_3 bitb_17_3 bitb_17_4 R_bl
Cb_17_3 bit_17_3 gnd C_bl
Cbb_17_3 bitb_17_3 gnd C_bl
Rb_17_4 bit_17_4 bit_17_5 R_bl
Rbb_17_4 bitb_17_4 bitb_17_5 R_bl
Cb_17_4 bit_17_4 gnd C_bl
Cbb_17_4 bitb_17_4 gnd C_bl
Rb_17_5 bit_17_5 bit_17_6 R_bl
Rbb_17_5 bitb_17_5 bitb_17_6 R_bl
Cb_17_5 bit_17_5 gnd C_bl
Cbb_17_5 bitb_17_5 gnd C_bl
Rb_17_6 bit_17_6 bit_17_7 R_bl
Rbb_17_6 bitb_17_6 bitb_17_7 R_bl
Cb_17_6 bit_17_6 gnd C_bl
Cbb_17_6 bitb_17_6 gnd C_bl
Rb_17_7 bit_17_7 bit_17_8 R_bl
Rbb_17_7 bitb_17_7 bitb_17_8 R_bl
Cb_17_7 bit_17_7 gnd C_bl
Cbb_17_7 bitb_17_7 gnd C_bl
Rb_17_8 bit_17_8 bit_17_9 R_bl
Rbb_17_8 bitb_17_8 bitb_17_9 R_bl
Cb_17_8 bit_17_8 gnd C_bl
Cbb_17_8 bitb_17_8 gnd C_bl
Rb_17_9 bit_17_9 bit_17_10 R_bl
Rbb_17_9 bitb_17_9 bitb_17_10 R_bl
Cb_17_9 bit_17_9 gnd C_bl
Cbb_17_9 bitb_17_9 gnd C_bl
Rb_17_10 bit_17_10 bit_17_11 R_bl
Rbb_17_10 bitb_17_10 bitb_17_11 R_bl
Cb_17_10 bit_17_10 gnd C_bl
Cbb_17_10 bitb_17_10 gnd C_bl
Rb_17_11 bit_17_11 bit_17_12 R_bl
Rbb_17_11 bitb_17_11 bitb_17_12 R_bl
Cb_17_11 bit_17_11 gnd C_bl
Cbb_17_11 bitb_17_11 gnd C_bl
Rb_17_12 bit_17_12 bit_17_13 R_bl
Rbb_17_12 bitb_17_12 bitb_17_13 R_bl
Cb_17_12 bit_17_12 gnd C_bl
Cbb_17_12 bitb_17_12 gnd C_bl
Rb_17_13 bit_17_13 bit_17_14 R_bl
Rbb_17_13 bitb_17_13 bitb_17_14 R_bl
Cb_17_13 bit_17_13 gnd C_bl
Cbb_17_13 bitb_17_13 gnd C_bl
Rb_17_14 bit_17_14 bit_17_15 R_bl
Rbb_17_14 bitb_17_14 bitb_17_15 R_bl
Cb_17_14 bit_17_14 gnd C_bl
Cbb_17_14 bitb_17_14 gnd C_bl
Rb_17_15 bit_17_15 bit_17_16 R_bl
Rbb_17_15 bitb_17_15 bitb_17_16 R_bl
Cb_17_15 bit_17_15 gnd C_bl
Cbb_17_15 bitb_17_15 gnd C_bl
Rb_17_16 bit_17_16 bit_17_17 R_bl
Rbb_17_16 bitb_17_16 bitb_17_17 R_bl
Cb_17_16 bit_17_16 gnd C_bl
Cbb_17_16 bitb_17_16 gnd C_bl
Rb_17_17 bit_17_17 bit_17_18 R_bl
Rbb_17_17 bitb_17_17 bitb_17_18 R_bl
Cb_17_17 bit_17_17 gnd C_bl
Cbb_17_17 bitb_17_17 gnd C_bl
Rb_17_18 bit_17_18 bit_17_19 R_bl
Rbb_17_18 bitb_17_18 bitb_17_19 R_bl
Cb_17_18 bit_17_18 gnd C_bl
Cbb_17_18 bitb_17_18 gnd C_bl
Rb_17_19 bit_17_19 bit_17_20 R_bl
Rbb_17_19 bitb_17_19 bitb_17_20 R_bl
Cb_17_19 bit_17_19 gnd C_bl
Cbb_17_19 bitb_17_19 gnd C_bl
Rb_17_20 bit_17_20 bit_17_21 R_bl
Rbb_17_20 bitb_17_20 bitb_17_21 R_bl
Cb_17_20 bit_17_20 gnd C_bl
Cbb_17_20 bitb_17_20 gnd C_bl
Rb_17_21 bit_17_21 bit_17_22 R_bl
Rbb_17_21 bitb_17_21 bitb_17_22 R_bl
Cb_17_21 bit_17_21 gnd C_bl
Cbb_17_21 bitb_17_21 gnd C_bl
Rb_17_22 bit_17_22 bit_17_23 R_bl
Rbb_17_22 bitb_17_22 bitb_17_23 R_bl
Cb_17_22 bit_17_22 gnd C_bl
Cbb_17_22 bitb_17_22 gnd C_bl
Rb_17_23 bit_17_23 bit_17_24 R_bl
Rbb_17_23 bitb_17_23 bitb_17_24 R_bl
Cb_17_23 bit_17_23 gnd C_bl
Cbb_17_23 bitb_17_23 gnd C_bl
Rb_17_24 bit_17_24 bit_17_25 R_bl
Rbb_17_24 bitb_17_24 bitb_17_25 R_bl
Cb_17_24 bit_17_24 gnd C_bl
Cbb_17_24 bitb_17_24 gnd C_bl
Rb_17_25 bit_17_25 bit_17_26 R_bl
Rbb_17_25 bitb_17_25 bitb_17_26 R_bl
Cb_17_25 bit_17_25 gnd C_bl
Cbb_17_25 bitb_17_25 gnd C_bl
Rb_17_26 bit_17_26 bit_17_27 R_bl
Rbb_17_26 bitb_17_26 bitb_17_27 R_bl
Cb_17_26 bit_17_26 gnd C_bl
Cbb_17_26 bitb_17_26 gnd C_bl
Rb_17_27 bit_17_27 bit_17_28 R_bl
Rbb_17_27 bitb_17_27 bitb_17_28 R_bl
Cb_17_27 bit_17_27 gnd C_bl
Cbb_17_27 bitb_17_27 gnd C_bl
Rb_17_28 bit_17_28 bit_17_29 R_bl
Rbb_17_28 bitb_17_28 bitb_17_29 R_bl
Cb_17_28 bit_17_28 gnd C_bl
Cbb_17_28 bitb_17_28 gnd C_bl
Rb_17_29 bit_17_29 bit_17_30 R_bl
Rbb_17_29 bitb_17_29 bitb_17_30 R_bl
Cb_17_29 bit_17_29 gnd C_bl
Cbb_17_29 bitb_17_29 gnd C_bl
Rb_17_30 bit_17_30 bit_17_31 R_bl
Rbb_17_30 bitb_17_30 bitb_17_31 R_bl
Cb_17_30 bit_17_30 gnd C_bl
Cbb_17_30 bitb_17_30 gnd C_bl
Rb_17_31 bit_17_31 bit_17_32 R_bl
Rbb_17_31 bitb_17_31 bitb_17_32 R_bl
Cb_17_31 bit_17_31 gnd C_bl
Cbb_17_31 bitb_17_31 gnd C_bl
Rb_17_32 bit_17_32 bit_17_33 R_bl
Rbb_17_32 bitb_17_32 bitb_17_33 R_bl
Cb_17_32 bit_17_32 gnd C_bl
Cbb_17_32 bitb_17_32 gnd C_bl
Rb_17_33 bit_17_33 bit_17_34 R_bl
Rbb_17_33 bitb_17_33 bitb_17_34 R_bl
Cb_17_33 bit_17_33 gnd C_bl
Cbb_17_33 bitb_17_33 gnd C_bl
Rb_17_34 bit_17_34 bit_17_35 R_bl
Rbb_17_34 bitb_17_34 bitb_17_35 R_bl
Cb_17_34 bit_17_34 gnd C_bl
Cbb_17_34 bitb_17_34 gnd C_bl
Rb_17_35 bit_17_35 bit_17_36 R_bl
Rbb_17_35 bitb_17_35 bitb_17_36 R_bl
Cb_17_35 bit_17_35 gnd C_bl
Cbb_17_35 bitb_17_35 gnd C_bl
Rb_17_36 bit_17_36 bit_17_37 R_bl
Rbb_17_36 bitb_17_36 bitb_17_37 R_bl
Cb_17_36 bit_17_36 gnd C_bl
Cbb_17_36 bitb_17_36 gnd C_bl
Rb_17_37 bit_17_37 bit_17_38 R_bl
Rbb_17_37 bitb_17_37 bitb_17_38 R_bl
Cb_17_37 bit_17_37 gnd C_bl
Cbb_17_37 bitb_17_37 gnd C_bl
Rb_17_38 bit_17_38 bit_17_39 R_bl
Rbb_17_38 bitb_17_38 bitb_17_39 R_bl
Cb_17_38 bit_17_38 gnd C_bl
Cbb_17_38 bitb_17_38 gnd C_bl
Rb_17_39 bit_17_39 bit_17_40 R_bl
Rbb_17_39 bitb_17_39 bitb_17_40 R_bl
Cb_17_39 bit_17_39 gnd C_bl
Cbb_17_39 bitb_17_39 gnd C_bl
Rb_17_40 bit_17_40 bit_17_41 R_bl
Rbb_17_40 bitb_17_40 bitb_17_41 R_bl
Cb_17_40 bit_17_40 gnd C_bl
Cbb_17_40 bitb_17_40 gnd C_bl
Rb_17_41 bit_17_41 bit_17_42 R_bl
Rbb_17_41 bitb_17_41 bitb_17_42 R_bl
Cb_17_41 bit_17_41 gnd C_bl
Cbb_17_41 bitb_17_41 gnd C_bl
Rb_17_42 bit_17_42 bit_17_43 R_bl
Rbb_17_42 bitb_17_42 bitb_17_43 R_bl
Cb_17_42 bit_17_42 gnd C_bl
Cbb_17_42 bitb_17_42 gnd C_bl
Rb_17_43 bit_17_43 bit_17_44 R_bl
Rbb_17_43 bitb_17_43 bitb_17_44 R_bl
Cb_17_43 bit_17_43 gnd C_bl
Cbb_17_43 bitb_17_43 gnd C_bl
Rb_17_44 bit_17_44 bit_17_45 R_bl
Rbb_17_44 bitb_17_44 bitb_17_45 R_bl
Cb_17_44 bit_17_44 gnd C_bl
Cbb_17_44 bitb_17_44 gnd C_bl
Rb_17_45 bit_17_45 bit_17_46 R_bl
Rbb_17_45 bitb_17_45 bitb_17_46 R_bl
Cb_17_45 bit_17_45 gnd C_bl
Cbb_17_45 bitb_17_45 gnd C_bl
Rb_17_46 bit_17_46 bit_17_47 R_bl
Rbb_17_46 bitb_17_46 bitb_17_47 R_bl
Cb_17_46 bit_17_46 gnd C_bl
Cbb_17_46 bitb_17_46 gnd C_bl
Rb_17_47 bit_17_47 bit_17_48 R_bl
Rbb_17_47 bitb_17_47 bitb_17_48 R_bl
Cb_17_47 bit_17_47 gnd C_bl
Cbb_17_47 bitb_17_47 gnd C_bl
Rb_17_48 bit_17_48 bit_17_49 R_bl
Rbb_17_48 bitb_17_48 bitb_17_49 R_bl
Cb_17_48 bit_17_48 gnd C_bl
Cbb_17_48 bitb_17_48 gnd C_bl
Rb_17_49 bit_17_49 bit_17_50 R_bl
Rbb_17_49 bitb_17_49 bitb_17_50 R_bl
Cb_17_49 bit_17_49 gnd C_bl
Cbb_17_49 bitb_17_49 gnd C_bl
Rb_17_50 bit_17_50 bit_17_51 R_bl
Rbb_17_50 bitb_17_50 bitb_17_51 R_bl
Cb_17_50 bit_17_50 gnd C_bl
Cbb_17_50 bitb_17_50 gnd C_bl
Rb_17_51 bit_17_51 bit_17_52 R_bl
Rbb_17_51 bitb_17_51 bitb_17_52 R_bl
Cb_17_51 bit_17_51 gnd C_bl
Cbb_17_51 bitb_17_51 gnd C_bl
Rb_17_52 bit_17_52 bit_17_53 R_bl
Rbb_17_52 bitb_17_52 bitb_17_53 R_bl
Cb_17_52 bit_17_52 gnd C_bl
Cbb_17_52 bitb_17_52 gnd C_bl
Rb_17_53 bit_17_53 bit_17_54 R_bl
Rbb_17_53 bitb_17_53 bitb_17_54 R_bl
Cb_17_53 bit_17_53 gnd C_bl
Cbb_17_53 bitb_17_53 gnd C_bl
Rb_17_54 bit_17_54 bit_17_55 R_bl
Rbb_17_54 bitb_17_54 bitb_17_55 R_bl
Cb_17_54 bit_17_54 gnd C_bl
Cbb_17_54 bitb_17_54 gnd C_bl
Rb_17_55 bit_17_55 bit_17_56 R_bl
Rbb_17_55 bitb_17_55 bitb_17_56 R_bl
Cb_17_55 bit_17_55 gnd C_bl
Cbb_17_55 bitb_17_55 gnd C_bl
Rb_17_56 bit_17_56 bit_17_57 R_bl
Rbb_17_56 bitb_17_56 bitb_17_57 R_bl
Cb_17_56 bit_17_56 gnd C_bl
Cbb_17_56 bitb_17_56 gnd C_bl
Rb_17_57 bit_17_57 bit_17_58 R_bl
Rbb_17_57 bitb_17_57 bitb_17_58 R_bl
Cb_17_57 bit_17_57 gnd C_bl
Cbb_17_57 bitb_17_57 gnd C_bl
Rb_17_58 bit_17_58 bit_17_59 R_bl
Rbb_17_58 bitb_17_58 bitb_17_59 R_bl
Cb_17_58 bit_17_58 gnd C_bl
Cbb_17_58 bitb_17_58 gnd C_bl
Rb_17_59 bit_17_59 bit_17_60 R_bl
Rbb_17_59 bitb_17_59 bitb_17_60 R_bl
Cb_17_59 bit_17_59 gnd C_bl
Cbb_17_59 bitb_17_59 gnd C_bl
Rb_17_60 bit_17_60 bit_17_61 R_bl
Rbb_17_60 bitb_17_60 bitb_17_61 R_bl
Cb_17_60 bit_17_60 gnd C_bl
Cbb_17_60 bitb_17_60 gnd C_bl
Rb_17_61 bit_17_61 bit_17_62 R_bl
Rbb_17_61 bitb_17_61 bitb_17_62 R_bl
Cb_17_61 bit_17_61 gnd C_bl
Cbb_17_61 bitb_17_61 gnd C_bl
Rb_17_62 bit_17_62 bit_17_63 R_bl
Rbb_17_62 bitb_17_62 bitb_17_63 R_bl
Cb_17_62 bit_17_62 gnd C_bl
Cbb_17_62 bitb_17_62 gnd C_bl
Rb_17_63 bit_17_63 bit_17_64 R_bl
Rbb_17_63 bitb_17_63 bitb_17_64 R_bl
Cb_17_63 bit_17_63 gnd C_bl
Cbb_17_63 bitb_17_63 gnd C_bl
Rb_17_64 bit_17_64 bit_17_65 R_bl
Rbb_17_64 bitb_17_64 bitb_17_65 R_bl
Cb_17_64 bit_17_64 gnd C_bl
Cbb_17_64 bitb_17_64 gnd C_bl
Rb_17_65 bit_17_65 bit_17_66 R_bl
Rbb_17_65 bitb_17_65 bitb_17_66 R_bl
Cb_17_65 bit_17_65 gnd C_bl
Cbb_17_65 bitb_17_65 gnd C_bl
Rb_17_66 bit_17_66 bit_17_67 R_bl
Rbb_17_66 bitb_17_66 bitb_17_67 R_bl
Cb_17_66 bit_17_66 gnd C_bl
Cbb_17_66 bitb_17_66 gnd C_bl
Rb_17_67 bit_17_67 bit_17_68 R_bl
Rbb_17_67 bitb_17_67 bitb_17_68 R_bl
Cb_17_67 bit_17_67 gnd C_bl
Cbb_17_67 bitb_17_67 gnd C_bl
Rb_17_68 bit_17_68 bit_17_69 R_bl
Rbb_17_68 bitb_17_68 bitb_17_69 R_bl
Cb_17_68 bit_17_68 gnd C_bl
Cbb_17_68 bitb_17_68 gnd C_bl
Rb_17_69 bit_17_69 bit_17_70 R_bl
Rbb_17_69 bitb_17_69 bitb_17_70 R_bl
Cb_17_69 bit_17_69 gnd C_bl
Cbb_17_69 bitb_17_69 gnd C_bl
Rb_17_70 bit_17_70 bit_17_71 R_bl
Rbb_17_70 bitb_17_70 bitb_17_71 R_bl
Cb_17_70 bit_17_70 gnd C_bl
Cbb_17_70 bitb_17_70 gnd C_bl
Rb_17_71 bit_17_71 bit_17_72 R_bl
Rbb_17_71 bitb_17_71 bitb_17_72 R_bl
Cb_17_71 bit_17_71 gnd C_bl
Cbb_17_71 bitb_17_71 gnd C_bl
Rb_17_72 bit_17_72 bit_17_73 R_bl
Rbb_17_72 bitb_17_72 bitb_17_73 R_bl
Cb_17_72 bit_17_72 gnd C_bl
Cbb_17_72 bitb_17_72 gnd C_bl
Rb_17_73 bit_17_73 bit_17_74 R_bl
Rbb_17_73 bitb_17_73 bitb_17_74 R_bl
Cb_17_73 bit_17_73 gnd C_bl
Cbb_17_73 bitb_17_73 gnd C_bl
Rb_17_74 bit_17_74 bit_17_75 R_bl
Rbb_17_74 bitb_17_74 bitb_17_75 R_bl
Cb_17_74 bit_17_74 gnd C_bl
Cbb_17_74 bitb_17_74 gnd C_bl
Rb_17_75 bit_17_75 bit_17_76 R_bl
Rbb_17_75 bitb_17_75 bitb_17_76 R_bl
Cb_17_75 bit_17_75 gnd C_bl
Cbb_17_75 bitb_17_75 gnd C_bl
Rb_17_76 bit_17_76 bit_17_77 R_bl
Rbb_17_76 bitb_17_76 bitb_17_77 R_bl
Cb_17_76 bit_17_76 gnd C_bl
Cbb_17_76 bitb_17_76 gnd C_bl
Rb_17_77 bit_17_77 bit_17_78 R_bl
Rbb_17_77 bitb_17_77 bitb_17_78 R_bl
Cb_17_77 bit_17_77 gnd C_bl
Cbb_17_77 bitb_17_77 gnd C_bl
Rb_17_78 bit_17_78 bit_17_79 R_bl
Rbb_17_78 bitb_17_78 bitb_17_79 R_bl
Cb_17_78 bit_17_78 gnd C_bl
Cbb_17_78 bitb_17_78 gnd C_bl
Rb_17_79 bit_17_79 bit_17_80 R_bl
Rbb_17_79 bitb_17_79 bitb_17_80 R_bl
Cb_17_79 bit_17_79 gnd C_bl
Cbb_17_79 bitb_17_79 gnd C_bl
Rb_17_80 bit_17_80 bit_17_81 R_bl
Rbb_17_80 bitb_17_80 bitb_17_81 R_bl
Cb_17_80 bit_17_80 gnd C_bl
Cbb_17_80 bitb_17_80 gnd C_bl
Rb_17_81 bit_17_81 bit_17_82 R_bl
Rbb_17_81 bitb_17_81 bitb_17_82 R_bl
Cb_17_81 bit_17_81 gnd C_bl
Cbb_17_81 bitb_17_81 gnd C_bl
Rb_17_82 bit_17_82 bit_17_83 R_bl
Rbb_17_82 bitb_17_82 bitb_17_83 R_bl
Cb_17_82 bit_17_82 gnd C_bl
Cbb_17_82 bitb_17_82 gnd C_bl
Rb_17_83 bit_17_83 bit_17_84 R_bl
Rbb_17_83 bitb_17_83 bitb_17_84 R_bl
Cb_17_83 bit_17_83 gnd C_bl
Cbb_17_83 bitb_17_83 gnd C_bl
Rb_17_84 bit_17_84 bit_17_85 R_bl
Rbb_17_84 bitb_17_84 bitb_17_85 R_bl
Cb_17_84 bit_17_84 gnd C_bl
Cbb_17_84 bitb_17_84 gnd C_bl
Rb_17_85 bit_17_85 bit_17_86 R_bl
Rbb_17_85 bitb_17_85 bitb_17_86 R_bl
Cb_17_85 bit_17_85 gnd C_bl
Cbb_17_85 bitb_17_85 gnd C_bl
Rb_17_86 bit_17_86 bit_17_87 R_bl
Rbb_17_86 bitb_17_86 bitb_17_87 R_bl
Cb_17_86 bit_17_86 gnd C_bl
Cbb_17_86 bitb_17_86 gnd C_bl
Rb_17_87 bit_17_87 bit_17_88 R_bl
Rbb_17_87 bitb_17_87 bitb_17_88 R_bl
Cb_17_87 bit_17_87 gnd C_bl
Cbb_17_87 bitb_17_87 gnd C_bl
Rb_17_88 bit_17_88 bit_17_89 R_bl
Rbb_17_88 bitb_17_88 bitb_17_89 R_bl
Cb_17_88 bit_17_88 gnd C_bl
Cbb_17_88 bitb_17_88 gnd C_bl
Rb_17_89 bit_17_89 bit_17_90 R_bl
Rbb_17_89 bitb_17_89 bitb_17_90 R_bl
Cb_17_89 bit_17_89 gnd C_bl
Cbb_17_89 bitb_17_89 gnd C_bl
Rb_17_90 bit_17_90 bit_17_91 R_bl
Rbb_17_90 bitb_17_90 bitb_17_91 R_bl
Cb_17_90 bit_17_90 gnd C_bl
Cbb_17_90 bitb_17_90 gnd C_bl
Rb_17_91 bit_17_91 bit_17_92 R_bl
Rbb_17_91 bitb_17_91 bitb_17_92 R_bl
Cb_17_91 bit_17_91 gnd C_bl
Cbb_17_91 bitb_17_91 gnd C_bl
Rb_17_92 bit_17_92 bit_17_93 R_bl
Rbb_17_92 bitb_17_92 bitb_17_93 R_bl
Cb_17_92 bit_17_92 gnd C_bl
Cbb_17_92 bitb_17_92 gnd C_bl
Rb_17_93 bit_17_93 bit_17_94 R_bl
Rbb_17_93 bitb_17_93 bitb_17_94 R_bl
Cb_17_93 bit_17_93 gnd C_bl
Cbb_17_93 bitb_17_93 gnd C_bl
Rb_17_94 bit_17_94 bit_17_95 R_bl
Rbb_17_94 bitb_17_94 bitb_17_95 R_bl
Cb_17_94 bit_17_94 gnd C_bl
Cbb_17_94 bitb_17_94 gnd C_bl
Rb_17_95 bit_17_95 bit_17_96 R_bl
Rbb_17_95 bitb_17_95 bitb_17_96 R_bl
Cb_17_95 bit_17_95 gnd C_bl
Cbb_17_95 bitb_17_95 gnd C_bl
Rb_17_96 bit_17_96 bit_17_97 R_bl
Rbb_17_96 bitb_17_96 bitb_17_97 R_bl
Cb_17_96 bit_17_96 gnd C_bl
Cbb_17_96 bitb_17_96 gnd C_bl
Rb_17_97 bit_17_97 bit_17_98 R_bl
Rbb_17_97 bitb_17_97 bitb_17_98 R_bl
Cb_17_97 bit_17_97 gnd C_bl
Cbb_17_97 bitb_17_97 gnd C_bl
Rb_17_98 bit_17_98 bit_17_99 R_bl
Rbb_17_98 bitb_17_98 bitb_17_99 R_bl
Cb_17_98 bit_17_98 gnd C_bl
Cbb_17_98 bitb_17_98 gnd C_bl
Rb_17_99 bit_17_99 bit_17_100 R_bl
Rbb_17_99 bitb_17_99 bitb_17_100 R_bl
Cb_17_99 bit_17_99 gnd C_bl
Cbb_17_99 bitb_17_99 gnd C_bl
Rb_18_0 bit_18_0 bit_18_1 R_bl
Rbb_18_0 bitb_18_0 bitb_18_1 R_bl
Cb_18_0 bit_18_0 gnd C_bl
Cbb_18_0 bitb_18_0 gnd C_bl
Rb_18_1 bit_18_1 bit_18_2 R_bl
Rbb_18_1 bitb_18_1 bitb_18_2 R_bl
Cb_18_1 bit_18_1 gnd C_bl
Cbb_18_1 bitb_18_1 gnd C_bl
Rb_18_2 bit_18_2 bit_18_3 R_bl
Rbb_18_2 bitb_18_2 bitb_18_3 R_bl
Cb_18_2 bit_18_2 gnd C_bl
Cbb_18_2 bitb_18_2 gnd C_bl
Rb_18_3 bit_18_3 bit_18_4 R_bl
Rbb_18_3 bitb_18_3 bitb_18_4 R_bl
Cb_18_3 bit_18_3 gnd C_bl
Cbb_18_3 bitb_18_3 gnd C_bl
Rb_18_4 bit_18_4 bit_18_5 R_bl
Rbb_18_4 bitb_18_4 bitb_18_5 R_bl
Cb_18_4 bit_18_4 gnd C_bl
Cbb_18_4 bitb_18_4 gnd C_bl
Rb_18_5 bit_18_5 bit_18_6 R_bl
Rbb_18_5 bitb_18_5 bitb_18_6 R_bl
Cb_18_5 bit_18_5 gnd C_bl
Cbb_18_5 bitb_18_5 gnd C_bl
Rb_18_6 bit_18_6 bit_18_7 R_bl
Rbb_18_6 bitb_18_6 bitb_18_7 R_bl
Cb_18_6 bit_18_6 gnd C_bl
Cbb_18_6 bitb_18_6 gnd C_bl
Rb_18_7 bit_18_7 bit_18_8 R_bl
Rbb_18_7 bitb_18_7 bitb_18_8 R_bl
Cb_18_7 bit_18_7 gnd C_bl
Cbb_18_7 bitb_18_7 gnd C_bl
Rb_18_8 bit_18_8 bit_18_9 R_bl
Rbb_18_8 bitb_18_8 bitb_18_9 R_bl
Cb_18_8 bit_18_8 gnd C_bl
Cbb_18_8 bitb_18_8 gnd C_bl
Rb_18_9 bit_18_9 bit_18_10 R_bl
Rbb_18_9 bitb_18_9 bitb_18_10 R_bl
Cb_18_9 bit_18_9 gnd C_bl
Cbb_18_9 bitb_18_9 gnd C_bl
Rb_18_10 bit_18_10 bit_18_11 R_bl
Rbb_18_10 bitb_18_10 bitb_18_11 R_bl
Cb_18_10 bit_18_10 gnd C_bl
Cbb_18_10 bitb_18_10 gnd C_bl
Rb_18_11 bit_18_11 bit_18_12 R_bl
Rbb_18_11 bitb_18_11 bitb_18_12 R_bl
Cb_18_11 bit_18_11 gnd C_bl
Cbb_18_11 bitb_18_11 gnd C_bl
Rb_18_12 bit_18_12 bit_18_13 R_bl
Rbb_18_12 bitb_18_12 bitb_18_13 R_bl
Cb_18_12 bit_18_12 gnd C_bl
Cbb_18_12 bitb_18_12 gnd C_bl
Rb_18_13 bit_18_13 bit_18_14 R_bl
Rbb_18_13 bitb_18_13 bitb_18_14 R_bl
Cb_18_13 bit_18_13 gnd C_bl
Cbb_18_13 bitb_18_13 gnd C_bl
Rb_18_14 bit_18_14 bit_18_15 R_bl
Rbb_18_14 bitb_18_14 bitb_18_15 R_bl
Cb_18_14 bit_18_14 gnd C_bl
Cbb_18_14 bitb_18_14 gnd C_bl
Rb_18_15 bit_18_15 bit_18_16 R_bl
Rbb_18_15 bitb_18_15 bitb_18_16 R_bl
Cb_18_15 bit_18_15 gnd C_bl
Cbb_18_15 bitb_18_15 gnd C_bl
Rb_18_16 bit_18_16 bit_18_17 R_bl
Rbb_18_16 bitb_18_16 bitb_18_17 R_bl
Cb_18_16 bit_18_16 gnd C_bl
Cbb_18_16 bitb_18_16 gnd C_bl
Rb_18_17 bit_18_17 bit_18_18 R_bl
Rbb_18_17 bitb_18_17 bitb_18_18 R_bl
Cb_18_17 bit_18_17 gnd C_bl
Cbb_18_17 bitb_18_17 gnd C_bl
Rb_18_18 bit_18_18 bit_18_19 R_bl
Rbb_18_18 bitb_18_18 bitb_18_19 R_bl
Cb_18_18 bit_18_18 gnd C_bl
Cbb_18_18 bitb_18_18 gnd C_bl
Rb_18_19 bit_18_19 bit_18_20 R_bl
Rbb_18_19 bitb_18_19 bitb_18_20 R_bl
Cb_18_19 bit_18_19 gnd C_bl
Cbb_18_19 bitb_18_19 gnd C_bl
Rb_18_20 bit_18_20 bit_18_21 R_bl
Rbb_18_20 bitb_18_20 bitb_18_21 R_bl
Cb_18_20 bit_18_20 gnd C_bl
Cbb_18_20 bitb_18_20 gnd C_bl
Rb_18_21 bit_18_21 bit_18_22 R_bl
Rbb_18_21 bitb_18_21 bitb_18_22 R_bl
Cb_18_21 bit_18_21 gnd C_bl
Cbb_18_21 bitb_18_21 gnd C_bl
Rb_18_22 bit_18_22 bit_18_23 R_bl
Rbb_18_22 bitb_18_22 bitb_18_23 R_bl
Cb_18_22 bit_18_22 gnd C_bl
Cbb_18_22 bitb_18_22 gnd C_bl
Rb_18_23 bit_18_23 bit_18_24 R_bl
Rbb_18_23 bitb_18_23 bitb_18_24 R_bl
Cb_18_23 bit_18_23 gnd C_bl
Cbb_18_23 bitb_18_23 gnd C_bl
Rb_18_24 bit_18_24 bit_18_25 R_bl
Rbb_18_24 bitb_18_24 bitb_18_25 R_bl
Cb_18_24 bit_18_24 gnd C_bl
Cbb_18_24 bitb_18_24 gnd C_bl
Rb_18_25 bit_18_25 bit_18_26 R_bl
Rbb_18_25 bitb_18_25 bitb_18_26 R_bl
Cb_18_25 bit_18_25 gnd C_bl
Cbb_18_25 bitb_18_25 gnd C_bl
Rb_18_26 bit_18_26 bit_18_27 R_bl
Rbb_18_26 bitb_18_26 bitb_18_27 R_bl
Cb_18_26 bit_18_26 gnd C_bl
Cbb_18_26 bitb_18_26 gnd C_bl
Rb_18_27 bit_18_27 bit_18_28 R_bl
Rbb_18_27 bitb_18_27 bitb_18_28 R_bl
Cb_18_27 bit_18_27 gnd C_bl
Cbb_18_27 bitb_18_27 gnd C_bl
Rb_18_28 bit_18_28 bit_18_29 R_bl
Rbb_18_28 bitb_18_28 bitb_18_29 R_bl
Cb_18_28 bit_18_28 gnd C_bl
Cbb_18_28 bitb_18_28 gnd C_bl
Rb_18_29 bit_18_29 bit_18_30 R_bl
Rbb_18_29 bitb_18_29 bitb_18_30 R_bl
Cb_18_29 bit_18_29 gnd C_bl
Cbb_18_29 bitb_18_29 gnd C_bl
Rb_18_30 bit_18_30 bit_18_31 R_bl
Rbb_18_30 bitb_18_30 bitb_18_31 R_bl
Cb_18_30 bit_18_30 gnd C_bl
Cbb_18_30 bitb_18_30 gnd C_bl
Rb_18_31 bit_18_31 bit_18_32 R_bl
Rbb_18_31 bitb_18_31 bitb_18_32 R_bl
Cb_18_31 bit_18_31 gnd C_bl
Cbb_18_31 bitb_18_31 gnd C_bl
Rb_18_32 bit_18_32 bit_18_33 R_bl
Rbb_18_32 bitb_18_32 bitb_18_33 R_bl
Cb_18_32 bit_18_32 gnd C_bl
Cbb_18_32 bitb_18_32 gnd C_bl
Rb_18_33 bit_18_33 bit_18_34 R_bl
Rbb_18_33 bitb_18_33 bitb_18_34 R_bl
Cb_18_33 bit_18_33 gnd C_bl
Cbb_18_33 bitb_18_33 gnd C_bl
Rb_18_34 bit_18_34 bit_18_35 R_bl
Rbb_18_34 bitb_18_34 bitb_18_35 R_bl
Cb_18_34 bit_18_34 gnd C_bl
Cbb_18_34 bitb_18_34 gnd C_bl
Rb_18_35 bit_18_35 bit_18_36 R_bl
Rbb_18_35 bitb_18_35 bitb_18_36 R_bl
Cb_18_35 bit_18_35 gnd C_bl
Cbb_18_35 bitb_18_35 gnd C_bl
Rb_18_36 bit_18_36 bit_18_37 R_bl
Rbb_18_36 bitb_18_36 bitb_18_37 R_bl
Cb_18_36 bit_18_36 gnd C_bl
Cbb_18_36 bitb_18_36 gnd C_bl
Rb_18_37 bit_18_37 bit_18_38 R_bl
Rbb_18_37 bitb_18_37 bitb_18_38 R_bl
Cb_18_37 bit_18_37 gnd C_bl
Cbb_18_37 bitb_18_37 gnd C_bl
Rb_18_38 bit_18_38 bit_18_39 R_bl
Rbb_18_38 bitb_18_38 bitb_18_39 R_bl
Cb_18_38 bit_18_38 gnd C_bl
Cbb_18_38 bitb_18_38 gnd C_bl
Rb_18_39 bit_18_39 bit_18_40 R_bl
Rbb_18_39 bitb_18_39 bitb_18_40 R_bl
Cb_18_39 bit_18_39 gnd C_bl
Cbb_18_39 bitb_18_39 gnd C_bl
Rb_18_40 bit_18_40 bit_18_41 R_bl
Rbb_18_40 bitb_18_40 bitb_18_41 R_bl
Cb_18_40 bit_18_40 gnd C_bl
Cbb_18_40 bitb_18_40 gnd C_bl
Rb_18_41 bit_18_41 bit_18_42 R_bl
Rbb_18_41 bitb_18_41 bitb_18_42 R_bl
Cb_18_41 bit_18_41 gnd C_bl
Cbb_18_41 bitb_18_41 gnd C_bl
Rb_18_42 bit_18_42 bit_18_43 R_bl
Rbb_18_42 bitb_18_42 bitb_18_43 R_bl
Cb_18_42 bit_18_42 gnd C_bl
Cbb_18_42 bitb_18_42 gnd C_bl
Rb_18_43 bit_18_43 bit_18_44 R_bl
Rbb_18_43 bitb_18_43 bitb_18_44 R_bl
Cb_18_43 bit_18_43 gnd C_bl
Cbb_18_43 bitb_18_43 gnd C_bl
Rb_18_44 bit_18_44 bit_18_45 R_bl
Rbb_18_44 bitb_18_44 bitb_18_45 R_bl
Cb_18_44 bit_18_44 gnd C_bl
Cbb_18_44 bitb_18_44 gnd C_bl
Rb_18_45 bit_18_45 bit_18_46 R_bl
Rbb_18_45 bitb_18_45 bitb_18_46 R_bl
Cb_18_45 bit_18_45 gnd C_bl
Cbb_18_45 bitb_18_45 gnd C_bl
Rb_18_46 bit_18_46 bit_18_47 R_bl
Rbb_18_46 bitb_18_46 bitb_18_47 R_bl
Cb_18_46 bit_18_46 gnd C_bl
Cbb_18_46 bitb_18_46 gnd C_bl
Rb_18_47 bit_18_47 bit_18_48 R_bl
Rbb_18_47 bitb_18_47 bitb_18_48 R_bl
Cb_18_47 bit_18_47 gnd C_bl
Cbb_18_47 bitb_18_47 gnd C_bl
Rb_18_48 bit_18_48 bit_18_49 R_bl
Rbb_18_48 bitb_18_48 bitb_18_49 R_bl
Cb_18_48 bit_18_48 gnd C_bl
Cbb_18_48 bitb_18_48 gnd C_bl
Rb_18_49 bit_18_49 bit_18_50 R_bl
Rbb_18_49 bitb_18_49 bitb_18_50 R_bl
Cb_18_49 bit_18_49 gnd C_bl
Cbb_18_49 bitb_18_49 gnd C_bl
Rb_18_50 bit_18_50 bit_18_51 R_bl
Rbb_18_50 bitb_18_50 bitb_18_51 R_bl
Cb_18_50 bit_18_50 gnd C_bl
Cbb_18_50 bitb_18_50 gnd C_bl
Rb_18_51 bit_18_51 bit_18_52 R_bl
Rbb_18_51 bitb_18_51 bitb_18_52 R_bl
Cb_18_51 bit_18_51 gnd C_bl
Cbb_18_51 bitb_18_51 gnd C_bl
Rb_18_52 bit_18_52 bit_18_53 R_bl
Rbb_18_52 bitb_18_52 bitb_18_53 R_bl
Cb_18_52 bit_18_52 gnd C_bl
Cbb_18_52 bitb_18_52 gnd C_bl
Rb_18_53 bit_18_53 bit_18_54 R_bl
Rbb_18_53 bitb_18_53 bitb_18_54 R_bl
Cb_18_53 bit_18_53 gnd C_bl
Cbb_18_53 bitb_18_53 gnd C_bl
Rb_18_54 bit_18_54 bit_18_55 R_bl
Rbb_18_54 bitb_18_54 bitb_18_55 R_bl
Cb_18_54 bit_18_54 gnd C_bl
Cbb_18_54 bitb_18_54 gnd C_bl
Rb_18_55 bit_18_55 bit_18_56 R_bl
Rbb_18_55 bitb_18_55 bitb_18_56 R_bl
Cb_18_55 bit_18_55 gnd C_bl
Cbb_18_55 bitb_18_55 gnd C_bl
Rb_18_56 bit_18_56 bit_18_57 R_bl
Rbb_18_56 bitb_18_56 bitb_18_57 R_bl
Cb_18_56 bit_18_56 gnd C_bl
Cbb_18_56 bitb_18_56 gnd C_bl
Rb_18_57 bit_18_57 bit_18_58 R_bl
Rbb_18_57 bitb_18_57 bitb_18_58 R_bl
Cb_18_57 bit_18_57 gnd C_bl
Cbb_18_57 bitb_18_57 gnd C_bl
Rb_18_58 bit_18_58 bit_18_59 R_bl
Rbb_18_58 bitb_18_58 bitb_18_59 R_bl
Cb_18_58 bit_18_58 gnd C_bl
Cbb_18_58 bitb_18_58 gnd C_bl
Rb_18_59 bit_18_59 bit_18_60 R_bl
Rbb_18_59 bitb_18_59 bitb_18_60 R_bl
Cb_18_59 bit_18_59 gnd C_bl
Cbb_18_59 bitb_18_59 gnd C_bl
Rb_18_60 bit_18_60 bit_18_61 R_bl
Rbb_18_60 bitb_18_60 bitb_18_61 R_bl
Cb_18_60 bit_18_60 gnd C_bl
Cbb_18_60 bitb_18_60 gnd C_bl
Rb_18_61 bit_18_61 bit_18_62 R_bl
Rbb_18_61 bitb_18_61 bitb_18_62 R_bl
Cb_18_61 bit_18_61 gnd C_bl
Cbb_18_61 bitb_18_61 gnd C_bl
Rb_18_62 bit_18_62 bit_18_63 R_bl
Rbb_18_62 bitb_18_62 bitb_18_63 R_bl
Cb_18_62 bit_18_62 gnd C_bl
Cbb_18_62 bitb_18_62 gnd C_bl
Rb_18_63 bit_18_63 bit_18_64 R_bl
Rbb_18_63 bitb_18_63 bitb_18_64 R_bl
Cb_18_63 bit_18_63 gnd C_bl
Cbb_18_63 bitb_18_63 gnd C_bl
Rb_18_64 bit_18_64 bit_18_65 R_bl
Rbb_18_64 bitb_18_64 bitb_18_65 R_bl
Cb_18_64 bit_18_64 gnd C_bl
Cbb_18_64 bitb_18_64 gnd C_bl
Rb_18_65 bit_18_65 bit_18_66 R_bl
Rbb_18_65 bitb_18_65 bitb_18_66 R_bl
Cb_18_65 bit_18_65 gnd C_bl
Cbb_18_65 bitb_18_65 gnd C_bl
Rb_18_66 bit_18_66 bit_18_67 R_bl
Rbb_18_66 bitb_18_66 bitb_18_67 R_bl
Cb_18_66 bit_18_66 gnd C_bl
Cbb_18_66 bitb_18_66 gnd C_bl
Rb_18_67 bit_18_67 bit_18_68 R_bl
Rbb_18_67 bitb_18_67 bitb_18_68 R_bl
Cb_18_67 bit_18_67 gnd C_bl
Cbb_18_67 bitb_18_67 gnd C_bl
Rb_18_68 bit_18_68 bit_18_69 R_bl
Rbb_18_68 bitb_18_68 bitb_18_69 R_bl
Cb_18_68 bit_18_68 gnd C_bl
Cbb_18_68 bitb_18_68 gnd C_bl
Rb_18_69 bit_18_69 bit_18_70 R_bl
Rbb_18_69 bitb_18_69 bitb_18_70 R_bl
Cb_18_69 bit_18_69 gnd C_bl
Cbb_18_69 bitb_18_69 gnd C_bl
Rb_18_70 bit_18_70 bit_18_71 R_bl
Rbb_18_70 bitb_18_70 bitb_18_71 R_bl
Cb_18_70 bit_18_70 gnd C_bl
Cbb_18_70 bitb_18_70 gnd C_bl
Rb_18_71 bit_18_71 bit_18_72 R_bl
Rbb_18_71 bitb_18_71 bitb_18_72 R_bl
Cb_18_71 bit_18_71 gnd C_bl
Cbb_18_71 bitb_18_71 gnd C_bl
Rb_18_72 bit_18_72 bit_18_73 R_bl
Rbb_18_72 bitb_18_72 bitb_18_73 R_bl
Cb_18_72 bit_18_72 gnd C_bl
Cbb_18_72 bitb_18_72 gnd C_bl
Rb_18_73 bit_18_73 bit_18_74 R_bl
Rbb_18_73 bitb_18_73 bitb_18_74 R_bl
Cb_18_73 bit_18_73 gnd C_bl
Cbb_18_73 bitb_18_73 gnd C_bl
Rb_18_74 bit_18_74 bit_18_75 R_bl
Rbb_18_74 bitb_18_74 bitb_18_75 R_bl
Cb_18_74 bit_18_74 gnd C_bl
Cbb_18_74 bitb_18_74 gnd C_bl
Rb_18_75 bit_18_75 bit_18_76 R_bl
Rbb_18_75 bitb_18_75 bitb_18_76 R_bl
Cb_18_75 bit_18_75 gnd C_bl
Cbb_18_75 bitb_18_75 gnd C_bl
Rb_18_76 bit_18_76 bit_18_77 R_bl
Rbb_18_76 bitb_18_76 bitb_18_77 R_bl
Cb_18_76 bit_18_76 gnd C_bl
Cbb_18_76 bitb_18_76 gnd C_bl
Rb_18_77 bit_18_77 bit_18_78 R_bl
Rbb_18_77 bitb_18_77 bitb_18_78 R_bl
Cb_18_77 bit_18_77 gnd C_bl
Cbb_18_77 bitb_18_77 gnd C_bl
Rb_18_78 bit_18_78 bit_18_79 R_bl
Rbb_18_78 bitb_18_78 bitb_18_79 R_bl
Cb_18_78 bit_18_78 gnd C_bl
Cbb_18_78 bitb_18_78 gnd C_bl
Rb_18_79 bit_18_79 bit_18_80 R_bl
Rbb_18_79 bitb_18_79 bitb_18_80 R_bl
Cb_18_79 bit_18_79 gnd C_bl
Cbb_18_79 bitb_18_79 gnd C_bl
Rb_18_80 bit_18_80 bit_18_81 R_bl
Rbb_18_80 bitb_18_80 bitb_18_81 R_bl
Cb_18_80 bit_18_80 gnd C_bl
Cbb_18_80 bitb_18_80 gnd C_bl
Rb_18_81 bit_18_81 bit_18_82 R_bl
Rbb_18_81 bitb_18_81 bitb_18_82 R_bl
Cb_18_81 bit_18_81 gnd C_bl
Cbb_18_81 bitb_18_81 gnd C_bl
Rb_18_82 bit_18_82 bit_18_83 R_bl
Rbb_18_82 bitb_18_82 bitb_18_83 R_bl
Cb_18_82 bit_18_82 gnd C_bl
Cbb_18_82 bitb_18_82 gnd C_bl
Rb_18_83 bit_18_83 bit_18_84 R_bl
Rbb_18_83 bitb_18_83 bitb_18_84 R_bl
Cb_18_83 bit_18_83 gnd C_bl
Cbb_18_83 bitb_18_83 gnd C_bl
Rb_18_84 bit_18_84 bit_18_85 R_bl
Rbb_18_84 bitb_18_84 bitb_18_85 R_bl
Cb_18_84 bit_18_84 gnd C_bl
Cbb_18_84 bitb_18_84 gnd C_bl
Rb_18_85 bit_18_85 bit_18_86 R_bl
Rbb_18_85 bitb_18_85 bitb_18_86 R_bl
Cb_18_85 bit_18_85 gnd C_bl
Cbb_18_85 bitb_18_85 gnd C_bl
Rb_18_86 bit_18_86 bit_18_87 R_bl
Rbb_18_86 bitb_18_86 bitb_18_87 R_bl
Cb_18_86 bit_18_86 gnd C_bl
Cbb_18_86 bitb_18_86 gnd C_bl
Rb_18_87 bit_18_87 bit_18_88 R_bl
Rbb_18_87 bitb_18_87 bitb_18_88 R_bl
Cb_18_87 bit_18_87 gnd C_bl
Cbb_18_87 bitb_18_87 gnd C_bl
Rb_18_88 bit_18_88 bit_18_89 R_bl
Rbb_18_88 bitb_18_88 bitb_18_89 R_bl
Cb_18_88 bit_18_88 gnd C_bl
Cbb_18_88 bitb_18_88 gnd C_bl
Rb_18_89 bit_18_89 bit_18_90 R_bl
Rbb_18_89 bitb_18_89 bitb_18_90 R_bl
Cb_18_89 bit_18_89 gnd C_bl
Cbb_18_89 bitb_18_89 gnd C_bl
Rb_18_90 bit_18_90 bit_18_91 R_bl
Rbb_18_90 bitb_18_90 bitb_18_91 R_bl
Cb_18_90 bit_18_90 gnd C_bl
Cbb_18_90 bitb_18_90 gnd C_bl
Rb_18_91 bit_18_91 bit_18_92 R_bl
Rbb_18_91 bitb_18_91 bitb_18_92 R_bl
Cb_18_91 bit_18_91 gnd C_bl
Cbb_18_91 bitb_18_91 gnd C_bl
Rb_18_92 bit_18_92 bit_18_93 R_bl
Rbb_18_92 bitb_18_92 bitb_18_93 R_bl
Cb_18_92 bit_18_92 gnd C_bl
Cbb_18_92 bitb_18_92 gnd C_bl
Rb_18_93 bit_18_93 bit_18_94 R_bl
Rbb_18_93 bitb_18_93 bitb_18_94 R_bl
Cb_18_93 bit_18_93 gnd C_bl
Cbb_18_93 bitb_18_93 gnd C_bl
Rb_18_94 bit_18_94 bit_18_95 R_bl
Rbb_18_94 bitb_18_94 bitb_18_95 R_bl
Cb_18_94 bit_18_94 gnd C_bl
Cbb_18_94 bitb_18_94 gnd C_bl
Rb_18_95 bit_18_95 bit_18_96 R_bl
Rbb_18_95 bitb_18_95 bitb_18_96 R_bl
Cb_18_95 bit_18_95 gnd C_bl
Cbb_18_95 bitb_18_95 gnd C_bl
Rb_18_96 bit_18_96 bit_18_97 R_bl
Rbb_18_96 bitb_18_96 bitb_18_97 R_bl
Cb_18_96 bit_18_96 gnd C_bl
Cbb_18_96 bitb_18_96 gnd C_bl
Rb_18_97 bit_18_97 bit_18_98 R_bl
Rbb_18_97 bitb_18_97 bitb_18_98 R_bl
Cb_18_97 bit_18_97 gnd C_bl
Cbb_18_97 bitb_18_97 gnd C_bl
Rb_18_98 bit_18_98 bit_18_99 R_bl
Rbb_18_98 bitb_18_98 bitb_18_99 R_bl
Cb_18_98 bit_18_98 gnd C_bl
Cbb_18_98 bitb_18_98 gnd C_bl
Rb_18_99 bit_18_99 bit_18_100 R_bl
Rbb_18_99 bitb_18_99 bitb_18_100 R_bl
Cb_18_99 bit_18_99 gnd C_bl
Cbb_18_99 bitb_18_99 gnd C_bl
Rb_19_0 bit_19_0 bit_19_1 R_bl
Rbb_19_0 bitb_19_0 bitb_19_1 R_bl
Cb_19_0 bit_19_0 gnd C_bl
Cbb_19_0 bitb_19_0 gnd C_bl
Rb_19_1 bit_19_1 bit_19_2 R_bl
Rbb_19_1 bitb_19_1 bitb_19_2 R_bl
Cb_19_1 bit_19_1 gnd C_bl
Cbb_19_1 bitb_19_1 gnd C_bl
Rb_19_2 bit_19_2 bit_19_3 R_bl
Rbb_19_2 bitb_19_2 bitb_19_3 R_bl
Cb_19_2 bit_19_2 gnd C_bl
Cbb_19_2 bitb_19_2 gnd C_bl
Rb_19_3 bit_19_3 bit_19_4 R_bl
Rbb_19_3 bitb_19_3 bitb_19_4 R_bl
Cb_19_3 bit_19_3 gnd C_bl
Cbb_19_3 bitb_19_3 gnd C_bl
Rb_19_4 bit_19_4 bit_19_5 R_bl
Rbb_19_4 bitb_19_4 bitb_19_5 R_bl
Cb_19_4 bit_19_4 gnd C_bl
Cbb_19_4 bitb_19_4 gnd C_bl
Rb_19_5 bit_19_5 bit_19_6 R_bl
Rbb_19_5 bitb_19_5 bitb_19_6 R_bl
Cb_19_5 bit_19_5 gnd C_bl
Cbb_19_5 bitb_19_5 gnd C_bl
Rb_19_6 bit_19_6 bit_19_7 R_bl
Rbb_19_6 bitb_19_6 bitb_19_7 R_bl
Cb_19_6 bit_19_6 gnd C_bl
Cbb_19_6 bitb_19_6 gnd C_bl
Rb_19_7 bit_19_7 bit_19_8 R_bl
Rbb_19_7 bitb_19_7 bitb_19_8 R_bl
Cb_19_7 bit_19_7 gnd C_bl
Cbb_19_7 bitb_19_7 gnd C_bl
Rb_19_8 bit_19_8 bit_19_9 R_bl
Rbb_19_8 bitb_19_8 bitb_19_9 R_bl
Cb_19_8 bit_19_8 gnd C_bl
Cbb_19_8 bitb_19_8 gnd C_bl
Rb_19_9 bit_19_9 bit_19_10 R_bl
Rbb_19_9 bitb_19_9 bitb_19_10 R_bl
Cb_19_9 bit_19_9 gnd C_bl
Cbb_19_9 bitb_19_9 gnd C_bl
Rb_19_10 bit_19_10 bit_19_11 R_bl
Rbb_19_10 bitb_19_10 bitb_19_11 R_bl
Cb_19_10 bit_19_10 gnd C_bl
Cbb_19_10 bitb_19_10 gnd C_bl
Rb_19_11 bit_19_11 bit_19_12 R_bl
Rbb_19_11 bitb_19_11 bitb_19_12 R_bl
Cb_19_11 bit_19_11 gnd C_bl
Cbb_19_11 bitb_19_11 gnd C_bl
Rb_19_12 bit_19_12 bit_19_13 R_bl
Rbb_19_12 bitb_19_12 bitb_19_13 R_bl
Cb_19_12 bit_19_12 gnd C_bl
Cbb_19_12 bitb_19_12 gnd C_bl
Rb_19_13 bit_19_13 bit_19_14 R_bl
Rbb_19_13 bitb_19_13 bitb_19_14 R_bl
Cb_19_13 bit_19_13 gnd C_bl
Cbb_19_13 bitb_19_13 gnd C_bl
Rb_19_14 bit_19_14 bit_19_15 R_bl
Rbb_19_14 bitb_19_14 bitb_19_15 R_bl
Cb_19_14 bit_19_14 gnd C_bl
Cbb_19_14 bitb_19_14 gnd C_bl
Rb_19_15 bit_19_15 bit_19_16 R_bl
Rbb_19_15 bitb_19_15 bitb_19_16 R_bl
Cb_19_15 bit_19_15 gnd C_bl
Cbb_19_15 bitb_19_15 gnd C_bl
Rb_19_16 bit_19_16 bit_19_17 R_bl
Rbb_19_16 bitb_19_16 bitb_19_17 R_bl
Cb_19_16 bit_19_16 gnd C_bl
Cbb_19_16 bitb_19_16 gnd C_bl
Rb_19_17 bit_19_17 bit_19_18 R_bl
Rbb_19_17 bitb_19_17 bitb_19_18 R_bl
Cb_19_17 bit_19_17 gnd C_bl
Cbb_19_17 bitb_19_17 gnd C_bl
Rb_19_18 bit_19_18 bit_19_19 R_bl
Rbb_19_18 bitb_19_18 bitb_19_19 R_bl
Cb_19_18 bit_19_18 gnd C_bl
Cbb_19_18 bitb_19_18 gnd C_bl
Rb_19_19 bit_19_19 bit_19_20 R_bl
Rbb_19_19 bitb_19_19 bitb_19_20 R_bl
Cb_19_19 bit_19_19 gnd C_bl
Cbb_19_19 bitb_19_19 gnd C_bl
Rb_19_20 bit_19_20 bit_19_21 R_bl
Rbb_19_20 bitb_19_20 bitb_19_21 R_bl
Cb_19_20 bit_19_20 gnd C_bl
Cbb_19_20 bitb_19_20 gnd C_bl
Rb_19_21 bit_19_21 bit_19_22 R_bl
Rbb_19_21 bitb_19_21 bitb_19_22 R_bl
Cb_19_21 bit_19_21 gnd C_bl
Cbb_19_21 bitb_19_21 gnd C_bl
Rb_19_22 bit_19_22 bit_19_23 R_bl
Rbb_19_22 bitb_19_22 bitb_19_23 R_bl
Cb_19_22 bit_19_22 gnd C_bl
Cbb_19_22 bitb_19_22 gnd C_bl
Rb_19_23 bit_19_23 bit_19_24 R_bl
Rbb_19_23 bitb_19_23 bitb_19_24 R_bl
Cb_19_23 bit_19_23 gnd C_bl
Cbb_19_23 bitb_19_23 gnd C_bl
Rb_19_24 bit_19_24 bit_19_25 R_bl
Rbb_19_24 bitb_19_24 bitb_19_25 R_bl
Cb_19_24 bit_19_24 gnd C_bl
Cbb_19_24 bitb_19_24 gnd C_bl
Rb_19_25 bit_19_25 bit_19_26 R_bl
Rbb_19_25 bitb_19_25 bitb_19_26 R_bl
Cb_19_25 bit_19_25 gnd C_bl
Cbb_19_25 bitb_19_25 gnd C_bl
Rb_19_26 bit_19_26 bit_19_27 R_bl
Rbb_19_26 bitb_19_26 bitb_19_27 R_bl
Cb_19_26 bit_19_26 gnd C_bl
Cbb_19_26 bitb_19_26 gnd C_bl
Rb_19_27 bit_19_27 bit_19_28 R_bl
Rbb_19_27 bitb_19_27 bitb_19_28 R_bl
Cb_19_27 bit_19_27 gnd C_bl
Cbb_19_27 bitb_19_27 gnd C_bl
Rb_19_28 bit_19_28 bit_19_29 R_bl
Rbb_19_28 bitb_19_28 bitb_19_29 R_bl
Cb_19_28 bit_19_28 gnd C_bl
Cbb_19_28 bitb_19_28 gnd C_bl
Rb_19_29 bit_19_29 bit_19_30 R_bl
Rbb_19_29 bitb_19_29 bitb_19_30 R_bl
Cb_19_29 bit_19_29 gnd C_bl
Cbb_19_29 bitb_19_29 gnd C_bl
Rb_19_30 bit_19_30 bit_19_31 R_bl
Rbb_19_30 bitb_19_30 bitb_19_31 R_bl
Cb_19_30 bit_19_30 gnd C_bl
Cbb_19_30 bitb_19_30 gnd C_bl
Rb_19_31 bit_19_31 bit_19_32 R_bl
Rbb_19_31 bitb_19_31 bitb_19_32 R_bl
Cb_19_31 bit_19_31 gnd C_bl
Cbb_19_31 bitb_19_31 gnd C_bl
Rb_19_32 bit_19_32 bit_19_33 R_bl
Rbb_19_32 bitb_19_32 bitb_19_33 R_bl
Cb_19_32 bit_19_32 gnd C_bl
Cbb_19_32 bitb_19_32 gnd C_bl
Rb_19_33 bit_19_33 bit_19_34 R_bl
Rbb_19_33 bitb_19_33 bitb_19_34 R_bl
Cb_19_33 bit_19_33 gnd C_bl
Cbb_19_33 bitb_19_33 gnd C_bl
Rb_19_34 bit_19_34 bit_19_35 R_bl
Rbb_19_34 bitb_19_34 bitb_19_35 R_bl
Cb_19_34 bit_19_34 gnd C_bl
Cbb_19_34 bitb_19_34 gnd C_bl
Rb_19_35 bit_19_35 bit_19_36 R_bl
Rbb_19_35 bitb_19_35 bitb_19_36 R_bl
Cb_19_35 bit_19_35 gnd C_bl
Cbb_19_35 bitb_19_35 gnd C_bl
Rb_19_36 bit_19_36 bit_19_37 R_bl
Rbb_19_36 bitb_19_36 bitb_19_37 R_bl
Cb_19_36 bit_19_36 gnd C_bl
Cbb_19_36 bitb_19_36 gnd C_bl
Rb_19_37 bit_19_37 bit_19_38 R_bl
Rbb_19_37 bitb_19_37 bitb_19_38 R_bl
Cb_19_37 bit_19_37 gnd C_bl
Cbb_19_37 bitb_19_37 gnd C_bl
Rb_19_38 bit_19_38 bit_19_39 R_bl
Rbb_19_38 bitb_19_38 bitb_19_39 R_bl
Cb_19_38 bit_19_38 gnd C_bl
Cbb_19_38 bitb_19_38 gnd C_bl
Rb_19_39 bit_19_39 bit_19_40 R_bl
Rbb_19_39 bitb_19_39 bitb_19_40 R_bl
Cb_19_39 bit_19_39 gnd C_bl
Cbb_19_39 bitb_19_39 gnd C_bl
Rb_19_40 bit_19_40 bit_19_41 R_bl
Rbb_19_40 bitb_19_40 bitb_19_41 R_bl
Cb_19_40 bit_19_40 gnd C_bl
Cbb_19_40 bitb_19_40 gnd C_bl
Rb_19_41 bit_19_41 bit_19_42 R_bl
Rbb_19_41 bitb_19_41 bitb_19_42 R_bl
Cb_19_41 bit_19_41 gnd C_bl
Cbb_19_41 bitb_19_41 gnd C_bl
Rb_19_42 bit_19_42 bit_19_43 R_bl
Rbb_19_42 bitb_19_42 bitb_19_43 R_bl
Cb_19_42 bit_19_42 gnd C_bl
Cbb_19_42 bitb_19_42 gnd C_bl
Rb_19_43 bit_19_43 bit_19_44 R_bl
Rbb_19_43 bitb_19_43 bitb_19_44 R_bl
Cb_19_43 bit_19_43 gnd C_bl
Cbb_19_43 bitb_19_43 gnd C_bl
Rb_19_44 bit_19_44 bit_19_45 R_bl
Rbb_19_44 bitb_19_44 bitb_19_45 R_bl
Cb_19_44 bit_19_44 gnd C_bl
Cbb_19_44 bitb_19_44 gnd C_bl
Rb_19_45 bit_19_45 bit_19_46 R_bl
Rbb_19_45 bitb_19_45 bitb_19_46 R_bl
Cb_19_45 bit_19_45 gnd C_bl
Cbb_19_45 bitb_19_45 gnd C_bl
Rb_19_46 bit_19_46 bit_19_47 R_bl
Rbb_19_46 bitb_19_46 bitb_19_47 R_bl
Cb_19_46 bit_19_46 gnd C_bl
Cbb_19_46 bitb_19_46 gnd C_bl
Rb_19_47 bit_19_47 bit_19_48 R_bl
Rbb_19_47 bitb_19_47 bitb_19_48 R_bl
Cb_19_47 bit_19_47 gnd C_bl
Cbb_19_47 bitb_19_47 gnd C_bl
Rb_19_48 bit_19_48 bit_19_49 R_bl
Rbb_19_48 bitb_19_48 bitb_19_49 R_bl
Cb_19_48 bit_19_48 gnd C_bl
Cbb_19_48 bitb_19_48 gnd C_bl
Rb_19_49 bit_19_49 bit_19_50 R_bl
Rbb_19_49 bitb_19_49 bitb_19_50 R_bl
Cb_19_49 bit_19_49 gnd C_bl
Cbb_19_49 bitb_19_49 gnd C_bl
Rb_19_50 bit_19_50 bit_19_51 R_bl
Rbb_19_50 bitb_19_50 bitb_19_51 R_bl
Cb_19_50 bit_19_50 gnd C_bl
Cbb_19_50 bitb_19_50 gnd C_bl
Rb_19_51 bit_19_51 bit_19_52 R_bl
Rbb_19_51 bitb_19_51 bitb_19_52 R_bl
Cb_19_51 bit_19_51 gnd C_bl
Cbb_19_51 bitb_19_51 gnd C_bl
Rb_19_52 bit_19_52 bit_19_53 R_bl
Rbb_19_52 bitb_19_52 bitb_19_53 R_bl
Cb_19_52 bit_19_52 gnd C_bl
Cbb_19_52 bitb_19_52 gnd C_bl
Rb_19_53 bit_19_53 bit_19_54 R_bl
Rbb_19_53 bitb_19_53 bitb_19_54 R_bl
Cb_19_53 bit_19_53 gnd C_bl
Cbb_19_53 bitb_19_53 gnd C_bl
Rb_19_54 bit_19_54 bit_19_55 R_bl
Rbb_19_54 bitb_19_54 bitb_19_55 R_bl
Cb_19_54 bit_19_54 gnd C_bl
Cbb_19_54 bitb_19_54 gnd C_bl
Rb_19_55 bit_19_55 bit_19_56 R_bl
Rbb_19_55 bitb_19_55 bitb_19_56 R_bl
Cb_19_55 bit_19_55 gnd C_bl
Cbb_19_55 bitb_19_55 gnd C_bl
Rb_19_56 bit_19_56 bit_19_57 R_bl
Rbb_19_56 bitb_19_56 bitb_19_57 R_bl
Cb_19_56 bit_19_56 gnd C_bl
Cbb_19_56 bitb_19_56 gnd C_bl
Rb_19_57 bit_19_57 bit_19_58 R_bl
Rbb_19_57 bitb_19_57 bitb_19_58 R_bl
Cb_19_57 bit_19_57 gnd C_bl
Cbb_19_57 bitb_19_57 gnd C_bl
Rb_19_58 bit_19_58 bit_19_59 R_bl
Rbb_19_58 bitb_19_58 bitb_19_59 R_bl
Cb_19_58 bit_19_58 gnd C_bl
Cbb_19_58 bitb_19_58 gnd C_bl
Rb_19_59 bit_19_59 bit_19_60 R_bl
Rbb_19_59 bitb_19_59 bitb_19_60 R_bl
Cb_19_59 bit_19_59 gnd C_bl
Cbb_19_59 bitb_19_59 gnd C_bl
Rb_19_60 bit_19_60 bit_19_61 R_bl
Rbb_19_60 bitb_19_60 bitb_19_61 R_bl
Cb_19_60 bit_19_60 gnd C_bl
Cbb_19_60 bitb_19_60 gnd C_bl
Rb_19_61 bit_19_61 bit_19_62 R_bl
Rbb_19_61 bitb_19_61 bitb_19_62 R_bl
Cb_19_61 bit_19_61 gnd C_bl
Cbb_19_61 bitb_19_61 gnd C_bl
Rb_19_62 bit_19_62 bit_19_63 R_bl
Rbb_19_62 bitb_19_62 bitb_19_63 R_bl
Cb_19_62 bit_19_62 gnd C_bl
Cbb_19_62 bitb_19_62 gnd C_bl
Rb_19_63 bit_19_63 bit_19_64 R_bl
Rbb_19_63 bitb_19_63 bitb_19_64 R_bl
Cb_19_63 bit_19_63 gnd C_bl
Cbb_19_63 bitb_19_63 gnd C_bl
Rb_19_64 bit_19_64 bit_19_65 R_bl
Rbb_19_64 bitb_19_64 bitb_19_65 R_bl
Cb_19_64 bit_19_64 gnd C_bl
Cbb_19_64 bitb_19_64 gnd C_bl
Rb_19_65 bit_19_65 bit_19_66 R_bl
Rbb_19_65 bitb_19_65 bitb_19_66 R_bl
Cb_19_65 bit_19_65 gnd C_bl
Cbb_19_65 bitb_19_65 gnd C_bl
Rb_19_66 bit_19_66 bit_19_67 R_bl
Rbb_19_66 bitb_19_66 bitb_19_67 R_bl
Cb_19_66 bit_19_66 gnd C_bl
Cbb_19_66 bitb_19_66 gnd C_bl
Rb_19_67 bit_19_67 bit_19_68 R_bl
Rbb_19_67 bitb_19_67 bitb_19_68 R_bl
Cb_19_67 bit_19_67 gnd C_bl
Cbb_19_67 bitb_19_67 gnd C_bl
Rb_19_68 bit_19_68 bit_19_69 R_bl
Rbb_19_68 bitb_19_68 bitb_19_69 R_bl
Cb_19_68 bit_19_68 gnd C_bl
Cbb_19_68 bitb_19_68 gnd C_bl
Rb_19_69 bit_19_69 bit_19_70 R_bl
Rbb_19_69 bitb_19_69 bitb_19_70 R_bl
Cb_19_69 bit_19_69 gnd C_bl
Cbb_19_69 bitb_19_69 gnd C_bl
Rb_19_70 bit_19_70 bit_19_71 R_bl
Rbb_19_70 bitb_19_70 bitb_19_71 R_bl
Cb_19_70 bit_19_70 gnd C_bl
Cbb_19_70 bitb_19_70 gnd C_bl
Rb_19_71 bit_19_71 bit_19_72 R_bl
Rbb_19_71 bitb_19_71 bitb_19_72 R_bl
Cb_19_71 bit_19_71 gnd C_bl
Cbb_19_71 bitb_19_71 gnd C_bl
Rb_19_72 bit_19_72 bit_19_73 R_bl
Rbb_19_72 bitb_19_72 bitb_19_73 R_bl
Cb_19_72 bit_19_72 gnd C_bl
Cbb_19_72 bitb_19_72 gnd C_bl
Rb_19_73 bit_19_73 bit_19_74 R_bl
Rbb_19_73 bitb_19_73 bitb_19_74 R_bl
Cb_19_73 bit_19_73 gnd C_bl
Cbb_19_73 bitb_19_73 gnd C_bl
Rb_19_74 bit_19_74 bit_19_75 R_bl
Rbb_19_74 bitb_19_74 bitb_19_75 R_bl
Cb_19_74 bit_19_74 gnd C_bl
Cbb_19_74 bitb_19_74 gnd C_bl
Rb_19_75 bit_19_75 bit_19_76 R_bl
Rbb_19_75 bitb_19_75 bitb_19_76 R_bl
Cb_19_75 bit_19_75 gnd C_bl
Cbb_19_75 bitb_19_75 gnd C_bl
Rb_19_76 bit_19_76 bit_19_77 R_bl
Rbb_19_76 bitb_19_76 bitb_19_77 R_bl
Cb_19_76 bit_19_76 gnd C_bl
Cbb_19_76 bitb_19_76 gnd C_bl
Rb_19_77 bit_19_77 bit_19_78 R_bl
Rbb_19_77 bitb_19_77 bitb_19_78 R_bl
Cb_19_77 bit_19_77 gnd C_bl
Cbb_19_77 bitb_19_77 gnd C_bl
Rb_19_78 bit_19_78 bit_19_79 R_bl
Rbb_19_78 bitb_19_78 bitb_19_79 R_bl
Cb_19_78 bit_19_78 gnd C_bl
Cbb_19_78 bitb_19_78 gnd C_bl
Rb_19_79 bit_19_79 bit_19_80 R_bl
Rbb_19_79 bitb_19_79 bitb_19_80 R_bl
Cb_19_79 bit_19_79 gnd C_bl
Cbb_19_79 bitb_19_79 gnd C_bl
Rb_19_80 bit_19_80 bit_19_81 R_bl
Rbb_19_80 bitb_19_80 bitb_19_81 R_bl
Cb_19_80 bit_19_80 gnd C_bl
Cbb_19_80 bitb_19_80 gnd C_bl
Rb_19_81 bit_19_81 bit_19_82 R_bl
Rbb_19_81 bitb_19_81 bitb_19_82 R_bl
Cb_19_81 bit_19_81 gnd C_bl
Cbb_19_81 bitb_19_81 gnd C_bl
Rb_19_82 bit_19_82 bit_19_83 R_bl
Rbb_19_82 bitb_19_82 bitb_19_83 R_bl
Cb_19_82 bit_19_82 gnd C_bl
Cbb_19_82 bitb_19_82 gnd C_bl
Rb_19_83 bit_19_83 bit_19_84 R_bl
Rbb_19_83 bitb_19_83 bitb_19_84 R_bl
Cb_19_83 bit_19_83 gnd C_bl
Cbb_19_83 bitb_19_83 gnd C_bl
Rb_19_84 bit_19_84 bit_19_85 R_bl
Rbb_19_84 bitb_19_84 bitb_19_85 R_bl
Cb_19_84 bit_19_84 gnd C_bl
Cbb_19_84 bitb_19_84 gnd C_bl
Rb_19_85 bit_19_85 bit_19_86 R_bl
Rbb_19_85 bitb_19_85 bitb_19_86 R_bl
Cb_19_85 bit_19_85 gnd C_bl
Cbb_19_85 bitb_19_85 gnd C_bl
Rb_19_86 bit_19_86 bit_19_87 R_bl
Rbb_19_86 bitb_19_86 bitb_19_87 R_bl
Cb_19_86 bit_19_86 gnd C_bl
Cbb_19_86 bitb_19_86 gnd C_bl
Rb_19_87 bit_19_87 bit_19_88 R_bl
Rbb_19_87 bitb_19_87 bitb_19_88 R_bl
Cb_19_87 bit_19_87 gnd C_bl
Cbb_19_87 bitb_19_87 gnd C_bl
Rb_19_88 bit_19_88 bit_19_89 R_bl
Rbb_19_88 bitb_19_88 bitb_19_89 R_bl
Cb_19_88 bit_19_88 gnd C_bl
Cbb_19_88 bitb_19_88 gnd C_bl
Rb_19_89 bit_19_89 bit_19_90 R_bl
Rbb_19_89 bitb_19_89 bitb_19_90 R_bl
Cb_19_89 bit_19_89 gnd C_bl
Cbb_19_89 bitb_19_89 gnd C_bl
Rb_19_90 bit_19_90 bit_19_91 R_bl
Rbb_19_90 bitb_19_90 bitb_19_91 R_bl
Cb_19_90 bit_19_90 gnd C_bl
Cbb_19_90 bitb_19_90 gnd C_bl
Rb_19_91 bit_19_91 bit_19_92 R_bl
Rbb_19_91 bitb_19_91 bitb_19_92 R_bl
Cb_19_91 bit_19_91 gnd C_bl
Cbb_19_91 bitb_19_91 gnd C_bl
Rb_19_92 bit_19_92 bit_19_93 R_bl
Rbb_19_92 bitb_19_92 bitb_19_93 R_bl
Cb_19_92 bit_19_92 gnd C_bl
Cbb_19_92 bitb_19_92 gnd C_bl
Rb_19_93 bit_19_93 bit_19_94 R_bl
Rbb_19_93 bitb_19_93 bitb_19_94 R_bl
Cb_19_93 bit_19_93 gnd C_bl
Cbb_19_93 bitb_19_93 gnd C_bl
Rb_19_94 bit_19_94 bit_19_95 R_bl
Rbb_19_94 bitb_19_94 bitb_19_95 R_bl
Cb_19_94 bit_19_94 gnd C_bl
Cbb_19_94 bitb_19_94 gnd C_bl
Rb_19_95 bit_19_95 bit_19_96 R_bl
Rbb_19_95 bitb_19_95 bitb_19_96 R_bl
Cb_19_95 bit_19_95 gnd C_bl
Cbb_19_95 bitb_19_95 gnd C_bl
Rb_19_96 bit_19_96 bit_19_97 R_bl
Rbb_19_96 bitb_19_96 bitb_19_97 R_bl
Cb_19_96 bit_19_96 gnd C_bl
Cbb_19_96 bitb_19_96 gnd C_bl
Rb_19_97 bit_19_97 bit_19_98 R_bl
Rbb_19_97 bitb_19_97 bitb_19_98 R_bl
Cb_19_97 bit_19_97 gnd C_bl
Cbb_19_97 bitb_19_97 gnd C_bl
Rb_19_98 bit_19_98 bit_19_99 R_bl
Rbb_19_98 bitb_19_98 bitb_19_99 R_bl
Cb_19_98 bit_19_98 gnd C_bl
Cbb_19_98 bitb_19_98 gnd C_bl
Rb_19_99 bit_19_99 bit_19_100 R_bl
Rbb_19_99 bitb_19_99 bitb_19_100 R_bl
Cb_19_99 bit_19_99 gnd C_bl
Cbb_19_99 bitb_19_99 gnd C_bl
Rb_20_0 bit_20_0 bit_20_1 R_bl
Rbb_20_0 bitb_20_0 bitb_20_1 R_bl
Cb_20_0 bit_20_0 gnd C_bl
Cbb_20_0 bitb_20_0 gnd C_bl
Rb_20_1 bit_20_1 bit_20_2 R_bl
Rbb_20_1 bitb_20_1 bitb_20_2 R_bl
Cb_20_1 bit_20_1 gnd C_bl
Cbb_20_1 bitb_20_1 gnd C_bl
Rb_20_2 bit_20_2 bit_20_3 R_bl
Rbb_20_2 bitb_20_2 bitb_20_3 R_bl
Cb_20_2 bit_20_2 gnd C_bl
Cbb_20_2 bitb_20_2 gnd C_bl
Rb_20_3 bit_20_3 bit_20_4 R_bl
Rbb_20_3 bitb_20_3 bitb_20_4 R_bl
Cb_20_3 bit_20_3 gnd C_bl
Cbb_20_3 bitb_20_3 gnd C_bl
Rb_20_4 bit_20_4 bit_20_5 R_bl
Rbb_20_4 bitb_20_4 bitb_20_5 R_bl
Cb_20_4 bit_20_4 gnd C_bl
Cbb_20_4 bitb_20_4 gnd C_bl
Rb_20_5 bit_20_5 bit_20_6 R_bl
Rbb_20_5 bitb_20_5 bitb_20_6 R_bl
Cb_20_5 bit_20_5 gnd C_bl
Cbb_20_5 bitb_20_5 gnd C_bl
Rb_20_6 bit_20_6 bit_20_7 R_bl
Rbb_20_6 bitb_20_6 bitb_20_7 R_bl
Cb_20_6 bit_20_6 gnd C_bl
Cbb_20_6 bitb_20_6 gnd C_bl
Rb_20_7 bit_20_7 bit_20_8 R_bl
Rbb_20_7 bitb_20_7 bitb_20_8 R_bl
Cb_20_7 bit_20_7 gnd C_bl
Cbb_20_7 bitb_20_7 gnd C_bl
Rb_20_8 bit_20_8 bit_20_9 R_bl
Rbb_20_8 bitb_20_8 bitb_20_9 R_bl
Cb_20_8 bit_20_8 gnd C_bl
Cbb_20_8 bitb_20_8 gnd C_bl
Rb_20_9 bit_20_9 bit_20_10 R_bl
Rbb_20_9 bitb_20_9 bitb_20_10 R_bl
Cb_20_9 bit_20_9 gnd C_bl
Cbb_20_9 bitb_20_9 gnd C_bl
Rb_20_10 bit_20_10 bit_20_11 R_bl
Rbb_20_10 bitb_20_10 bitb_20_11 R_bl
Cb_20_10 bit_20_10 gnd C_bl
Cbb_20_10 bitb_20_10 gnd C_bl
Rb_20_11 bit_20_11 bit_20_12 R_bl
Rbb_20_11 bitb_20_11 bitb_20_12 R_bl
Cb_20_11 bit_20_11 gnd C_bl
Cbb_20_11 bitb_20_11 gnd C_bl
Rb_20_12 bit_20_12 bit_20_13 R_bl
Rbb_20_12 bitb_20_12 bitb_20_13 R_bl
Cb_20_12 bit_20_12 gnd C_bl
Cbb_20_12 bitb_20_12 gnd C_bl
Rb_20_13 bit_20_13 bit_20_14 R_bl
Rbb_20_13 bitb_20_13 bitb_20_14 R_bl
Cb_20_13 bit_20_13 gnd C_bl
Cbb_20_13 bitb_20_13 gnd C_bl
Rb_20_14 bit_20_14 bit_20_15 R_bl
Rbb_20_14 bitb_20_14 bitb_20_15 R_bl
Cb_20_14 bit_20_14 gnd C_bl
Cbb_20_14 bitb_20_14 gnd C_bl
Rb_20_15 bit_20_15 bit_20_16 R_bl
Rbb_20_15 bitb_20_15 bitb_20_16 R_bl
Cb_20_15 bit_20_15 gnd C_bl
Cbb_20_15 bitb_20_15 gnd C_bl
Rb_20_16 bit_20_16 bit_20_17 R_bl
Rbb_20_16 bitb_20_16 bitb_20_17 R_bl
Cb_20_16 bit_20_16 gnd C_bl
Cbb_20_16 bitb_20_16 gnd C_bl
Rb_20_17 bit_20_17 bit_20_18 R_bl
Rbb_20_17 bitb_20_17 bitb_20_18 R_bl
Cb_20_17 bit_20_17 gnd C_bl
Cbb_20_17 bitb_20_17 gnd C_bl
Rb_20_18 bit_20_18 bit_20_19 R_bl
Rbb_20_18 bitb_20_18 bitb_20_19 R_bl
Cb_20_18 bit_20_18 gnd C_bl
Cbb_20_18 bitb_20_18 gnd C_bl
Rb_20_19 bit_20_19 bit_20_20 R_bl
Rbb_20_19 bitb_20_19 bitb_20_20 R_bl
Cb_20_19 bit_20_19 gnd C_bl
Cbb_20_19 bitb_20_19 gnd C_bl
Rb_20_20 bit_20_20 bit_20_21 R_bl
Rbb_20_20 bitb_20_20 bitb_20_21 R_bl
Cb_20_20 bit_20_20 gnd C_bl
Cbb_20_20 bitb_20_20 gnd C_bl
Rb_20_21 bit_20_21 bit_20_22 R_bl
Rbb_20_21 bitb_20_21 bitb_20_22 R_bl
Cb_20_21 bit_20_21 gnd C_bl
Cbb_20_21 bitb_20_21 gnd C_bl
Rb_20_22 bit_20_22 bit_20_23 R_bl
Rbb_20_22 bitb_20_22 bitb_20_23 R_bl
Cb_20_22 bit_20_22 gnd C_bl
Cbb_20_22 bitb_20_22 gnd C_bl
Rb_20_23 bit_20_23 bit_20_24 R_bl
Rbb_20_23 bitb_20_23 bitb_20_24 R_bl
Cb_20_23 bit_20_23 gnd C_bl
Cbb_20_23 bitb_20_23 gnd C_bl
Rb_20_24 bit_20_24 bit_20_25 R_bl
Rbb_20_24 bitb_20_24 bitb_20_25 R_bl
Cb_20_24 bit_20_24 gnd C_bl
Cbb_20_24 bitb_20_24 gnd C_bl
Rb_20_25 bit_20_25 bit_20_26 R_bl
Rbb_20_25 bitb_20_25 bitb_20_26 R_bl
Cb_20_25 bit_20_25 gnd C_bl
Cbb_20_25 bitb_20_25 gnd C_bl
Rb_20_26 bit_20_26 bit_20_27 R_bl
Rbb_20_26 bitb_20_26 bitb_20_27 R_bl
Cb_20_26 bit_20_26 gnd C_bl
Cbb_20_26 bitb_20_26 gnd C_bl
Rb_20_27 bit_20_27 bit_20_28 R_bl
Rbb_20_27 bitb_20_27 bitb_20_28 R_bl
Cb_20_27 bit_20_27 gnd C_bl
Cbb_20_27 bitb_20_27 gnd C_bl
Rb_20_28 bit_20_28 bit_20_29 R_bl
Rbb_20_28 bitb_20_28 bitb_20_29 R_bl
Cb_20_28 bit_20_28 gnd C_bl
Cbb_20_28 bitb_20_28 gnd C_bl
Rb_20_29 bit_20_29 bit_20_30 R_bl
Rbb_20_29 bitb_20_29 bitb_20_30 R_bl
Cb_20_29 bit_20_29 gnd C_bl
Cbb_20_29 bitb_20_29 gnd C_bl
Rb_20_30 bit_20_30 bit_20_31 R_bl
Rbb_20_30 bitb_20_30 bitb_20_31 R_bl
Cb_20_30 bit_20_30 gnd C_bl
Cbb_20_30 bitb_20_30 gnd C_bl
Rb_20_31 bit_20_31 bit_20_32 R_bl
Rbb_20_31 bitb_20_31 bitb_20_32 R_bl
Cb_20_31 bit_20_31 gnd C_bl
Cbb_20_31 bitb_20_31 gnd C_bl
Rb_20_32 bit_20_32 bit_20_33 R_bl
Rbb_20_32 bitb_20_32 bitb_20_33 R_bl
Cb_20_32 bit_20_32 gnd C_bl
Cbb_20_32 bitb_20_32 gnd C_bl
Rb_20_33 bit_20_33 bit_20_34 R_bl
Rbb_20_33 bitb_20_33 bitb_20_34 R_bl
Cb_20_33 bit_20_33 gnd C_bl
Cbb_20_33 bitb_20_33 gnd C_bl
Rb_20_34 bit_20_34 bit_20_35 R_bl
Rbb_20_34 bitb_20_34 bitb_20_35 R_bl
Cb_20_34 bit_20_34 gnd C_bl
Cbb_20_34 bitb_20_34 gnd C_bl
Rb_20_35 bit_20_35 bit_20_36 R_bl
Rbb_20_35 bitb_20_35 bitb_20_36 R_bl
Cb_20_35 bit_20_35 gnd C_bl
Cbb_20_35 bitb_20_35 gnd C_bl
Rb_20_36 bit_20_36 bit_20_37 R_bl
Rbb_20_36 bitb_20_36 bitb_20_37 R_bl
Cb_20_36 bit_20_36 gnd C_bl
Cbb_20_36 bitb_20_36 gnd C_bl
Rb_20_37 bit_20_37 bit_20_38 R_bl
Rbb_20_37 bitb_20_37 bitb_20_38 R_bl
Cb_20_37 bit_20_37 gnd C_bl
Cbb_20_37 bitb_20_37 gnd C_bl
Rb_20_38 bit_20_38 bit_20_39 R_bl
Rbb_20_38 bitb_20_38 bitb_20_39 R_bl
Cb_20_38 bit_20_38 gnd C_bl
Cbb_20_38 bitb_20_38 gnd C_bl
Rb_20_39 bit_20_39 bit_20_40 R_bl
Rbb_20_39 bitb_20_39 bitb_20_40 R_bl
Cb_20_39 bit_20_39 gnd C_bl
Cbb_20_39 bitb_20_39 gnd C_bl
Rb_20_40 bit_20_40 bit_20_41 R_bl
Rbb_20_40 bitb_20_40 bitb_20_41 R_bl
Cb_20_40 bit_20_40 gnd C_bl
Cbb_20_40 bitb_20_40 gnd C_bl
Rb_20_41 bit_20_41 bit_20_42 R_bl
Rbb_20_41 bitb_20_41 bitb_20_42 R_bl
Cb_20_41 bit_20_41 gnd C_bl
Cbb_20_41 bitb_20_41 gnd C_bl
Rb_20_42 bit_20_42 bit_20_43 R_bl
Rbb_20_42 bitb_20_42 bitb_20_43 R_bl
Cb_20_42 bit_20_42 gnd C_bl
Cbb_20_42 bitb_20_42 gnd C_bl
Rb_20_43 bit_20_43 bit_20_44 R_bl
Rbb_20_43 bitb_20_43 bitb_20_44 R_bl
Cb_20_43 bit_20_43 gnd C_bl
Cbb_20_43 bitb_20_43 gnd C_bl
Rb_20_44 bit_20_44 bit_20_45 R_bl
Rbb_20_44 bitb_20_44 bitb_20_45 R_bl
Cb_20_44 bit_20_44 gnd C_bl
Cbb_20_44 bitb_20_44 gnd C_bl
Rb_20_45 bit_20_45 bit_20_46 R_bl
Rbb_20_45 bitb_20_45 bitb_20_46 R_bl
Cb_20_45 bit_20_45 gnd C_bl
Cbb_20_45 bitb_20_45 gnd C_bl
Rb_20_46 bit_20_46 bit_20_47 R_bl
Rbb_20_46 bitb_20_46 bitb_20_47 R_bl
Cb_20_46 bit_20_46 gnd C_bl
Cbb_20_46 bitb_20_46 gnd C_bl
Rb_20_47 bit_20_47 bit_20_48 R_bl
Rbb_20_47 bitb_20_47 bitb_20_48 R_bl
Cb_20_47 bit_20_47 gnd C_bl
Cbb_20_47 bitb_20_47 gnd C_bl
Rb_20_48 bit_20_48 bit_20_49 R_bl
Rbb_20_48 bitb_20_48 bitb_20_49 R_bl
Cb_20_48 bit_20_48 gnd C_bl
Cbb_20_48 bitb_20_48 gnd C_bl
Rb_20_49 bit_20_49 bit_20_50 R_bl
Rbb_20_49 bitb_20_49 bitb_20_50 R_bl
Cb_20_49 bit_20_49 gnd C_bl
Cbb_20_49 bitb_20_49 gnd C_bl
Rb_20_50 bit_20_50 bit_20_51 R_bl
Rbb_20_50 bitb_20_50 bitb_20_51 R_bl
Cb_20_50 bit_20_50 gnd C_bl
Cbb_20_50 bitb_20_50 gnd C_bl
Rb_20_51 bit_20_51 bit_20_52 R_bl
Rbb_20_51 bitb_20_51 bitb_20_52 R_bl
Cb_20_51 bit_20_51 gnd C_bl
Cbb_20_51 bitb_20_51 gnd C_bl
Rb_20_52 bit_20_52 bit_20_53 R_bl
Rbb_20_52 bitb_20_52 bitb_20_53 R_bl
Cb_20_52 bit_20_52 gnd C_bl
Cbb_20_52 bitb_20_52 gnd C_bl
Rb_20_53 bit_20_53 bit_20_54 R_bl
Rbb_20_53 bitb_20_53 bitb_20_54 R_bl
Cb_20_53 bit_20_53 gnd C_bl
Cbb_20_53 bitb_20_53 gnd C_bl
Rb_20_54 bit_20_54 bit_20_55 R_bl
Rbb_20_54 bitb_20_54 bitb_20_55 R_bl
Cb_20_54 bit_20_54 gnd C_bl
Cbb_20_54 bitb_20_54 gnd C_bl
Rb_20_55 bit_20_55 bit_20_56 R_bl
Rbb_20_55 bitb_20_55 bitb_20_56 R_bl
Cb_20_55 bit_20_55 gnd C_bl
Cbb_20_55 bitb_20_55 gnd C_bl
Rb_20_56 bit_20_56 bit_20_57 R_bl
Rbb_20_56 bitb_20_56 bitb_20_57 R_bl
Cb_20_56 bit_20_56 gnd C_bl
Cbb_20_56 bitb_20_56 gnd C_bl
Rb_20_57 bit_20_57 bit_20_58 R_bl
Rbb_20_57 bitb_20_57 bitb_20_58 R_bl
Cb_20_57 bit_20_57 gnd C_bl
Cbb_20_57 bitb_20_57 gnd C_bl
Rb_20_58 bit_20_58 bit_20_59 R_bl
Rbb_20_58 bitb_20_58 bitb_20_59 R_bl
Cb_20_58 bit_20_58 gnd C_bl
Cbb_20_58 bitb_20_58 gnd C_bl
Rb_20_59 bit_20_59 bit_20_60 R_bl
Rbb_20_59 bitb_20_59 bitb_20_60 R_bl
Cb_20_59 bit_20_59 gnd C_bl
Cbb_20_59 bitb_20_59 gnd C_bl
Rb_20_60 bit_20_60 bit_20_61 R_bl
Rbb_20_60 bitb_20_60 bitb_20_61 R_bl
Cb_20_60 bit_20_60 gnd C_bl
Cbb_20_60 bitb_20_60 gnd C_bl
Rb_20_61 bit_20_61 bit_20_62 R_bl
Rbb_20_61 bitb_20_61 bitb_20_62 R_bl
Cb_20_61 bit_20_61 gnd C_bl
Cbb_20_61 bitb_20_61 gnd C_bl
Rb_20_62 bit_20_62 bit_20_63 R_bl
Rbb_20_62 bitb_20_62 bitb_20_63 R_bl
Cb_20_62 bit_20_62 gnd C_bl
Cbb_20_62 bitb_20_62 gnd C_bl
Rb_20_63 bit_20_63 bit_20_64 R_bl
Rbb_20_63 bitb_20_63 bitb_20_64 R_bl
Cb_20_63 bit_20_63 gnd C_bl
Cbb_20_63 bitb_20_63 gnd C_bl
Rb_20_64 bit_20_64 bit_20_65 R_bl
Rbb_20_64 bitb_20_64 bitb_20_65 R_bl
Cb_20_64 bit_20_64 gnd C_bl
Cbb_20_64 bitb_20_64 gnd C_bl
Rb_20_65 bit_20_65 bit_20_66 R_bl
Rbb_20_65 bitb_20_65 bitb_20_66 R_bl
Cb_20_65 bit_20_65 gnd C_bl
Cbb_20_65 bitb_20_65 gnd C_bl
Rb_20_66 bit_20_66 bit_20_67 R_bl
Rbb_20_66 bitb_20_66 bitb_20_67 R_bl
Cb_20_66 bit_20_66 gnd C_bl
Cbb_20_66 bitb_20_66 gnd C_bl
Rb_20_67 bit_20_67 bit_20_68 R_bl
Rbb_20_67 bitb_20_67 bitb_20_68 R_bl
Cb_20_67 bit_20_67 gnd C_bl
Cbb_20_67 bitb_20_67 gnd C_bl
Rb_20_68 bit_20_68 bit_20_69 R_bl
Rbb_20_68 bitb_20_68 bitb_20_69 R_bl
Cb_20_68 bit_20_68 gnd C_bl
Cbb_20_68 bitb_20_68 gnd C_bl
Rb_20_69 bit_20_69 bit_20_70 R_bl
Rbb_20_69 bitb_20_69 bitb_20_70 R_bl
Cb_20_69 bit_20_69 gnd C_bl
Cbb_20_69 bitb_20_69 gnd C_bl
Rb_20_70 bit_20_70 bit_20_71 R_bl
Rbb_20_70 bitb_20_70 bitb_20_71 R_bl
Cb_20_70 bit_20_70 gnd C_bl
Cbb_20_70 bitb_20_70 gnd C_bl
Rb_20_71 bit_20_71 bit_20_72 R_bl
Rbb_20_71 bitb_20_71 bitb_20_72 R_bl
Cb_20_71 bit_20_71 gnd C_bl
Cbb_20_71 bitb_20_71 gnd C_bl
Rb_20_72 bit_20_72 bit_20_73 R_bl
Rbb_20_72 bitb_20_72 bitb_20_73 R_bl
Cb_20_72 bit_20_72 gnd C_bl
Cbb_20_72 bitb_20_72 gnd C_bl
Rb_20_73 bit_20_73 bit_20_74 R_bl
Rbb_20_73 bitb_20_73 bitb_20_74 R_bl
Cb_20_73 bit_20_73 gnd C_bl
Cbb_20_73 bitb_20_73 gnd C_bl
Rb_20_74 bit_20_74 bit_20_75 R_bl
Rbb_20_74 bitb_20_74 bitb_20_75 R_bl
Cb_20_74 bit_20_74 gnd C_bl
Cbb_20_74 bitb_20_74 gnd C_bl
Rb_20_75 bit_20_75 bit_20_76 R_bl
Rbb_20_75 bitb_20_75 bitb_20_76 R_bl
Cb_20_75 bit_20_75 gnd C_bl
Cbb_20_75 bitb_20_75 gnd C_bl
Rb_20_76 bit_20_76 bit_20_77 R_bl
Rbb_20_76 bitb_20_76 bitb_20_77 R_bl
Cb_20_76 bit_20_76 gnd C_bl
Cbb_20_76 bitb_20_76 gnd C_bl
Rb_20_77 bit_20_77 bit_20_78 R_bl
Rbb_20_77 bitb_20_77 bitb_20_78 R_bl
Cb_20_77 bit_20_77 gnd C_bl
Cbb_20_77 bitb_20_77 gnd C_bl
Rb_20_78 bit_20_78 bit_20_79 R_bl
Rbb_20_78 bitb_20_78 bitb_20_79 R_bl
Cb_20_78 bit_20_78 gnd C_bl
Cbb_20_78 bitb_20_78 gnd C_bl
Rb_20_79 bit_20_79 bit_20_80 R_bl
Rbb_20_79 bitb_20_79 bitb_20_80 R_bl
Cb_20_79 bit_20_79 gnd C_bl
Cbb_20_79 bitb_20_79 gnd C_bl
Rb_20_80 bit_20_80 bit_20_81 R_bl
Rbb_20_80 bitb_20_80 bitb_20_81 R_bl
Cb_20_80 bit_20_80 gnd C_bl
Cbb_20_80 bitb_20_80 gnd C_bl
Rb_20_81 bit_20_81 bit_20_82 R_bl
Rbb_20_81 bitb_20_81 bitb_20_82 R_bl
Cb_20_81 bit_20_81 gnd C_bl
Cbb_20_81 bitb_20_81 gnd C_bl
Rb_20_82 bit_20_82 bit_20_83 R_bl
Rbb_20_82 bitb_20_82 bitb_20_83 R_bl
Cb_20_82 bit_20_82 gnd C_bl
Cbb_20_82 bitb_20_82 gnd C_bl
Rb_20_83 bit_20_83 bit_20_84 R_bl
Rbb_20_83 bitb_20_83 bitb_20_84 R_bl
Cb_20_83 bit_20_83 gnd C_bl
Cbb_20_83 bitb_20_83 gnd C_bl
Rb_20_84 bit_20_84 bit_20_85 R_bl
Rbb_20_84 bitb_20_84 bitb_20_85 R_bl
Cb_20_84 bit_20_84 gnd C_bl
Cbb_20_84 bitb_20_84 gnd C_bl
Rb_20_85 bit_20_85 bit_20_86 R_bl
Rbb_20_85 bitb_20_85 bitb_20_86 R_bl
Cb_20_85 bit_20_85 gnd C_bl
Cbb_20_85 bitb_20_85 gnd C_bl
Rb_20_86 bit_20_86 bit_20_87 R_bl
Rbb_20_86 bitb_20_86 bitb_20_87 R_bl
Cb_20_86 bit_20_86 gnd C_bl
Cbb_20_86 bitb_20_86 gnd C_bl
Rb_20_87 bit_20_87 bit_20_88 R_bl
Rbb_20_87 bitb_20_87 bitb_20_88 R_bl
Cb_20_87 bit_20_87 gnd C_bl
Cbb_20_87 bitb_20_87 gnd C_bl
Rb_20_88 bit_20_88 bit_20_89 R_bl
Rbb_20_88 bitb_20_88 bitb_20_89 R_bl
Cb_20_88 bit_20_88 gnd C_bl
Cbb_20_88 bitb_20_88 gnd C_bl
Rb_20_89 bit_20_89 bit_20_90 R_bl
Rbb_20_89 bitb_20_89 bitb_20_90 R_bl
Cb_20_89 bit_20_89 gnd C_bl
Cbb_20_89 bitb_20_89 gnd C_bl
Rb_20_90 bit_20_90 bit_20_91 R_bl
Rbb_20_90 bitb_20_90 bitb_20_91 R_bl
Cb_20_90 bit_20_90 gnd C_bl
Cbb_20_90 bitb_20_90 gnd C_bl
Rb_20_91 bit_20_91 bit_20_92 R_bl
Rbb_20_91 bitb_20_91 bitb_20_92 R_bl
Cb_20_91 bit_20_91 gnd C_bl
Cbb_20_91 bitb_20_91 gnd C_bl
Rb_20_92 bit_20_92 bit_20_93 R_bl
Rbb_20_92 bitb_20_92 bitb_20_93 R_bl
Cb_20_92 bit_20_92 gnd C_bl
Cbb_20_92 bitb_20_92 gnd C_bl
Rb_20_93 bit_20_93 bit_20_94 R_bl
Rbb_20_93 bitb_20_93 bitb_20_94 R_bl
Cb_20_93 bit_20_93 gnd C_bl
Cbb_20_93 bitb_20_93 gnd C_bl
Rb_20_94 bit_20_94 bit_20_95 R_bl
Rbb_20_94 bitb_20_94 bitb_20_95 R_bl
Cb_20_94 bit_20_94 gnd C_bl
Cbb_20_94 bitb_20_94 gnd C_bl
Rb_20_95 bit_20_95 bit_20_96 R_bl
Rbb_20_95 bitb_20_95 bitb_20_96 R_bl
Cb_20_95 bit_20_95 gnd C_bl
Cbb_20_95 bitb_20_95 gnd C_bl
Rb_20_96 bit_20_96 bit_20_97 R_bl
Rbb_20_96 bitb_20_96 bitb_20_97 R_bl
Cb_20_96 bit_20_96 gnd C_bl
Cbb_20_96 bitb_20_96 gnd C_bl
Rb_20_97 bit_20_97 bit_20_98 R_bl
Rbb_20_97 bitb_20_97 bitb_20_98 R_bl
Cb_20_97 bit_20_97 gnd C_bl
Cbb_20_97 bitb_20_97 gnd C_bl
Rb_20_98 bit_20_98 bit_20_99 R_bl
Rbb_20_98 bitb_20_98 bitb_20_99 R_bl
Cb_20_98 bit_20_98 gnd C_bl
Cbb_20_98 bitb_20_98 gnd C_bl
Rb_20_99 bit_20_99 bit_20_100 R_bl
Rbb_20_99 bitb_20_99 bitb_20_100 R_bl
Cb_20_99 bit_20_99 gnd C_bl
Cbb_20_99 bitb_20_99 gnd C_bl
Rb_21_0 bit_21_0 bit_21_1 R_bl
Rbb_21_0 bitb_21_0 bitb_21_1 R_bl
Cb_21_0 bit_21_0 gnd C_bl
Cbb_21_0 bitb_21_0 gnd C_bl
Rb_21_1 bit_21_1 bit_21_2 R_bl
Rbb_21_1 bitb_21_1 bitb_21_2 R_bl
Cb_21_1 bit_21_1 gnd C_bl
Cbb_21_1 bitb_21_1 gnd C_bl
Rb_21_2 bit_21_2 bit_21_3 R_bl
Rbb_21_2 bitb_21_2 bitb_21_3 R_bl
Cb_21_2 bit_21_2 gnd C_bl
Cbb_21_2 bitb_21_2 gnd C_bl
Rb_21_3 bit_21_3 bit_21_4 R_bl
Rbb_21_3 bitb_21_3 bitb_21_4 R_bl
Cb_21_3 bit_21_3 gnd C_bl
Cbb_21_3 bitb_21_3 gnd C_bl
Rb_21_4 bit_21_4 bit_21_5 R_bl
Rbb_21_4 bitb_21_4 bitb_21_5 R_bl
Cb_21_4 bit_21_4 gnd C_bl
Cbb_21_4 bitb_21_4 gnd C_bl
Rb_21_5 bit_21_5 bit_21_6 R_bl
Rbb_21_5 bitb_21_5 bitb_21_6 R_bl
Cb_21_5 bit_21_5 gnd C_bl
Cbb_21_5 bitb_21_5 gnd C_bl
Rb_21_6 bit_21_6 bit_21_7 R_bl
Rbb_21_6 bitb_21_6 bitb_21_7 R_bl
Cb_21_6 bit_21_6 gnd C_bl
Cbb_21_6 bitb_21_6 gnd C_bl
Rb_21_7 bit_21_7 bit_21_8 R_bl
Rbb_21_7 bitb_21_7 bitb_21_8 R_bl
Cb_21_7 bit_21_7 gnd C_bl
Cbb_21_7 bitb_21_7 gnd C_bl
Rb_21_8 bit_21_8 bit_21_9 R_bl
Rbb_21_8 bitb_21_8 bitb_21_9 R_bl
Cb_21_8 bit_21_8 gnd C_bl
Cbb_21_8 bitb_21_8 gnd C_bl
Rb_21_9 bit_21_9 bit_21_10 R_bl
Rbb_21_9 bitb_21_9 bitb_21_10 R_bl
Cb_21_9 bit_21_9 gnd C_bl
Cbb_21_9 bitb_21_9 gnd C_bl
Rb_21_10 bit_21_10 bit_21_11 R_bl
Rbb_21_10 bitb_21_10 bitb_21_11 R_bl
Cb_21_10 bit_21_10 gnd C_bl
Cbb_21_10 bitb_21_10 gnd C_bl
Rb_21_11 bit_21_11 bit_21_12 R_bl
Rbb_21_11 bitb_21_11 bitb_21_12 R_bl
Cb_21_11 bit_21_11 gnd C_bl
Cbb_21_11 bitb_21_11 gnd C_bl
Rb_21_12 bit_21_12 bit_21_13 R_bl
Rbb_21_12 bitb_21_12 bitb_21_13 R_bl
Cb_21_12 bit_21_12 gnd C_bl
Cbb_21_12 bitb_21_12 gnd C_bl
Rb_21_13 bit_21_13 bit_21_14 R_bl
Rbb_21_13 bitb_21_13 bitb_21_14 R_bl
Cb_21_13 bit_21_13 gnd C_bl
Cbb_21_13 bitb_21_13 gnd C_bl
Rb_21_14 bit_21_14 bit_21_15 R_bl
Rbb_21_14 bitb_21_14 bitb_21_15 R_bl
Cb_21_14 bit_21_14 gnd C_bl
Cbb_21_14 bitb_21_14 gnd C_bl
Rb_21_15 bit_21_15 bit_21_16 R_bl
Rbb_21_15 bitb_21_15 bitb_21_16 R_bl
Cb_21_15 bit_21_15 gnd C_bl
Cbb_21_15 bitb_21_15 gnd C_bl
Rb_21_16 bit_21_16 bit_21_17 R_bl
Rbb_21_16 bitb_21_16 bitb_21_17 R_bl
Cb_21_16 bit_21_16 gnd C_bl
Cbb_21_16 bitb_21_16 gnd C_bl
Rb_21_17 bit_21_17 bit_21_18 R_bl
Rbb_21_17 bitb_21_17 bitb_21_18 R_bl
Cb_21_17 bit_21_17 gnd C_bl
Cbb_21_17 bitb_21_17 gnd C_bl
Rb_21_18 bit_21_18 bit_21_19 R_bl
Rbb_21_18 bitb_21_18 bitb_21_19 R_bl
Cb_21_18 bit_21_18 gnd C_bl
Cbb_21_18 bitb_21_18 gnd C_bl
Rb_21_19 bit_21_19 bit_21_20 R_bl
Rbb_21_19 bitb_21_19 bitb_21_20 R_bl
Cb_21_19 bit_21_19 gnd C_bl
Cbb_21_19 bitb_21_19 gnd C_bl
Rb_21_20 bit_21_20 bit_21_21 R_bl
Rbb_21_20 bitb_21_20 bitb_21_21 R_bl
Cb_21_20 bit_21_20 gnd C_bl
Cbb_21_20 bitb_21_20 gnd C_bl
Rb_21_21 bit_21_21 bit_21_22 R_bl
Rbb_21_21 bitb_21_21 bitb_21_22 R_bl
Cb_21_21 bit_21_21 gnd C_bl
Cbb_21_21 bitb_21_21 gnd C_bl
Rb_21_22 bit_21_22 bit_21_23 R_bl
Rbb_21_22 bitb_21_22 bitb_21_23 R_bl
Cb_21_22 bit_21_22 gnd C_bl
Cbb_21_22 bitb_21_22 gnd C_bl
Rb_21_23 bit_21_23 bit_21_24 R_bl
Rbb_21_23 bitb_21_23 bitb_21_24 R_bl
Cb_21_23 bit_21_23 gnd C_bl
Cbb_21_23 bitb_21_23 gnd C_bl
Rb_21_24 bit_21_24 bit_21_25 R_bl
Rbb_21_24 bitb_21_24 bitb_21_25 R_bl
Cb_21_24 bit_21_24 gnd C_bl
Cbb_21_24 bitb_21_24 gnd C_bl
Rb_21_25 bit_21_25 bit_21_26 R_bl
Rbb_21_25 bitb_21_25 bitb_21_26 R_bl
Cb_21_25 bit_21_25 gnd C_bl
Cbb_21_25 bitb_21_25 gnd C_bl
Rb_21_26 bit_21_26 bit_21_27 R_bl
Rbb_21_26 bitb_21_26 bitb_21_27 R_bl
Cb_21_26 bit_21_26 gnd C_bl
Cbb_21_26 bitb_21_26 gnd C_bl
Rb_21_27 bit_21_27 bit_21_28 R_bl
Rbb_21_27 bitb_21_27 bitb_21_28 R_bl
Cb_21_27 bit_21_27 gnd C_bl
Cbb_21_27 bitb_21_27 gnd C_bl
Rb_21_28 bit_21_28 bit_21_29 R_bl
Rbb_21_28 bitb_21_28 bitb_21_29 R_bl
Cb_21_28 bit_21_28 gnd C_bl
Cbb_21_28 bitb_21_28 gnd C_bl
Rb_21_29 bit_21_29 bit_21_30 R_bl
Rbb_21_29 bitb_21_29 bitb_21_30 R_bl
Cb_21_29 bit_21_29 gnd C_bl
Cbb_21_29 bitb_21_29 gnd C_bl
Rb_21_30 bit_21_30 bit_21_31 R_bl
Rbb_21_30 bitb_21_30 bitb_21_31 R_bl
Cb_21_30 bit_21_30 gnd C_bl
Cbb_21_30 bitb_21_30 gnd C_bl
Rb_21_31 bit_21_31 bit_21_32 R_bl
Rbb_21_31 bitb_21_31 bitb_21_32 R_bl
Cb_21_31 bit_21_31 gnd C_bl
Cbb_21_31 bitb_21_31 gnd C_bl
Rb_21_32 bit_21_32 bit_21_33 R_bl
Rbb_21_32 bitb_21_32 bitb_21_33 R_bl
Cb_21_32 bit_21_32 gnd C_bl
Cbb_21_32 bitb_21_32 gnd C_bl
Rb_21_33 bit_21_33 bit_21_34 R_bl
Rbb_21_33 bitb_21_33 bitb_21_34 R_bl
Cb_21_33 bit_21_33 gnd C_bl
Cbb_21_33 bitb_21_33 gnd C_bl
Rb_21_34 bit_21_34 bit_21_35 R_bl
Rbb_21_34 bitb_21_34 bitb_21_35 R_bl
Cb_21_34 bit_21_34 gnd C_bl
Cbb_21_34 bitb_21_34 gnd C_bl
Rb_21_35 bit_21_35 bit_21_36 R_bl
Rbb_21_35 bitb_21_35 bitb_21_36 R_bl
Cb_21_35 bit_21_35 gnd C_bl
Cbb_21_35 bitb_21_35 gnd C_bl
Rb_21_36 bit_21_36 bit_21_37 R_bl
Rbb_21_36 bitb_21_36 bitb_21_37 R_bl
Cb_21_36 bit_21_36 gnd C_bl
Cbb_21_36 bitb_21_36 gnd C_bl
Rb_21_37 bit_21_37 bit_21_38 R_bl
Rbb_21_37 bitb_21_37 bitb_21_38 R_bl
Cb_21_37 bit_21_37 gnd C_bl
Cbb_21_37 bitb_21_37 gnd C_bl
Rb_21_38 bit_21_38 bit_21_39 R_bl
Rbb_21_38 bitb_21_38 bitb_21_39 R_bl
Cb_21_38 bit_21_38 gnd C_bl
Cbb_21_38 bitb_21_38 gnd C_bl
Rb_21_39 bit_21_39 bit_21_40 R_bl
Rbb_21_39 bitb_21_39 bitb_21_40 R_bl
Cb_21_39 bit_21_39 gnd C_bl
Cbb_21_39 bitb_21_39 gnd C_bl
Rb_21_40 bit_21_40 bit_21_41 R_bl
Rbb_21_40 bitb_21_40 bitb_21_41 R_bl
Cb_21_40 bit_21_40 gnd C_bl
Cbb_21_40 bitb_21_40 gnd C_bl
Rb_21_41 bit_21_41 bit_21_42 R_bl
Rbb_21_41 bitb_21_41 bitb_21_42 R_bl
Cb_21_41 bit_21_41 gnd C_bl
Cbb_21_41 bitb_21_41 gnd C_bl
Rb_21_42 bit_21_42 bit_21_43 R_bl
Rbb_21_42 bitb_21_42 bitb_21_43 R_bl
Cb_21_42 bit_21_42 gnd C_bl
Cbb_21_42 bitb_21_42 gnd C_bl
Rb_21_43 bit_21_43 bit_21_44 R_bl
Rbb_21_43 bitb_21_43 bitb_21_44 R_bl
Cb_21_43 bit_21_43 gnd C_bl
Cbb_21_43 bitb_21_43 gnd C_bl
Rb_21_44 bit_21_44 bit_21_45 R_bl
Rbb_21_44 bitb_21_44 bitb_21_45 R_bl
Cb_21_44 bit_21_44 gnd C_bl
Cbb_21_44 bitb_21_44 gnd C_bl
Rb_21_45 bit_21_45 bit_21_46 R_bl
Rbb_21_45 bitb_21_45 bitb_21_46 R_bl
Cb_21_45 bit_21_45 gnd C_bl
Cbb_21_45 bitb_21_45 gnd C_bl
Rb_21_46 bit_21_46 bit_21_47 R_bl
Rbb_21_46 bitb_21_46 bitb_21_47 R_bl
Cb_21_46 bit_21_46 gnd C_bl
Cbb_21_46 bitb_21_46 gnd C_bl
Rb_21_47 bit_21_47 bit_21_48 R_bl
Rbb_21_47 bitb_21_47 bitb_21_48 R_bl
Cb_21_47 bit_21_47 gnd C_bl
Cbb_21_47 bitb_21_47 gnd C_bl
Rb_21_48 bit_21_48 bit_21_49 R_bl
Rbb_21_48 bitb_21_48 bitb_21_49 R_bl
Cb_21_48 bit_21_48 gnd C_bl
Cbb_21_48 bitb_21_48 gnd C_bl
Rb_21_49 bit_21_49 bit_21_50 R_bl
Rbb_21_49 bitb_21_49 bitb_21_50 R_bl
Cb_21_49 bit_21_49 gnd C_bl
Cbb_21_49 bitb_21_49 gnd C_bl
Rb_21_50 bit_21_50 bit_21_51 R_bl
Rbb_21_50 bitb_21_50 bitb_21_51 R_bl
Cb_21_50 bit_21_50 gnd C_bl
Cbb_21_50 bitb_21_50 gnd C_bl
Rb_21_51 bit_21_51 bit_21_52 R_bl
Rbb_21_51 bitb_21_51 bitb_21_52 R_bl
Cb_21_51 bit_21_51 gnd C_bl
Cbb_21_51 bitb_21_51 gnd C_bl
Rb_21_52 bit_21_52 bit_21_53 R_bl
Rbb_21_52 bitb_21_52 bitb_21_53 R_bl
Cb_21_52 bit_21_52 gnd C_bl
Cbb_21_52 bitb_21_52 gnd C_bl
Rb_21_53 bit_21_53 bit_21_54 R_bl
Rbb_21_53 bitb_21_53 bitb_21_54 R_bl
Cb_21_53 bit_21_53 gnd C_bl
Cbb_21_53 bitb_21_53 gnd C_bl
Rb_21_54 bit_21_54 bit_21_55 R_bl
Rbb_21_54 bitb_21_54 bitb_21_55 R_bl
Cb_21_54 bit_21_54 gnd C_bl
Cbb_21_54 bitb_21_54 gnd C_bl
Rb_21_55 bit_21_55 bit_21_56 R_bl
Rbb_21_55 bitb_21_55 bitb_21_56 R_bl
Cb_21_55 bit_21_55 gnd C_bl
Cbb_21_55 bitb_21_55 gnd C_bl
Rb_21_56 bit_21_56 bit_21_57 R_bl
Rbb_21_56 bitb_21_56 bitb_21_57 R_bl
Cb_21_56 bit_21_56 gnd C_bl
Cbb_21_56 bitb_21_56 gnd C_bl
Rb_21_57 bit_21_57 bit_21_58 R_bl
Rbb_21_57 bitb_21_57 bitb_21_58 R_bl
Cb_21_57 bit_21_57 gnd C_bl
Cbb_21_57 bitb_21_57 gnd C_bl
Rb_21_58 bit_21_58 bit_21_59 R_bl
Rbb_21_58 bitb_21_58 bitb_21_59 R_bl
Cb_21_58 bit_21_58 gnd C_bl
Cbb_21_58 bitb_21_58 gnd C_bl
Rb_21_59 bit_21_59 bit_21_60 R_bl
Rbb_21_59 bitb_21_59 bitb_21_60 R_bl
Cb_21_59 bit_21_59 gnd C_bl
Cbb_21_59 bitb_21_59 gnd C_bl
Rb_21_60 bit_21_60 bit_21_61 R_bl
Rbb_21_60 bitb_21_60 bitb_21_61 R_bl
Cb_21_60 bit_21_60 gnd C_bl
Cbb_21_60 bitb_21_60 gnd C_bl
Rb_21_61 bit_21_61 bit_21_62 R_bl
Rbb_21_61 bitb_21_61 bitb_21_62 R_bl
Cb_21_61 bit_21_61 gnd C_bl
Cbb_21_61 bitb_21_61 gnd C_bl
Rb_21_62 bit_21_62 bit_21_63 R_bl
Rbb_21_62 bitb_21_62 bitb_21_63 R_bl
Cb_21_62 bit_21_62 gnd C_bl
Cbb_21_62 bitb_21_62 gnd C_bl
Rb_21_63 bit_21_63 bit_21_64 R_bl
Rbb_21_63 bitb_21_63 bitb_21_64 R_bl
Cb_21_63 bit_21_63 gnd C_bl
Cbb_21_63 bitb_21_63 gnd C_bl
Rb_21_64 bit_21_64 bit_21_65 R_bl
Rbb_21_64 bitb_21_64 bitb_21_65 R_bl
Cb_21_64 bit_21_64 gnd C_bl
Cbb_21_64 bitb_21_64 gnd C_bl
Rb_21_65 bit_21_65 bit_21_66 R_bl
Rbb_21_65 bitb_21_65 bitb_21_66 R_bl
Cb_21_65 bit_21_65 gnd C_bl
Cbb_21_65 bitb_21_65 gnd C_bl
Rb_21_66 bit_21_66 bit_21_67 R_bl
Rbb_21_66 bitb_21_66 bitb_21_67 R_bl
Cb_21_66 bit_21_66 gnd C_bl
Cbb_21_66 bitb_21_66 gnd C_bl
Rb_21_67 bit_21_67 bit_21_68 R_bl
Rbb_21_67 bitb_21_67 bitb_21_68 R_bl
Cb_21_67 bit_21_67 gnd C_bl
Cbb_21_67 bitb_21_67 gnd C_bl
Rb_21_68 bit_21_68 bit_21_69 R_bl
Rbb_21_68 bitb_21_68 bitb_21_69 R_bl
Cb_21_68 bit_21_68 gnd C_bl
Cbb_21_68 bitb_21_68 gnd C_bl
Rb_21_69 bit_21_69 bit_21_70 R_bl
Rbb_21_69 bitb_21_69 bitb_21_70 R_bl
Cb_21_69 bit_21_69 gnd C_bl
Cbb_21_69 bitb_21_69 gnd C_bl
Rb_21_70 bit_21_70 bit_21_71 R_bl
Rbb_21_70 bitb_21_70 bitb_21_71 R_bl
Cb_21_70 bit_21_70 gnd C_bl
Cbb_21_70 bitb_21_70 gnd C_bl
Rb_21_71 bit_21_71 bit_21_72 R_bl
Rbb_21_71 bitb_21_71 bitb_21_72 R_bl
Cb_21_71 bit_21_71 gnd C_bl
Cbb_21_71 bitb_21_71 gnd C_bl
Rb_21_72 bit_21_72 bit_21_73 R_bl
Rbb_21_72 bitb_21_72 bitb_21_73 R_bl
Cb_21_72 bit_21_72 gnd C_bl
Cbb_21_72 bitb_21_72 gnd C_bl
Rb_21_73 bit_21_73 bit_21_74 R_bl
Rbb_21_73 bitb_21_73 bitb_21_74 R_bl
Cb_21_73 bit_21_73 gnd C_bl
Cbb_21_73 bitb_21_73 gnd C_bl
Rb_21_74 bit_21_74 bit_21_75 R_bl
Rbb_21_74 bitb_21_74 bitb_21_75 R_bl
Cb_21_74 bit_21_74 gnd C_bl
Cbb_21_74 bitb_21_74 gnd C_bl
Rb_21_75 bit_21_75 bit_21_76 R_bl
Rbb_21_75 bitb_21_75 bitb_21_76 R_bl
Cb_21_75 bit_21_75 gnd C_bl
Cbb_21_75 bitb_21_75 gnd C_bl
Rb_21_76 bit_21_76 bit_21_77 R_bl
Rbb_21_76 bitb_21_76 bitb_21_77 R_bl
Cb_21_76 bit_21_76 gnd C_bl
Cbb_21_76 bitb_21_76 gnd C_bl
Rb_21_77 bit_21_77 bit_21_78 R_bl
Rbb_21_77 bitb_21_77 bitb_21_78 R_bl
Cb_21_77 bit_21_77 gnd C_bl
Cbb_21_77 bitb_21_77 gnd C_bl
Rb_21_78 bit_21_78 bit_21_79 R_bl
Rbb_21_78 bitb_21_78 bitb_21_79 R_bl
Cb_21_78 bit_21_78 gnd C_bl
Cbb_21_78 bitb_21_78 gnd C_bl
Rb_21_79 bit_21_79 bit_21_80 R_bl
Rbb_21_79 bitb_21_79 bitb_21_80 R_bl
Cb_21_79 bit_21_79 gnd C_bl
Cbb_21_79 bitb_21_79 gnd C_bl
Rb_21_80 bit_21_80 bit_21_81 R_bl
Rbb_21_80 bitb_21_80 bitb_21_81 R_bl
Cb_21_80 bit_21_80 gnd C_bl
Cbb_21_80 bitb_21_80 gnd C_bl
Rb_21_81 bit_21_81 bit_21_82 R_bl
Rbb_21_81 bitb_21_81 bitb_21_82 R_bl
Cb_21_81 bit_21_81 gnd C_bl
Cbb_21_81 bitb_21_81 gnd C_bl
Rb_21_82 bit_21_82 bit_21_83 R_bl
Rbb_21_82 bitb_21_82 bitb_21_83 R_bl
Cb_21_82 bit_21_82 gnd C_bl
Cbb_21_82 bitb_21_82 gnd C_bl
Rb_21_83 bit_21_83 bit_21_84 R_bl
Rbb_21_83 bitb_21_83 bitb_21_84 R_bl
Cb_21_83 bit_21_83 gnd C_bl
Cbb_21_83 bitb_21_83 gnd C_bl
Rb_21_84 bit_21_84 bit_21_85 R_bl
Rbb_21_84 bitb_21_84 bitb_21_85 R_bl
Cb_21_84 bit_21_84 gnd C_bl
Cbb_21_84 bitb_21_84 gnd C_bl
Rb_21_85 bit_21_85 bit_21_86 R_bl
Rbb_21_85 bitb_21_85 bitb_21_86 R_bl
Cb_21_85 bit_21_85 gnd C_bl
Cbb_21_85 bitb_21_85 gnd C_bl
Rb_21_86 bit_21_86 bit_21_87 R_bl
Rbb_21_86 bitb_21_86 bitb_21_87 R_bl
Cb_21_86 bit_21_86 gnd C_bl
Cbb_21_86 bitb_21_86 gnd C_bl
Rb_21_87 bit_21_87 bit_21_88 R_bl
Rbb_21_87 bitb_21_87 bitb_21_88 R_bl
Cb_21_87 bit_21_87 gnd C_bl
Cbb_21_87 bitb_21_87 gnd C_bl
Rb_21_88 bit_21_88 bit_21_89 R_bl
Rbb_21_88 bitb_21_88 bitb_21_89 R_bl
Cb_21_88 bit_21_88 gnd C_bl
Cbb_21_88 bitb_21_88 gnd C_bl
Rb_21_89 bit_21_89 bit_21_90 R_bl
Rbb_21_89 bitb_21_89 bitb_21_90 R_bl
Cb_21_89 bit_21_89 gnd C_bl
Cbb_21_89 bitb_21_89 gnd C_bl
Rb_21_90 bit_21_90 bit_21_91 R_bl
Rbb_21_90 bitb_21_90 bitb_21_91 R_bl
Cb_21_90 bit_21_90 gnd C_bl
Cbb_21_90 bitb_21_90 gnd C_bl
Rb_21_91 bit_21_91 bit_21_92 R_bl
Rbb_21_91 bitb_21_91 bitb_21_92 R_bl
Cb_21_91 bit_21_91 gnd C_bl
Cbb_21_91 bitb_21_91 gnd C_bl
Rb_21_92 bit_21_92 bit_21_93 R_bl
Rbb_21_92 bitb_21_92 bitb_21_93 R_bl
Cb_21_92 bit_21_92 gnd C_bl
Cbb_21_92 bitb_21_92 gnd C_bl
Rb_21_93 bit_21_93 bit_21_94 R_bl
Rbb_21_93 bitb_21_93 bitb_21_94 R_bl
Cb_21_93 bit_21_93 gnd C_bl
Cbb_21_93 bitb_21_93 gnd C_bl
Rb_21_94 bit_21_94 bit_21_95 R_bl
Rbb_21_94 bitb_21_94 bitb_21_95 R_bl
Cb_21_94 bit_21_94 gnd C_bl
Cbb_21_94 bitb_21_94 gnd C_bl
Rb_21_95 bit_21_95 bit_21_96 R_bl
Rbb_21_95 bitb_21_95 bitb_21_96 R_bl
Cb_21_95 bit_21_95 gnd C_bl
Cbb_21_95 bitb_21_95 gnd C_bl
Rb_21_96 bit_21_96 bit_21_97 R_bl
Rbb_21_96 bitb_21_96 bitb_21_97 R_bl
Cb_21_96 bit_21_96 gnd C_bl
Cbb_21_96 bitb_21_96 gnd C_bl
Rb_21_97 bit_21_97 bit_21_98 R_bl
Rbb_21_97 bitb_21_97 bitb_21_98 R_bl
Cb_21_97 bit_21_97 gnd C_bl
Cbb_21_97 bitb_21_97 gnd C_bl
Rb_21_98 bit_21_98 bit_21_99 R_bl
Rbb_21_98 bitb_21_98 bitb_21_99 R_bl
Cb_21_98 bit_21_98 gnd C_bl
Cbb_21_98 bitb_21_98 gnd C_bl
Rb_21_99 bit_21_99 bit_21_100 R_bl
Rbb_21_99 bitb_21_99 bitb_21_100 R_bl
Cb_21_99 bit_21_99 gnd C_bl
Cbb_21_99 bitb_21_99 gnd C_bl
Rb_22_0 bit_22_0 bit_22_1 R_bl
Rbb_22_0 bitb_22_0 bitb_22_1 R_bl
Cb_22_0 bit_22_0 gnd C_bl
Cbb_22_0 bitb_22_0 gnd C_bl
Rb_22_1 bit_22_1 bit_22_2 R_bl
Rbb_22_1 bitb_22_1 bitb_22_2 R_bl
Cb_22_1 bit_22_1 gnd C_bl
Cbb_22_1 bitb_22_1 gnd C_bl
Rb_22_2 bit_22_2 bit_22_3 R_bl
Rbb_22_2 bitb_22_2 bitb_22_3 R_bl
Cb_22_2 bit_22_2 gnd C_bl
Cbb_22_2 bitb_22_2 gnd C_bl
Rb_22_3 bit_22_3 bit_22_4 R_bl
Rbb_22_3 bitb_22_3 bitb_22_4 R_bl
Cb_22_3 bit_22_3 gnd C_bl
Cbb_22_3 bitb_22_3 gnd C_bl
Rb_22_4 bit_22_4 bit_22_5 R_bl
Rbb_22_4 bitb_22_4 bitb_22_5 R_bl
Cb_22_4 bit_22_4 gnd C_bl
Cbb_22_4 bitb_22_4 gnd C_bl
Rb_22_5 bit_22_5 bit_22_6 R_bl
Rbb_22_5 bitb_22_5 bitb_22_6 R_bl
Cb_22_5 bit_22_5 gnd C_bl
Cbb_22_5 bitb_22_5 gnd C_bl
Rb_22_6 bit_22_6 bit_22_7 R_bl
Rbb_22_6 bitb_22_6 bitb_22_7 R_bl
Cb_22_6 bit_22_6 gnd C_bl
Cbb_22_6 bitb_22_6 gnd C_bl
Rb_22_7 bit_22_7 bit_22_8 R_bl
Rbb_22_7 bitb_22_7 bitb_22_8 R_bl
Cb_22_7 bit_22_7 gnd C_bl
Cbb_22_7 bitb_22_7 gnd C_bl
Rb_22_8 bit_22_8 bit_22_9 R_bl
Rbb_22_8 bitb_22_8 bitb_22_9 R_bl
Cb_22_8 bit_22_8 gnd C_bl
Cbb_22_8 bitb_22_8 gnd C_bl
Rb_22_9 bit_22_9 bit_22_10 R_bl
Rbb_22_9 bitb_22_9 bitb_22_10 R_bl
Cb_22_9 bit_22_9 gnd C_bl
Cbb_22_9 bitb_22_9 gnd C_bl
Rb_22_10 bit_22_10 bit_22_11 R_bl
Rbb_22_10 bitb_22_10 bitb_22_11 R_bl
Cb_22_10 bit_22_10 gnd C_bl
Cbb_22_10 bitb_22_10 gnd C_bl
Rb_22_11 bit_22_11 bit_22_12 R_bl
Rbb_22_11 bitb_22_11 bitb_22_12 R_bl
Cb_22_11 bit_22_11 gnd C_bl
Cbb_22_11 bitb_22_11 gnd C_bl
Rb_22_12 bit_22_12 bit_22_13 R_bl
Rbb_22_12 bitb_22_12 bitb_22_13 R_bl
Cb_22_12 bit_22_12 gnd C_bl
Cbb_22_12 bitb_22_12 gnd C_bl
Rb_22_13 bit_22_13 bit_22_14 R_bl
Rbb_22_13 bitb_22_13 bitb_22_14 R_bl
Cb_22_13 bit_22_13 gnd C_bl
Cbb_22_13 bitb_22_13 gnd C_bl
Rb_22_14 bit_22_14 bit_22_15 R_bl
Rbb_22_14 bitb_22_14 bitb_22_15 R_bl
Cb_22_14 bit_22_14 gnd C_bl
Cbb_22_14 bitb_22_14 gnd C_bl
Rb_22_15 bit_22_15 bit_22_16 R_bl
Rbb_22_15 bitb_22_15 bitb_22_16 R_bl
Cb_22_15 bit_22_15 gnd C_bl
Cbb_22_15 bitb_22_15 gnd C_bl
Rb_22_16 bit_22_16 bit_22_17 R_bl
Rbb_22_16 bitb_22_16 bitb_22_17 R_bl
Cb_22_16 bit_22_16 gnd C_bl
Cbb_22_16 bitb_22_16 gnd C_bl
Rb_22_17 bit_22_17 bit_22_18 R_bl
Rbb_22_17 bitb_22_17 bitb_22_18 R_bl
Cb_22_17 bit_22_17 gnd C_bl
Cbb_22_17 bitb_22_17 gnd C_bl
Rb_22_18 bit_22_18 bit_22_19 R_bl
Rbb_22_18 bitb_22_18 bitb_22_19 R_bl
Cb_22_18 bit_22_18 gnd C_bl
Cbb_22_18 bitb_22_18 gnd C_bl
Rb_22_19 bit_22_19 bit_22_20 R_bl
Rbb_22_19 bitb_22_19 bitb_22_20 R_bl
Cb_22_19 bit_22_19 gnd C_bl
Cbb_22_19 bitb_22_19 gnd C_bl
Rb_22_20 bit_22_20 bit_22_21 R_bl
Rbb_22_20 bitb_22_20 bitb_22_21 R_bl
Cb_22_20 bit_22_20 gnd C_bl
Cbb_22_20 bitb_22_20 gnd C_bl
Rb_22_21 bit_22_21 bit_22_22 R_bl
Rbb_22_21 bitb_22_21 bitb_22_22 R_bl
Cb_22_21 bit_22_21 gnd C_bl
Cbb_22_21 bitb_22_21 gnd C_bl
Rb_22_22 bit_22_22 bit_22_23 R_bl
Rbb_22_22 bitb_22_22 bitb_22_23 R_bl
Cb_22_22 bit_22_22 gnd C_bl
Cbb_22_22 bitb_22_22 gnd C_bl
Rb_22_23 bit_22_23 bit_22_24 R_bl
Rbb_22_23 bitb_22_23 bitb_22_24 R_bl
Cb_22_23 bit_22_23 gnd C_bl
Cbb_22_23 bitb_22_23 gnd C_bl
Rb_22_24 bit_22_24 bit_22_25 R_bl
Rbb_22_24 bitb_22_24 bitb_22_25 R_bl
Cb_22_24 bit_22_24 gnd C_bl
Cbb_22_24 bitb_22_24 gnd C_bl
Rb_22_25 bit_22_25 bit_22_26 R_bl
Rbb_22_25 bitb_22_25 bitb_22_26 R_bl
Cb_22_25 bit_22_25 gnd C_bl
Cbb_22_25 bitb_22_25 gnd C_bl
Rb_22_26 bit_22_26 bit_22_27 R_bl
Rbb_22_26 bitb_22_26 bitb_22_27 R_bl
Cb_22_26 bit_22_26 gnd C_bl
Cbb_22_26 bitb_22_26 gnd C_bl
Rb_22_27 bit_22_27 bit_22_28 R_bl
Rbb_22_27 bitb_22_27 bitb_22_28 R_bl
Cb_22_27 bit_22_27 gnd C_bl
Cbb_22_27 bitb_22_27 gnd C_bl
Rb_22_28 bit_22_28 bit_22_29 R_bl
Rbb_22_28 bitb_22_28 bitb_22_29 R_bl
Cb_22_28 bit_22_28 gnd C_bl
Cbb_22_28 bitb_22_28 gnd C_bl
Rb_22_29 bit_22_29 bit_22_30 R_bl
Rbb_22_29 bitb_22_29 bitb_22_30 R_bl
Cb_22_29 bit_22_29 gnd C_bl
Cbb_22_29 bitb_22_29 gnd C_bl
Rb_22_30 bit_22_30 bit_22_31 R_bl
Rbb_22_30 bitb_22_30 bitb_22_31 R_bl
Cb_22_30 bit_22_30 gnd C_bl
Cbb_22_30 bitb_22_30 gnd C_bl
Rb_22_31 bit_22_31 bit_22_32 R_bl
Rbb_22_31 bitb_22_31 bitb_22_32 R_bl
Cb_22_31 bit_22_31 gnd C_bl
Cbb_22_31 bitb_22_31 gnd C_bl
Rb_22_32 bit_22_32 bit_22_33 R_bl
Rbb_22_32 bitb_22_32 bitb_22_33 R_bl
Cb_22_32 bit_22_32 gnd C_bl
Cbb_22_32 bitb_22_32 gnd C_bl
Rb_22_33 bit_22_33 bit_22_34 R_bl
Rbb_22_33 bitb_22_33 bitb_22_34 R_bl
Cb_22_33 bit_22_33 gnd C_bl
Cbb_22_33 bitb_22_33 gnd C_bl
Rb_22_34 bit_22_34 bit_22_35 R_bl
Rbb_22_34 bitb_22_34 bitb_22_35 R_bl
Cb_22_34 bit_22_34 gnd C_bl
Cbb_22_34 bitb_22_34 gnd C_bl
Rb_22_35 bit_22_35 bit_22_36 R_bl
Rbb_22_35 bitb_22_35 bitb_22_36 R_bl
Cb_22_35 bit_22_35 gnd C_bl
Cbb_22_35 bitb_22_35 gnd C_bl
Rb_22_36 bit_22_36 bit_22_37 R_bl
Rbb_22_36 bitb_22_36 bitb_22_37 R_bl
Cb_22_36 bit_22_36 gnd C_bl
Cbb_22_36 bitb_22_36 gnd C_bl
Rb_22_37 bit_22_37 bit_22_38 R_bl
Rbb_22_37 bitb_22_37 bitb_22_38 R_bl
Cb_22_37 bit_22_37 gnd C_bl
Cbb_22_37 bitb_22_37 gnd C_bl
Rb_22_38 bit_22_38 bit_22_39 R_bl
Rbb_22_38 bitb_22_38 bitb_22_39 R_bl
Cb_22_38 bit_22_38 gnd C_bl
Cbb_22_38 bitb_22_38 gnd C_bl
Rb_22_39 bit_22_39 bit_22_40 R_bl
Rbb_22_39 bitb_22_39 bitb_22_40 R_bl
Cb_22_39 bit_22_39 gnd C_bl
Cbb_22_39 bitb_22_39 gnd C_bl
Rb_22_40 bit_22_40 bit_22_41 R_bl
Rbb_22_40 bitb_22_40 bitb_22_41 R_bl
Cb_22_40 bit_22_40 gnd C_bl
Cbb_22_40 bitb_22_40 gnd C_bl
Rb_22_41 bit_22_41 bit_22_42 R_bl
Rbb_22_41 bitb_22_41 bitb_22_42 R_bl
Cb_22_41 bit_22_41 gnd C_bl
Cbb_22_41 bitb_22_41 gnd C_bl
Rb_22_42 bit_22_42 bit_22_43 R_bl
Rbb_22_42 bitb_22_42 bitb_22_43 R_bl
Cb_22_42 bit_22_42 gnd C_bl
Cbb_22_42 bitb_22_42 gnd C_bl
Rb_22_43 bit_22_43 bit_22_44 R_bl
Rbb_22_43 bitb_22_43 bitb_22_44 R_bl
Cb_22_43 bit_22_43 gnd C_bl
Cbb_22_43 bitb_22_43 gnd C_bl
Rb_22_44 bit_22_44 bit_22_45 R_bl
Rbb_22_44 bitb_22_44 bitb_22_45 R_bl
Cb_22_44 bit_22_44 gnd C_bl
Cbb_22_44 bitb_22_44 gnd C_bl
Rb_22_45 bit_22_45 bit_22_46 R_bl
Rbb_22_45 bitb_22_45 bitb_22_46 R_bl
Cb_22_45 bit_22_45 gnd C_bl
Cbb_22_45 bitb_22_45 gnd C_bl
Rb_22_46 bit_22_46 bit_22_47 R_bl
Rbb_22_46 bitb_22_46 bitb_22_47 R_bl
Cb_22_46 bit_22_46 gnd C_bl
Cbb_22_46 bitb_22_46 gnd C_bl
Rb_22_47 bit_22_47 bit_22_48 R_bl
Rbb_22_47 bitb_22_47 bitb_22_48 R_bl
Cb_22_47 bit_22_47 gnd C_bl
Cbb_22_47 bitb_22_47 gnd C_bl
Rb_22_48 bit_22_48 bit_22_49 R_bl
Rbb_22_48 bitb_22_48 bitb_22_49 R_bl
Cb_22_48 bit_22_48 gnd C_bl
Cbb_22_48 bitb_22_48 gnd C_bl
Rb_22_49 bit_22_49 bit_22_50 R_bl
Rbb_22_49 bitb_22_49 bitb_22_50 R_bl
Cb_22_49 bit_22_49 gnd C_bl
Cbb_22_49 bitb_22_49 gnd C_bl
Rb_22_50 bit_22_50 bit_22_51 R_bl
Rbb_22_50 bitb_22_50 bitb_22_51 R_bl
Cb_22_50 bit_22_50 gnd C_bl
Cbb_22_50 bitb_22_50 gnd C_bl
Rb_22_51 bit_22_51 bit_22_52 R_bl
Rbb_22_51 bitb_22_51 bitb_22_52 R_bl
Cb_22_51 bit_22_51 gnd C_bl
Cbb_22_51 bitb_22_51 gnd C_bl
Rb_22_52 bit_22_52 bit_22_53 R_bl
Rbb_22_52 bitb_22_52 bitb_22_53 R_bl
Cb_22_52 bit_22_52 gnd C_bl
Cbb_22_52 bitb_22_52 gnd C_bl
Rb_22_53 bit_22_53 bit_22_54 R_bl
Rbb_22_53 bitb_22_53 bitb_22_54 R_bl
Cb_22_53 bit_22_53 gnd C_bl
Cbb_22_53 bitb_22_53 gnd C_bl
Rb_22_54 bit_22_54 bit_22_55 R_bl
Rbb_22_54 bitb_22_54 bitb_22_55 R_bl
Cb_22_54 bit_22_54 gnd C_bl
Cbb_22_54 bitb_22_54 gnd C_bl
Rb_22_55 bit_22_55 bit_22_56 R_bl
Rbb_22_55 bitb_22_55 bitb_22_56 R_bl
Cb_22_55 bit_22_55 gnd C_bl
Cbb_22_55 bitb_22_55 gnd C_bl
Rb_22_56 bit_22_56 bit_22_57 R_bl
Rbb_22_56 bitb_22_56 bitb_22_57 R_bl
Cb_22_56 bit_22_56 gnd C_bl
Cbb_22_56 bitb_22_56 gnd C_bl
Rb_22_57 bit_22_57 bit_22_58 R_bl
Rbb_22_57 bitb_22_57 bitb_22_58 R_bl
Cb_22_57 bit_22_57 gnd C_bl
Cbb_22_57 bitb_22_57 gnd C_bl
Rb_22_58 bit_22_58 bit_22_59 R_bl
Rbb_22_58 bitb_22_58 bitb_22_59 R_bl
Cb_22_58 bit_22_58 gnd C_bl
Cbb_22_58 bitb_22_58 gnd C_bl
Rb_22_59 bit_22_59 bit_22_60 R_bl
Rbb_22_59 bitb_22_59 bitb_22_60 R_bl
Cb_22_59 bit_22_59 gnd C_bl
Cbb_22_59 bitb_22_59 gnd C_bl
Rb_22_60 bit_22_60 bit_22_61 R_bl
Rbb_22_60 bitb_22_60 bitb_22_61 R_bl
Cb_22_60 bit_22_60 gnd C_bl
Cbb_22_60 bitb_22_60 gnd C_bl
Rb_22_61 bit_22_61 bit_22_62 R_bl
Rbb_22_61 bitb_22_61 bitb_22_62 R_bl
Cb_22_61 bit_22_61 gnd C_bl
Cbb_22_61 bitb_22_61 gnd C_bl
Rb_22_62 bit_22_62 bit_22_63 R_bl
Rbb_22_62 bitb_22_62 bitb_22_63 R_bl
Cb_22_62 bit_22_62 gnd C_bl
Cbb_22_62 bitb_22_62 gnd C_bl
Rb_22_63 bit_22_63 bit_22_64 R_bl
Rbb_22_63 bitb_22_63 bitb_22_64 R_bl
Cb_22_63 bit_22_63 gnd C_bl
Cbb_22_63 bitb_22_63 gnd C_bl
Rb_22_64 bit_22_64 bit_22_65 R_bl
Rbb_22_64 bitb_22_64 bitb_22_65 R_bl
Cb_22_64 bit_22_64 gnd C_bl
Cbb_22_64 bitb_22_64 gnd C_bl
Rb_22_65 bit_22_65 bit_22_66 R_bl
Rbb_22_65 bitb_22_65 bitb_22_66 R_bl
Cb_22_65 bit_22_65 gnd C_bl
Cbb_22_65 bitb_22_65 gnd C_bl
Rb_22_66 bit_22_66 bit_22_67 R_bl
Rbb_22_66 bitb_22_66 bitb_22_67 R_bl
Cb_22_66 bit_22_66 gnd C_bl
Cbb_22_66 bitb_22_66 gnd C_bl
Rb_22_67 bit_22_67 bit_22_68 R_bl
Rbb_22_67 bitb_22_67 bitb_22_68 R_bl
Cb_22_67 bit_22_67 gnd C_bl
Cbb_22_67 bitb_22_67 gnd C_bl
Rb_22_68 bit_22_68 bit_22_69 R_bl
Rbb_22_68 bitb_22_68 bitb_22_69 R_bl
Cb_22_68 bit_22_68 gnd C_bl
Cbb_22_68 bitb_22_68 gnd C_bl
Rb_22_69 bit_22_69 bit_22_70 R_bl
Rbb_22_69 bitb_22_69 bitb_22_70 R_bl
Cb_22_69 bit_22_69 gnd C_bl
Cbb_22_69 bitb_22_69 gnd C_bl
Rb_22_70 bit_22_70 bit_22_71 R_bl
Rbb_22_70 bitb_22_70 bitb_22_71 R_bl
Cb_22_70 bit_22_70 gnd C_bl
Cbb_22_70 bitb_22_70 gnd C_bl
Rb_22_71 bit_22_71 bit_22_72 R_bl
Rbb_22_71 bitb_22_71 bitb_22_72 R_bl
Cb_22_71 bit_22_71 gnd C_bl
Cbb_22_71 bitb_22_71 gnd C_bl
Rb_22_72 bit_22_72 bit_22_73 R_bl
Rbb_22_72 bitb_22_72 bitb_22_73 R_bl
Cb_22_72 bit_22_72 gnd C_bl
Cbb_22_72 bitb_22_72 gnd C_bl
Rb_22_73 bit_22_73 bit_22_74 R_bl
Rbb_22_73 bitb_22_73 bitb_22_74 R_bl
Cb_22_73 bit_22_73 gnd C_bl
Cbb_22_73 bitb_22_73 gnd C_bl
Rb_22_74 bit_22_74 bit_22_75 R_bl
Rbb_22_74 bitb_22_74 bitb_22_75 R_bl
Cb_22_74 bit_22_74 gnd C_bl
Cbb_22_74 bitb_22_74 gnd C_bl
Rb_22_75 bit_22_75 bit_22_76 R_bl
Rbb_22_75 bitb_22_75 bitb_22_76 R_bl
Cb_22_75 bit_22_75 gnd C_bl
Cbb_22_75 bitb_22_75 gnd C_bl
Rb_22_76 bit_22_76 bit_22_77 R_bl
Rbb_22_76 bitb_22_76 bitb_22_77 R_bl
Cb_22_76 bit_22_76 gnd C_bl
Cbb_22_76 bitb_22_76 gnd C_bl
Rb_22_77 bit_22_77 bit_22_78 R_bl
Rbb_22_77 bitb_22_77 bitb_22_78 R_bl
Cb_22_77 bit_22_77 gnd C_bl
Cbb_22_77 bitb_22_77 gnd C_bl
Rb_22_78 bit_22_78 bit_22_79 R_bl
Rbb_22_78 bitb_22_78 bitb_22_79 R_bl
Cb_22_78 bit_22_78 gnd C_bl
Cbb_22_78 bitb_22_78 gnd C_bl
Rb_22_79 bit_22_79 bit_22_80 R_bl
Rbb_22_79 bitb_22_79 bitb_22_80 R_bl
Cb_22_79 bit_22_79 gnd C_bl
Cbb_22_79 bitb_22_79 gnd C_bl
Rb_22_80 bit_22_80 bit_22_81 R_bl
Rbb_22_80 bitb_22_80 bitb_22_81 R_bl
Cb_22_80 bit_22_80 gnd C_bl
Cbb_22_80 bitb_22_80 gnd C_bl
Rb_22_81 bit_22_81 bit_22_82 R_bl
Rbb_22_81 bitb_22_81 bitb_22_82 R_bl
Cb_22_81 bit_22_81 gnd C_bl
Cbb_22_81 bitb_22_81 gnd C_bl
Rb_22_82 bit_22_82 bit_22_83 R_bl
Rbb_22_82 bitb_22_82 bitb_22_83 R_bl
Cb_22_82 bit_22_82 gnd C_bl
Cbb_22_82 bitb_22_82 gnd C_bl
Rb_22_83 bit_22_83 bit_22_84 R_bl
Rbb_22_83 bitb_22_83 bitb_22_84 R_bl
Cb_22_83 bit_22_83 gnd C_bl
Cbb_22_83 bitb_22_83 gnd C_bl
Rb_22_84 bit_22_84 bit_22_85 R_bl
Rbb_22_84 bitb_22_84 bitb_22_85 R_bl
Cb_22_84 bit_22_84 gnd C_bl
Cbb_22_84 bitb_22_84 gnd C_bl
Rb_22_85 bit_22_85 bit_22_86 R_bl
Rbb_22_85 bitb_22_85 bitb_22_86 R_bl
Cb_22_85 bit_22_85 gnd C_bl
Cbb_22_85 bitb_22_85 gnd C_bl
Rb_22_86 bit_22_86 bit_22_87 R_bl
Rbb_22_86 bitb_22_86 bitb_22_87 R_bl
Cb_22_86 bit_22_86 gnd C_bl
Cbb_22_86 bitb_22_86 gnd C_bl
Rb_22_87 bit_22_87 bit_22_88 R_bl
Rbb_22_87 bitb_22_87 bitb_22_88 R_bl
Cb_22_87 bit_22_87 gnd C_bl
Cbb_22_87 bitb_22_87 gnd C_bl
Rb_22_88 bit_22_88 bit_22_89 R_bl
Rbb_22_88 bitb_22_88 bitb_22_89 R_bl
Cb_22_88 bit_22_88 gnd C_bl
Cbb_22_88 bitb_22_88 gnd C_bl
Rb_22_89 bit_22_89 bit_22_90 R_bl
Rbb_22_89 bitb_22_89 bitb_22_90 R_bl
Cb_22_89 bit_22_89 gnd C_bl
Cbb_22_89 bitb_22_89 gnd C_bl
Rb_22_90 bit_22_90 bit_22_91 R_bl
Rbb_22_90 bitb_22_90 bitb_22_91 R_bl
Cb_22_90 bit_22_90 gnd C_bl
Cbb_22_90 bitb_22_90 gnd C_bl
Rb_22_91 bit_22_91 bit_22_92 R_bl
Rbb_22_91 bitb_22_91 bitb_22_92 R_bl
Cb_22_91 bit_22_91 gnd C_bl
Cbb_22_91 bitb_22_91 gnd C_bl
Rb_22_92 bit_22_92 bit_22_93 R_bl
Rbb_22_92 bitb_22_92 bitb_22_93 R_bl
Cb_22_92 bit_22_92 gnd C_bl
Cbb_22_92 bitb_22_92 gnd C_bl
Rb_22_93 bit_22_93 bit_22_94 R_bl
Rbb_22_93 bitb_22_93 bitb_22_94 R_bl
Cb_22_93 bit_22_93 gnd C_bl
Cbb_22_93 bitb_22_93 gnd C_bl
Rb_22_94 bit_22_94 bit_22_95 R_bl
Rbb_22_94 bitb_22_94 bitb_22_95 R_bl
Cb_22_94 bit_22_94 gnd C_bl
Cbb_22_94 bitb_22_94 gnd C_bl
Rb_22_95 bit_22_95 bit_22_96 R_bl
Rbb_22_95 bitb_22_95 bitb_22_96 R_bl
Cb_22_95 bit_22_95 gnd C_bl
Cbb_22_95 bitb_22_95 gnd C_bl
Rb_22_96 bit_22_96 bit_22_97 R_bl
Rbb_22_96 bitb_22_96 bitb_22_97 R_bl
Cb_22_96 bit_22_96 gnd C_bl
Cbb_22_96 bitb_22_96 gnd C_bl
Rb_22_97 bit_22_97 bit_22_98 R_bl
Rbb_22_97 bitb_22_97 bitb_22_98 R_bl
Cb_22_97 bit_22_97 gnd C_bl
Cbb_22_97 bitb_22_97 gnd C_bl
Rb_22_98 bit_22_98 bit_22_99 R_bl
Rbb_22_98 bitb_22_98 bitb_22_99 R_bl
Cb_22_98 bit_22_98 gnd C_bl
Cbb_22_98 bitb_22_98 gnd C_bl
Rb_22_99 bit_22_99 bit_22_100 R_bl
Rbb_22_99 bitb_22_99 bitb_22_100 R_bl
Cb_22_99 bit_22_99 gnd C_bl
Cbb_22_99 bitb_22_99 gnd C_bl
Rb_23_0 bit_23_0 bit_23_1 R_bl
Rbb_23_0 bitb_23_0 bitb_23_1 R_bl
Cb_23_0 bit_23_0 gnd C_bl
Cbb_23_0 bitb_23_0 gnd C_bl
Rb_23_1 bit_23_1 bit_23_2 R_bl
Rbb_23_1 bitb_23_1 bitb_23_2 R_bl
Cb_23_1 bit_23_1 gnd C_bl
Cbb_23_1 bitb_23_1 gnd C_bl
Rb_23_2 bit_23_2 bit_23_3 R_bl
Rbb_23_2 bitb_23_2 bitb_23_3 R_bl
Cb_23_2 bit_23_2 gnd C_bl
Cbb_23_2 bitb_23_2 gnd C_bl
Rb_23_3 bit_23_3 bit_23_4 R_bl
Rbb_23_3 bitb_23_3 bitb_23_4 R_bl
Cb_23_3 bit_23_3 gnd C_bl
Cbb_23_3 bitb_23_3 gnd C_bl
Rb_23_4 bit_23_4 bit_23_5 R_bl
Rbb_23_4 bitb_23_4 bitb_23_5 R_bl
Cb_23_4 bit_23_4 gnd C_bl
Cbb_23_4 bitb_23_4 gnd C_bl
Rb_23_5 bit_23_5 bit_23_6 R_bl
Rbb_23_5 bitb_23_5 bitb_23_6 R_bl
Cb_23_5 bit_23_5 gnd C_bl
Cbb_23_5 bitb_23_5 gnd C_bl
Rb_23_6 bit_23_6 bit_23_7 R_bl
Rbb_23_6 bitb_23_6 bitb_23_7 R_bl
Cb_23_6 bit_23_6 gnd C_bl
Cbb_23_6 bitb_23_6 gnd C_bl
Rb_23_7 bit_23_7 bit_23_8 R_bl
Rbb_23_7 bitb_23_7 bitb_23_8 R_bl
Cb_23_7 bit_23_7 gnd C_bl
Cbb_23_7 bitb_23_7 gnd C_bl
Rb_23_8 bit_23_8 bit_23_9 R_bl
Rbb_23_8 bitb_23_8 bitb_23_9 R_bl
Cb_23_8 bit_23_8 gnd C_bl
Cbb_23_8 bitb_23_8 gnd C_bl
Rb_23_9 bit_23_9 bit_23_10 R_bl
Rbb_23_9 bitb_23_9 bitb_23_10 R_bl
Cb_23_9 bit_23_9 gnd C_bl
Cbb_23_9 bitb_23_9 gnd C_bl
Rb_23_10 bit_23_10 bit_23_11 R_bl
Rbb_23_10 bitb_23_10 bitb_23_11 R_bl
Cb_23_10 bit_23_10 gnd C_bl
Cbb_23_10 bitb_23_10 gnd C_bl
Rb_23_11 bit_23_11 bit_23_12 R_bl
Rbb_23_11 bitb_23_11 bitb_23_12 R_bl
Cb_23_11 bit_23_11 gnd C_bl
Cbb_23_11 bitb_23_11 gnd C_bl
Rb_23_12 bit_23_12 bit_23_13 R_bl
Rbb_23_12 bitb_23_12 bitb_23_13 R_bl
Cb_23_12 bit_23_12 gnd C_bl
Cbb_23_12 bitb_23_12 gnd C_bl
Rb_23_13 bit_23_13 bit_23_14 R_bl
Rbb_23_13 bitb_23_13 bitb_23_14 R_bl
Cb_23_13 bit_23_13 gnd C_bl
Cbb_23_13 bitb_23_13 gnd C_bl
Rb_23_14 bit_23_14 bit_23_15 R_bl
Rbb_23_14 bitb_23_14 bitb_23_15 R_bl
Cb_23_14 bit_23_14 gnd C_bl
Cbb_23_14 bitb_23_14 gnd C_bl
Rb_23_15 bit_23_15 bit_23_16 R_bl
Rbb_23_15 bitb_23_15 bitb_23_16 R_bl
Cb_23_15 bit_23_15 gnd C_bl
Cbb_23_15 bitb_23_15 gnd C_bl
Rb_23_16 bit_23_16 bit_23_17 R_bl
Rbb_23_16 bitb_23_16 bitb_23_17 R_bl
Cb_23_16 bit_23_16 gnd C_bl
Cbb_23_16 bitb_23_16 gnd C_bl
Rb_23_17 bit_23_17 bit_23_18 R_bl
Rbb_23_17 bitb_23_17 bitb_23_18 R_bl
Cb_23_17 bit_23_17 gnd C_bl
Cbb_23_17 bitb_23_17 gnd C_bl
Rb_23_18 bit_23_18 bit_23_19 R_bl
Rbb_23_18 bitb_23_18 bitb_23_19 R_bl
Cb_23_18 bit_23_18 gnd C_bl
Cbb_23_18 bitb_23_18 gnd C_bl
Rb_23_19 bit_23_19 bit_23_20 R_bl
Rbb_23_19 bitb_23_19 bitb_23_20 R_bl
Cb_23_19 bit_23_19 gnd C_bl
Cbb_23_19 bitb_23_19 gnd C_bl
Rb_23_20 bit_23_20 bit_23_21 R_bl
Rbb_23_20 bitb_23_20 bitb_23_21 R_bl
Cb_23_20 bit_23_20 gnd C_bl
Cbb_23_20 bitb_23_20 gnd C_bl
Rb_23_21 bit_23_21 bit_23_22 R_bl
Rbb_23_21 bitb_23_21 bitb_23_22 R_bl
Cb_23_21 bit_23_21 gnd C_bl
Cbb_23_21 bitb_23_21 gnd C_bl
Rb_23_22 bit_23_22 bit_23_23 R_bl
Rbb_23_22 bitb_23_22 bitb_23_23 R_bl
Cb_23_22 bit_23_22 gnd C_bl
Cbb_23_22 bitb_23_22 gnd C_bl
Rb_23_23 bit_23_23 bit_23_24 R_bl
Rbb_23_23 bitb_23_23 bitb_23_24 R_bl
Cb_23_23 bit_23_23 gnd C_bl
Cbb_23_23 bitb_23_23 gnd C_bl
Rb_23_24 bit_23_24 bit_23_25 R_bl
Rbb_23_24 bitb_23_24 bitb_23_25 R_bl
Cb_23_24 bit_23_24 gnd C_bl
Cbb_23_24 bitb_23_24 gnd C_bl
Rb_23_25 bit_23_25 bit_23_26 R_bl
Rbb_23_25 bitb_23_25 bitb_23_26 R_bl
Cb_23_25 bit_23_25 gnd C_bl
Cbb_23_25 bitb_23_25 gnd C_bl
Rb_23_26 bit_23_26 bit_23_27 R_bl
Rbb_23_26 bitb_23_26 bitb_23_27 R_bl
Cb_23_26 bit_23_26 gnd C_bl
Cbb_23_26 bitb_23_26 gnd C_bl
Rb_23_27 bit_23_27 bit_23_28 R_bl
Rbb_23_27 bitb_23_27 bitb_23_28 R_bl
Cb_23_27 bit_23_27 gnd C_bl
Cbb_23_27 bitb_23_27 gnd C_bl
Rb_23_28 bit_23_28 bit_23_29 R_bl
Rbb_23_28 bitb_23_28 bitb_23_29 R_bl
Cb_23_28 bit_23_28 gnd C_bl
Cbb_23_28 bitb_23_28 gnd C_bl
Rb_23_29 bit_23_29 bit_23_30 R_bl
Rbb_23_29 bitb_23_29 bitb_23_30 R_bl
Cb_23_29 bit_23_29 gnd C_bl
Cbb_23_29 bitb_23_29 gnd C_bl
Rb_23_30 bit_23_30 bit_23_31 R_bl
Rbb_23_30 bitb_23_30 bitb_23_31 R_bl
Cb_23_30 bit_23_30 gnd C_bl
Cbb_23_30 bitb_23_30 gnd C_bl
Rb_23_31 bit_23_31 bit_23_32 R_bl
Rbb_23_31 bitb_23_31 bitb_23_32 R_bl
Cb_23_31 bit_23_31 gnd C_bl
Cbb_23_31 bitb_23_31 gnd C_bl
Rb_23_32 bit_23_32 bit_23_33 R_bl
Rbb_23_32 bitb_23_32 bitb_23_33 R_bl
Cb_23_32 bit_23_32 gnd C_bl
Cbb_23_32 bitb_23_32 gnd C_bl
Rb_23_33 bit_23_33 bit_23_34 R_bl
Rbb_23_33 bitb_23_33 bitb_23_34 R_bl
Cb_23_33 bit_23_33 gnd C_bl
Cbb_23_33 bitb_23_33 gnd C_bl
Rb_23_34 bit_23_34 bit_23_35 R_bl
Rbb_23_34 bitb_23_34 bitb_23_35 R_bl
Cb_23_34 bit_23_34 gnd C_bl
Cbb_23_34 bitb_23_34 gnd C_bl
Rb_23_35 bit_23_35 bit_23_36 R_bl
Rbb_23_35 bitb_23_35 bitb_23_36 R_bl
Cb_23_35 bit_23_35 gnd C_bl
Cbb_23_35 bitb_23_35 gnd C_bl
Rb_23_36 bit_23_36 bit_23_37 R_bl
Rbb_23_36 bitb_23_36 bitb_23_37 R_bl
Cb_23_36 bit_23_36 gnd C_bl
Cbb_23_36 bitb_23_36 gnd C_bl
Rb_23_37 bit_23_37 bit_23_38 R_bl
Rbb_23_37 bitb_23_37 bitb_23_38 R_bl
Cb_23_37 bit_23_37 gnd C_bl
Cbb_23_37 bitb_23_37 gnd C_bl
Rb_23_38 bit_23_38 bit_23_39 R_bl
Rbb_23_38 bitb_23_38 bitb_23_39 R_bl
Cb_23_38 bit_23_38 gnd C_bl
Cbb_23_38 bitb_23_38 gnd C_bl
Rb_23_39 bit_23_39 bit_23_40 R_bl
Rbb_23_39 bitb_23_39 bitb_23_40 R_bl
Cb_23_39 bit_23_39 gnd C_bl
Cbb_23_39 bitb_23_39 gnd C_bl
Rb_23_40 bit_23_40 bit_23_41 R_bl
Rbb_23_40 bitb_23_40 bitb_23_41 R_bl
Cb_23_40 bit_23_40 gnd C_bl
Cbb_23_40 bitb_23_40 gnd C_bl
Rb_23_41 bit_23_41 bit_23_42 R_bl
Rbb_23_41 bitb_23_41 bitb_23_42 R_bl
Cb_23_41 bit_23_41 gnd C_bl
Cbb_23_41 bitb_23_41 gnd C_bl
Rb_23_42 bit_23_42 bit_23_43 R_bl
Rbb_23_42 bitb_23_42 bitb_23_43 R_bl
Cb_23_42 bit_23_42 gnd C_bl
Cbb_23_42 bitb_23_42 gnd C_bl
Rb_23_43 bit_23_43 bit_23_44 R_bl
Rbb_23_43 bitb_23_43 bitb_23_44 R_bl
Cb_23_43 bit_23_43 gnd C_bl
Cbb_23_43 bitb_23_43 gnd C_bl
Rb_23_44 bit_23_44 bit_23_45 R_bl
Rbb_23_44 bitb_23_44 bitb_23_45 R_bl
Cb_23_44 bit_23_44 gnd C_bl
Cbb_23_44 bitb_23_44 gnd C_bl
Rb_23_45 bit_23_45 bit_23_46 R_bl
Rbb_23_45 bitb_23_45 bitb_23_46 R_bl
Cb_23_45 bit_23_45 gnd C_bl
Cbb_23_45 bitb_23_45 gnd C_bl
Rb_23_46 bit_23_46 bit_23_47 R_bl
Rbb_23_46 bitb_23_46 bitb_23_47 R_bl
Cb_23_46 bit_23_46 gnd C_bl
Cbb_23_46 bitb_23_46 gnd C_bl
Rb_23_47 bit_23_47 bit_23_48 R_bl
Rbb_23_47 bitb_23_47 bitb_23_48 R_bl
Cb_23_47 bit_23_47 gnd C_bl
Cbb_23_47 bitb_23_47 gnd C_bl
Rb_23_48 bit_23_48 bit_23_49 R_bl
Rbb_23_48 bitb_23_48 bitb_23_49 R_bl
Cb_23_48 bit_23_48 gnd C_bl
Cbb_23_48 bitb_23_48 gnd C_bl
Rb_23_49 bit_23_49 bit_23_50 R_bl
Rbb_23_49 bitb_23_49 bitb_23_50 R_bl
Cb_23_49 bit_23_49 gnd C_bl
Cbb_23_49 bitb_23_49 gnd C_bl
Rb_23_50 bit_23_50 bit_23_51 R_bl
Rbb_23_50 bitb_23_50 bitb_23_51 R_bl
Cb_23_50 bit_23_50 gnd C_bl
Cbb_23_50 bitb_23_50 gnd C_bl
Rb_23_51 bit_23_51 bit_23_52 R_bl
Rbb_23_51 bitb_23_51 bitb_23_52 R_bl
Cb_23_51 bit_23_51 gnd C_bl
Cbb_23_51 bitb_23_51 gnd C_bl
Rb_23_52 bit_23_52 bit_23_53 R_bl
Rbb_23_52 bitb_23_52 bitb_23_53 R_bl
Cb_23_52 bit_23_52 gnd C_bl
Cbb_23_52 bitb_23_52 gnd C_bl
Rb_23_53 bit_23_53 bit_23_54 R_bl
Rbb_23_53 bitb_23_53 bitb_23_54 R_bl
Cb_23_53 bit_23_53 gnd C_bl
Cbb_23_53 bitb_23_53 gnd C_bl
Rb_23_54 bit_23_54 bit_23_55 R_bl
Rbb_23_54 bitb_23_54 bitb_23_55 R_bl
Cb_23_54 bit_23_54 gnd C_bl
Cbb_23_54 bitb_23_54 gnd C_bl
Rb_23_55 bit_23_55 bit_23_56 R_bl
Rbb_23_55 bitb_23_55 bitb_23_56 R_bl
Cb_23_55 bit_23_55 gnd C_bl
Cbb_23_55 bitb_23_55 gnd C_bl
Rb_23_56 bit_23_56 bit_23_57 R_bl
Rbb_23_56 bitb_23_56 bitb_23_57 R_bl
Cb_23_56 bit_23_56 gnd C_bl
Cbb_23_56 bitb_23_56 gnd C_bl
Rb_23_57 bit_23_57 bit_23_58 R_bl
Rbb_23_57 bitb_23_57 bitb_23_58 R_bl
Cb_23_57 bit_23_57 gnd C_bl
Cbb_23_57 bitb_23_57 gnd C_bl
Rb_23_58 bit_23_58 bit_23_59 R_bl
Rbb_23_58 bitb_23_58 bitb_23_59 R_bl
Cb_23_58 bit_23_58 gnd C_bl
Cbb_23_58 bitb_23_58 gnd C_bl
Rb_23_59 bit_23_59 bit_23_60 R_bl
Rbb_23_59 bitb_23_59 bitb_23_60 R_bl
Cb_23_59 bit_23_59 gnd C_bl
Cbb_23_59 bitb_23_59 gnd C_bl
Rb_23_60 bit_23_60 bit_23_61 R_bl
Rbb_23_60 bitb_23_60 bitb_23_61 R_bl
Cb_23_60 bit_23_60 gnd C_bl
Cbb_23_60 bitb_23_60 gnd C_bl
Rb_23_61 bit_23_61 bit_23_62 R_bl
Rbb_23_61 bitb_23_61 bitb_23_62 R_bl
Cb_23_61 bit_23_61 gnd C_bl
Cbb_23_61 bitb_23_61 gnd C_bl
Rb_23_62 bit_23_62 bit_23_63 R_bl
Rbb_23_62 bitb_23_62 bitb_23_63 R_bl
Cb_23_62 bit_23_62 gnd C_bl
Cbb_23_62 bitb_23_62 gnd C_bl
Rb_23_63 bit_23_63 bit_23_64 R_bl
Rbb_23_63 bitb_23_63 bitb_23_64 R_bl
Cb_23_63 bit_23_63 gnd C_bl
Cbb_23_63 bitb_23_63 gnd C_bl
Rb_23_64 bit_23_64 bit_23_65 R_bl
Rbb_23_64 bitb_23_64 bitb_23_65 R_bl
Cb_23_64 bit_23_64 gnd C_bl
Cbb_23_64 bitb_23_64 gnd C_bl
Rb_23_65 bit_23_65 bit_23_66 R_bl
Rbb_23_65 bitb_23_65 bitb_23_66 R_bl
Cb_23_65 bit_23_65 gnd C_bl
Cbb_23_65 bitb_23_65 gnd C_bl
Rb_23_66 bit_23_66 bit_23_67 R_bl
Rbb_23_66 bitb_23_66 bitb_23_67 R_bl
Cb_23_66 bit_23_66 gnd C_bl
Cbb_23_66 bitb_23_66 gnd C_bl
Rb_23_67 bit_23_67 bit_23_68 R_bl
Rbb_23_67 bitb_23_67 bitb_23_68 R_bl
Cb_23_67 bit_23_67 gnd C_bl
Cbb_23_67 bitb_23_67 gnd C_bl
Rb_23_68 bit_23_68 bit_23_69 R_bl
Rbb_23_68 bitb_23_68 bitb_23_69 R_bl
Cb_23_68 bit_23_68 gnd C_bl
Cbb_23_68 bitb_23_68 gnd C_bl
Rb_23_69 bit_23_69 bit_23_70 R_bl
Rbb_23_69 bitb_23_69 bitb_23_70 R_bl
Cb_23_69 bit_23_69 gnd C_bl
Cbb_23_69 bitb_23_69 gnd C_bl
Rb_23_70 bit_23_70 bit_23_71 R_bl
Rbb_23_70 bitb_23_70 bitb_23_71 R_bl
Cb_23_70 bit_23_70 gnd C_bl
Cbb_23_70 bitb_23_70 gnd C_bl
Rb_23_71 bit_23_71 bit_23_72 R_bl
Rbb_23_71 bitb_23_71 bitb_23_72 R_bl
Cb_23_71 bit_23_71 gnd C_bl
Cbb_23_71 bitb_23_71 gnd C_bl
Rb_23_72 bit_23_72 bit_23_73 R_bl
Rbb_23_72 bitb_23_72 bitb_23_73 R_bl
Cb_23_72 bit_23_72 gnd C_bl
Cbb_23_72 bitb_23_72 gnd C_bl
Rb_23_73 bit_23_73 bit_23_74 R_bl
Rbb_23_73 bitb_23_73 bitb_23_74 R_bl
Cb_23_73 bit_23_73 gnd C_bl
Cbb_23_73 bitb_23_73 gnd C_bl
Rb_23_74 bit_23_74 bit_23_75 R_bl
Rbb_23_74 bitb_23_74 bitb_23_75 R_bl
Cb_23_74 bit_23_74 gnd C_bl
Cbb_23_74 bitb_23_74 gnd C_bl
Rb_23_75 bit_23_75 bit_23_76 R_bl
Rbb_23_75 bitb_23_75 bitb_23_76 R_bl
Cb_23_75 bit_23_75 gnd C_bl
Cbb_23_75 bitb_23_75 gnd C_bl
Rb_23_76 bit_23_76 bit_23_77 R_bl
Rbb_23_76 bitb_23_76 bitb_23_77 R_bl
Cb_23_76 bit_23_76 gnd C_bl
Cbb_23_76 bitb_23_76 gnd C_bl
Rb_23_77 bit_23_77 bit_23_78 R_bl
Rbb_23_77 bitb_23_77 bitb_23_78 R_bl
Cb_23_77 bit_23_77 gnd C_bl
Cbb_23_77 bitb_23_77 gnd C_bl
Rb_23_78 bit_23_78 bit_23_79 R_bl
Rbb_23_78 bitb_23_78 bitb_23_79 R_bl
Cb_23_78 bit_23_78 gnd C_bl
Cbb_23_78 bitb_23_78 gnd C_bl
Rb_23_79 bit_23_79 bit_23_80 R_bl
Rbb_23_79 bitb_23_79 bitb_23_80 R_bl
Cb_23_79 bit_23_79 gnd C_bl
Cbb_23_79 bitb_23_79 gnd C_bl
Rb_23_80 bit_23_80 bit_23_81 R_bl
Rbb_23_80 bitb_23_80 bitb_23_81 R_bl
Cb_23_80 bit_23_80 gnd C_bl
Cbb_23_80 bitb_23_80 gnd C_bl
Rb_23_81 bit_23_81 bit_23_82 R_bl
Rbb_23_81 bitb_23_81 bitb_23_82 R_bl
Cb_23_81 bit_23_81 gnd C_bl
Cbb_23_81 bitb_23_81 gnd C_bl
Rb_23_82 bit_23_82 bit_23_83 R_bl
Rbb_23_82 bitb_23_82 bitb_23_83 R_bl
Cb_23_82 bit_23_82 gnd C_bl
Cbb_23_82 bitb_23_82 gnd C_bl
Rb_23_83 bit_23_83 bit_23_84 R_bl
Rbb_23_83 bitb_23_83 bitb_23_84 R_bl
Cb_23_83 bit_23_83 gnd C_bl
Cbb_23_83 bitb_23_83 gnd C_bl
Rb_23_84 bit_23_84 bit_23_85 R_bl
Rbb_23_84 bitb_23_84 bitb_23_85 R_bl
Cb_23_84 bit_23_84 gnd C_bl
Cbb_23_84 bitb_23_84 gnd C_bl
Rb_23_85 bit_23_85 bit_23_86 R_bl
Rbb_23_85 bitb_23_85 bitb_23_86 R_bl
Cb_23_85 bit_23_85 gnd C_bl
Cbb_23_85 bitb_23_85 gnd C_bl
Rb_23_86 bit_23_86 bit_23_87 R_bl
Rbb_23_86 bitb_23_86 bitb_23_87 R_bl
Cb_23_86 bit_23_86 gnd C_bl
Cbb_23_86 bitb_23_86 gnd C_bl
Rb_23_87 bit_23_87 bit_23_88 R_bl
Rbb_23_87 bitb_23_87 bitb_23_88 R_bl
Cb_23_87 bit_23_87 gnd C_bl
Cbb_23_87 bitb_23_87 gnd C_bl
Rb_23_88 bit_23_88 bit_23_89 R_bl
Rbb_23_88 bitb_23_88 bitb_23_89 R_bl
Cb_23_88 bit_23_88 gnd C_bl
Cbb_23_88 bitb_23_88 gnd C_bl
Rb_23_89 bit_23_89 bit_23_90 R_bl
Rbb_23_89 bitb_23_89 bitb_23_90 R_bl
Cb_23_89 bit_23_89 gnd C_bl
Cbb_23_89 bitb_23_89 gnd C_bl
Rb_23_90 bit_23_90 bit_23_91 R_bl
Rbb_23_90 bitb_23_90 bitb_23_91 R_bl
Cb_23_90 bit_23_90 gnd C_bl
Cbb_23_90 bitb_23_90 gnd C_bl
Rb_23_91 bit_23_91 bit_23_92 R_bl
Rbb_23_91 bitb_23_91 bitb_23_92 R_bl
Cb_23_91 bit_23_91 gnd C_bl
Cbb_23_91 bitb_23_91 gnd C_bl
Rb_23_92 bit_23_92 bit_23_93 R_bl
Rbb_23_92 bitb_23_92 bitb_23_93 R_bl
Cb_23_92 bit_23_92 gnd C_bl
Cbb_23_92 bitb_23_92 gnd C_bl
Rb_23_93 bit_23_93 bit_23_94 R_bl
Rbb_23_93 bitb_23_93 bitb_23_94 R_bl
Cb_23_93 bit_23_93 gnd C_bl
Cbb_23_93 bitb_23_93 gnd C_bl
Rb_23_94 bit_23_94 bit_23_95 R_bl
Rbb_23_94 bitb_23_94 bitb_23_95 R_bl
Cb_23_94 bit_23_94 gnd C_bl
Cbb_23_94 bitb_23_94 gnd C_bl
Rb_23_95 bit_23_95 bit_23_96 R_bl
Rbb_23_95 bitb_23_95 bitb_23_96 R_bl
Cb_23_95 bit_23_95 gnd C_bl
Cbb_23_95 bitb_23_95 gnd C_bl
Rb_23_96 bit_23_96 bit_23_97 R_bl
Rbb_23_96 bitb_23_96 bitb_23_97 R_bl
Cb_23_96 bit_23_96 gnd C_bl
Cbb_23_96 bitb_23_96 gnd C_bl
Rb_23_97 bit_23_97 bit_23_98 R_bl
Rbb_23_97 bitb_23_97 bitb_23_98 R_bl
Cb_23_97 bit_23_97 gnd C_bl
Cbb_23_97 bitb_23_97 gnd C_bl
Rb_23_98 bit_23_98 bit_23_99 R_bl
Rbb_23_98 bitb_23_98 bitb_23_99 R_bl
Cb_23_98 bit_23_98 gnd C_bl
Cbb_23_98 bitb_23_98 gnd C_bl
Rb_23_99 bit_23_99 bit_23_100 R_bl
Rbb_23_99 bitb_23_99 bitb_23_100 R_bl
Cb_23_99 bit_23_99 gnd C_bl
Cbb_23_99 bitb_23_99 gnd C_bl
Rb_24_0 bit_24_0 bit_24_1 R_bl
Rbb_24_0 bitb_24_0 bitb_24_1 R_bl
Cb_24_0 bit_24_0 gnd C_bl
Cbb_24_0 bitb_24_0 gnd C_bl
Rb_24_1 bit_24_1 bit_24_2 R_bl
Rbb_24_1 bitb_24_1 bitb_24_2 R_bl
Cb_24_1 bit_24_1 gnd C_bl
Cbb_24_1 bitb_24_1 gnd C_bl
Rb_24_2 bit_24_2 bit_24_3 R_bl
Rbb_24_2 bitb_24_2 bitb_24_3 R_bl
Cb_24_2 bit_24_2 gnd C_bl
Cbb_24_2 bitb_24_2 gnd C_bl
Rb_24_3 bit_24_3 bit_24_4 R_bl
Rbb_24_3 bitb_24_3 bitb_24_4 R_bl
Cb_24_3 bit_24_3 gnd C_bl
Cbb_24_3 bitb_24_3 gnd C_bl
Rb_24_4 bit_24_4 bit_24_5 R_bl
Rbb_24_4 bitb_24_4 bitb_24_5 R_bl
Cb_24_4 bit_24_4 gnd C_bl
Cbb_24_4 bitb_24_4 gnd C_bl
Rb_24_5 bit_24_5 bit_24_6 R_bl
Rbb_24_5 bitb_24_5 bitb_24_6 R_bl
Cb_24_5 bit_24_5 gnd C_bl
Cbb_24_5 bitb_24_5 gnd C_bl
Rb_24_6 bit_24_6 bit_24_7 R_bl
Rbb_24_6 bitb_24_6 bitb_24_7 R_bl
Cb_24_6 bit_24_6 gnd C_bl
Cbb_24_6 bitb_24_6 gnd C_bl
Rb_24_7 bit_24_7 bit_24_8 R_bl
Rbb_24_7 bitb_24_7 bitb_24_8 R_bl
Cb_24_7 bit_24_7 gnd C_bl
Cbb_24_7 bitb_24_7 gnd C_bl
Rb_24_8 bit_24_8 bit_24_9 R_bl
Rbb_24_8 bitb_24_8 bitb_24_9 R_bl
Cb_24_8 bit_24_8 gnd C_bl
Cbb_24_8 bitb_24_8 gnd C_bl
Rb_24_9 bit_24_9 bit_24_10 R_bl
Rbb_24_9 bitb_24_9 bitb_24_10 R_bl
Cb_24_9 bit_24_9 gnd C_bl
Cbb_24_9 bitb_24_9 gnd C_bl
Rb_24_10 bit_24_10 bit_24_11 R_bl
Rbb_24_10 bitb_24_10 bitb_24_11 R_bl
Cb_24_10 bit_24_10 gnd C_bl
Cbb_24_10 bitb_24_10 gnd C_bl
Rb_24_11 bit_24_11 bit_24_12 R_bl
Rbb_24_11 bitb_24_11 bitb_24_12 R_bl
Cb_24_11 bit_24_11 gnd C_bl
Cbb_24_11 bitb_24_11 gnd C_bl
Rb_24_12 bit_24_12 bit_24_13 R_bl
Rbb_24_12 bitb_24_12 bitb_24_13 R_bl
Cb_24_12 bit_24_12 gnd C_bl
Cbb_24_12 bitb_24_12 gnd C_bl
Rb_24_13 bit_24_13 bit_24_14 R_bl
Rbb_24_13 bitb_24_13 bitb_24_14 R_bl
Cb_24_13 bit_24_13 gnd C_bl
Cbb_24_13 bitb_24_13 gnd C_bl
Rb_24_14 bit_24_14 bit_24_15 R_bl
Rbb_24_14 bitb_24_14 bitb_24_15 R_bl
Cb_24_14 bit_24_14 gnd C_bl
Cbb_24_14 bitb_24_14 gnd C_bl
Rb_24_15 bit_24_15 bit_24_16 R_bl
Rbb_24_15 bitb_24_15 bitb_24_16 R_bl
Cb_24_15 bit_24_15 gnd C_bl
Cbb_24_15 bitb_24_15 gnd C_bl
Rb_24_16 bit_24_16 bit_24_17 R_bl
Rbb_24_16 bitb_24_16 bitb_24_17 R_bl
Cb_24_16 bit_24_16 gnd C_bl
Cbb_24_16 bitb_24_16 gnd C_bl
Rb_24_17 bit_24_17 bit_24_18 R_bl
Rbb_24_17 bitb_24_17 bitb_24_18 R_bl
Cb_24_17 bit_24_17 gnd C_bl
Cbb_24_17 bitb_24_17 gnd C_bl
Rb_24_18 bit_24_18 bit_24_19 R_bl
Rbb_24_18 bitb_24_18 bitb_24_19 R_bl
Cb_24_18 bit_24_18 gnd C_bl
Cbb_24_18 bitb_24_18 gnd C_bl
Rb_24_19 bit_24_19 bit_24_20 R_bl
Rbb_24_19 bitb_24_19 bitb_24_20 R_bl
Cb_24_19 bit_24_19 gnd C_bl
Cbb_24_19 bitb_24_19 gnd C_bl
Rb_24_20 bit_24_20 bit_24_21 R_bl
Rbb_24_20 bitb_24_20 bitb_24_21 R_bl
Cb_24_20 bit_24_20 gnd C_bl
Cbb_24_20 bitb_24_20 gnd C_bl
Rb_24_21 bit_24_21 bit_24_22 R_bl
Rbb_24_21 bitb_24_21 bitb_24_22 R_bl
Cb_24_21 bit_24_21 gnd C_bl
Cbb_24_21 bitb_24_21 gnd C_bl
Rb_24_22 bit_24_22 bit_24_23 R_bl
Rbb_24_22 bitb_24_22 bitb_24_23 R_bl
Cb_24_22 bit_24_22 gnd C_bl
Cbb_24_22 bitb_24_22 gnd C_bl
Rb_24_23 bit_24_23 bit_24_24 R_bl
Rbb_24_23 bitb_24_23 bitb_24_24 R_bl
Cb_24_23 bit_24_23 gnd C_bl
Cbb_24_23 bitb_24_23 gnd C_bl
Rb_24_24 bit_24_24 bit_24_25 R_bl
Rbb_24_24 bitb_24_24 bitb_24_25 R_bl
Cb_24_24 bit_24_24 gnd C_bl
Cbb_24_24 bitb_24_24 gnd C_bl
Rb_24_25 bit_24_25 bit_24_26 R_bl
Rbb_24_25 bitb_24_25 bitb_24_26 R_bl
Cb_24_25 bit_24_25 gnd C_bl
Cbb_24_25 bitb_24_25 gnd C_bl
Rb_24_26 bit_24_26 bit_24_27 R_bl
Rbb_24_26 bitb_24_26 bitb_24_27 R_bl
Cb_24_26 bit_24_26 gnd C_bl
Cbb_24_26 bitb_24_26 gnd C_bl
Rb_24_27 bit_24_27 bit_24_28 R_bl
Rbb_24_27 bitb_24_27 bitb_24_28 R_bl
Cb_24_27 bit_24_27 gnd C_bl
Cbb_24_27 bitb_24_27 gnd C_bl
Rb_24_28 bit_24_28 bit_24_29 R_bl
Rbb_24_28 bitb_24_28 bitb_24_29 R_bl
Cb_24_28 bit_24_28 gnd C_bl
Cbb_24_28 bitb_24_28 gnd C_bl
Rb_24_29 bit_24_29 bit_24_30 R_bl
Rbb_24_29 bitb_24_29 bitb_24_30 R_bl
Cb_24_29 bit_24_29 gnd C_bl
Cbb_24_29 bitb_24_29 gnd C_bl
Rb_24_30 bit_24_30 bit_24_31 R_bl
Rbb_24_30 bitb_24_30 bitb_24_31 R_bl
Cb_24_30 bit_24_30 gnd C_bl
Cbb_24_30 bitb_24_30 gnd C_bl
Rb_24_31 bit_24_31 bit_24_32 R_bl
Rbb_24_31 bitb_24_31 bitb_24_32 R_bl
Cb_24_31 bit_24_31 gnd C_bl
Cbb_24_31 bitb_24_31 gnd C_bl
Rb_24_32 bit_24_32 bit_24_33 R_bl
Rbb_24_32 bitb_24_32 bitb_24_33 R_bl
Cb_24_32 bit_24_32 gnd C_bl
Cbb_24_32 bitb_24_32 gnd C_bl
Rb_24_33 bit_24_33 bit_24_34 R_bl
Rbb_24_33 bitb_24_33 bitb_24_34 R_bl
Cb_24_33 bit_24_33 gnd C_bl
Cbb_24_33 bitb_24_33 gnd C_bl
Rb_24_34 bit_24_34 bit_24_35 R_bl
Rbb_24_34 bitb_24_34 bitb_24_35 R_bl
Cb_24_34 bit_24_34 gnd C_bl
Cbb_24_34 bitb_24_34 gnd C_bl
Rb_24_35 bit_24_35 bit_24_36 R_bl
Rbb_24_35 bitb_24_35 bitb_24_36 R_bl
Cb_24_35 bit_24_35 gnd C_bl
Cbb_24_35 bitb_24_35 gnd C_bl
Rb_24_36 bit_24_36 bit_24_37 R_bl
Rbb_24_36 bitb_24_36 bitb_24_37 R_bl
Cb_24_36 bit_24_36 gnd C_bl
Cbb_24_36 bitb_24_36 gnd C_bl
Rb_24_37 bit_24_37 bit_24_38 R_bl
Rbb_24_37 bitb_24_37 bitb_24_38 R_bl
Cb_24_37 bit_24_37 gnd C_bl
Cbb_24_37 bitb_24_37 gnd C_bl
Rb_24_38 bit_24_38 bit_24_39 R_bl
Rbb_24_38 bitb_24_38 bitb_24_39 R_bl
Cb_24_38 bit_24_38 gnd C_bl
Cbb_24_38 bitb_24_38 gnd C_bl
Rb_24_39 bit_24_39 bit_24_40 R_bl
Rbb_24_39 bitb_24_39 bitb_24_40 R_bl
Cb_24_39 bit_24_39 gnd C_bl
Cbb_24_39 bitb_24_39 gnd C_bl
Rb_24_40 bit_24_40 bit_24_41 R_bl
Rbb_24_40 bitb_24_40 bitb_24_41 R_bl
Cb_24_40 bit_24_40 gnd C_bl
Cbb_24_40 bitb_24_40 gnd C_bl
Rb_24_41 bit_24_41 bit_24_42 R_bl
Rbb_24_41 bitb_24_41 bitb_24_42 R_bl
Cb_24_41 bit_24_41 gnd C_bl
Cbb_24_41 bitb_24_41 gnd C_bl
Rb_24_42 bit_24_42 bit_24_43 R_bl
Rbb_24_42 bitb_24_42 bitb_24_43 R_bl
Cb_24_42 bit_24_42 gnd C_bl
Cbb_24_42 bitb_24_42 gnd C_bl
Rb_24_43 bit_24_43 bit_24_44 R_bl
Rbb_24_43 bitb_24_43 bitb_24_44 R_bl
Cb_24_43 bit_24_43 gnd C_bl
Cbb_24_43 bitb_24_43 gnd C_bl
Rb_24_44 bit_24_44 bit_24_45 R_bl
Rbb_24_44 bitb_24_44 bitb_24_45 R_bl
Cb_24_44 bit_24_44 gnd C_bl
Cbb_24_44 bitb_24_44 gnd C_bl
Rb_24_45 bit_24_45 bit_24_46 R_bl
Rbb_24_45 bitb_24_45 bitb_24_46 R_bl
Cb_24_45 bit_24_45 gnd C_bl
Cbb_24_45 bitb_24_45 gnd C_bl
Rb_24_46 bit_24_46 bit_24_47 R_bl
Rbb_24_46 bitb_24_46 bitb_24_47 R_bl
Cb_24_46 bit_24_46 gnd C_bl
Cbb_24_46 bitb_24_46 gnd C_bl
Rb_24_47 bit_24_47 bit_24_48 R_bl
Rbb_24_47 bitb_24_47 bitb_24_48 R_bl
Cb_24_47 bit_24_47 gnd C_bl
Cbb_24_47 bitb_24_47 gnd C_bl
Rb_24_48 bit_24_48 bit_24_49 R_bl
Rbb_24_48 bitb_24_48 bitb_24_49 R_bl
Cb_24_48 bit_24_48 gnd C_bl
Cbb_24_48 bitb_24_48 gnd C_bl
Rb_24_49 bit_24_49 bit_24_50 R_bl
Rbb_24_49 bitb_24_49 bitb_24_50 R_bl
Cb_24_49 bit_24_49 gnd C_bl
Cbb_24_49 bitb_24_49 gnd C_bl
Rb_24_50 bit_24_50 bit_24_51 R_bl
Rbb_24_50 bitb_24_50 bitb_24_51 R_bl
Cb_24_50 bit_24_50 gnd C_bl
Cbb_24_50 bitb_24_50 gnd C_bl
Rb_24_51 bit_24_51 bit_24_52 R_bl
Rbb_24_51 bitb_24_51 bitb_24_52 R_bl
Cb_24_51 bit_24_51 gnd C_bl
Cbb_24_51 bitb_24_51 gnd C_bl
Rb_24_52 bit_24_52 bit_24_53 R_bl
Rbb_24_52 bitb_24_52 bitb_24_53 R_bl
Cb_24_52 bit_24_52 gnd C_bl
Cbb_24_52 bitb_24_52 gnd C_bl
Rb_24_53 bit_24_53 bit_24_54 R_bl
Rbb_24_53 bitb_24_53 bitb_24_54 R_bl
Cb_24_53 bit_24_53 gnd C_bl
Cbb_24_53 bitb_24_53 gnd C_bl
Rb_24_54 bit_24_54 bit_24_55 R_bl
Rbb_24_54 bitb_24_54 bitb_24_55 R_bl
Cb_24_54 bit_24_54 gnd C_bl
Cbb_24_54 bitb_24_54 gnd C_bl
Rb_24_55 bit_24_55 bit_24_56 R_bl
Rbb_24_55 bitb_24_55 bitb_24_56 R_bl
Cb_24_55 bit_24_55 gnd C_bl
Cbb_24_55 bitb_24_55 gnd C_bl
Rb_24_56 bit_24_56 bit_24_57 R_bl
Rbb_24_56 bitb_24_56 bitb_24_57 R_bl
Cb_24_56 bit_24_56 gnd C_bl
Cbb_24_56 bitb_24_56 gnd C_bl
Rb_24_57 bit_24_57 bit_24_58 R_bl
Rbb_24_57 bitb_24_57 bitb_24_58 R_bl
Cb_24_57 bit_24_57 gnd C_bl
Cbb_24_57 bitb_24_57 gnd C_bl
Rb_24_58 bit_24_58 bit_24_59 R_bl
Rbb_24_58 bitb_24_58 bitb_24_59 R_bl
Cb_24_58 bit_24_58 gnd C_bl
Cbb_24_58 bitb_24_58 gnd C_bl
Rb_24_59 bit_24_59 bit_24_60 R_bl
Rbb_24_59 bitb_24_59 bitb_24_60 R_bl
Cb_24_59 bit_24_59 gnd C_bl
Cbb_24_59 bitb_24_59 gnd C_bl
Rb_24_60 bit_24_60 bit_24_61 R_bl
Rbb_24_60 bitb_24_60 bitb_24_61 R_bl
Cb_24_60 bit_24_60 gnd C_bl
Cbb_24_60 bitb_24_60 gnd C_bl
Rb_24_61 bit_24_61 bit_24_62 R_bl
Rbb_24_61 bitb_24_61 bitb_24_62 R_bl
Cb_24_61 bit_24_61 gnd C_bl
Cbb_24_61 bitb_24_61 gnd C_bl
Rb_24_62 bit_24_62 bit_24_63 R_bl
Rbb_24_62 bitb_24_62 bitb_24_63 R_bl
Cb_24_62 bit_24_62 gnd C_bl
Cbb_24_62 bitb_24_62 gnd C_bl
Rb_24_63 bit_24_63 bit_24_64 R_bl
Rbb_24_63 bitb_24_63 bitb_24_64 R_bl
Cb_24_63 bit_24_63 gnd C_bl
Cbb_24_63 bitb_24_63 gnd C_bl
Rb_24_64 bit_24_64 bit_24_65 R_bl
Rbb_24_64 bitb_24_64 bitb_24_65 R_bl
Cb_24_64 bit_24_64 gnd C_bl
Cbb_24_64 bitb_24_64 gnd C_bl
Rb_24_65 bit_24_65 bit_24_66 R_bl
Rbb_24_65 bitb_24_65 bitb_24_66 R_bl
Cb_24_65 bit_24_65 gnd C_bl
Cbb_24_65 bitb_24_65 gnd C_bl
Rb_24_66 bit_24_66 bit_24_67 R_bl
Rbb_24_66 bitb_24_66 bitb_24_67 R_bl
Cb_24_66 bit_24_66 gnd C_bl
Cbb_24_66 bitb_24_66 gnd C_bl
Rb_24_67 bit_24_67 bit_24_68 R_bl
Rbb_24_67 bitb_24_67 bitb_24_68 R_bl
Cb_24_67 bit_24_67 gnd C_bl
Cbb_24_67 bitb_24_67 gnd C_bl
Rb_24_68 bit_24_68 bit_24_69 R_bl
Rbb_24_68 bitb_24_68 bitb_24_69 R_bl
Cb_24_68 bit_24_68 gnd C_bl
Cbb_24_68 bitb_24_68 gnd C_bl
Rb_24_69 bit_24_69 bit_24_70 R_bl
Rbb_24_69 bitb_24_69 bitb_24_70 R_bl
Cb_24_69 bit_24_69 gnd C_bl
Cbb_24_69 bitb_24_69 gnd C_bl
Rb_24_70 bit_24_70 bit_24_71 R_bl
Rbb_24_70 bitb_24_70 bitb_24_71 R_bl
Cb_24_70 bit_24_70 gnd C_bl
Cbb_24_70 bitb_24_70 gnd C_bl
Rb_24_71 bit_24_71 bit_24_72 R_bl
Rbb_24_71 bitb_24_71 bitb_24_72 R_bl
Cb_24_71 bit_24_71 gnd C_bl
Cbb_24_71 bitb_24_71 gnd C_bl
Rb_24_72 bit_24_72 bit_24_73 R_bl
Rbb_24_72 bitb_24_72 bitb_24_73 R_bl
Cb_24_72 bit_24_72 gnd C_bl
Cbb_24_72 bitb_24_72 gnd C_bl
Rb_24_73 bit_24_73 bit_24_74 R_bl
Rbb_24_73 bitb_24_73 bitb_24_74 R_bl
Cb_24_73 bit_24_73 gnd C_bl
Cbb_24_73 bitb_24_73 gnd C_bl
Rb_24_74 bit_24_74 bit_24_75 R_bl
Rbb_24_74 bitb_24_74 bitb_24_75 R_bl
Cb_24_74 bit_24_74 gnd C_bl
Cbb_24_74 bitb_24_74 gnd C_bl
Rb_24_75 bit_24_75 bit_24_76 R_bl
Rbb_24_75 bitb_24_75 bitb_24_76 R_bl
Cb_24_75 bit_24_75 gnd C_bl
Cbb_24_75 bitb_24_75 gnd C_bl
Rb_24_76 bit_24_76 bit_24_77 R_bl
Rbb_24_76 bitb_24_76 bitb_24_77 R_bl
Cb_24_76 bit_24_76 gnd C_bl
Cbb_24_76 bitb_24_76 gnd C_bl
Rb_24_77 bit_24_77 bit_24_78 R_bl
Rbb_24_77 bitb_24_77 bitb_24_78 R_bl
Cb_24_77 bit_24_77 gnd C_bl
Cbb_24_77 bitb_24_77 gnd C_bl
Rb_24_78 bit_24_78 bit_24_79 R_bl
Rbb_24_78 bitb_24_78 bitb_24_79 R_bl
Cb_24_78 bit_24_78 gnd C_bl
Cbb_24_78 bitb_24_78 gnd C_bl
Rb_24_79 bit_24_79 bit_24_80 R_bl
Rbb_24_79 bitb_24_79 bitb_24_80 R_bl
Cb_24_79 bit_24_79 gnd C_bl
Cbb_24_79 bitb_24_79 gnd C_bl
Rb_24_80 bit_24_80 bit_24_81 R_bl
Rbb_24_80 bitb_24_80 bitb_24_81 R_bl
Cb_24_80 bit_24_80 gnd C_bl
Cbb_24_80 bitb_24_80 gnd C_bl
Rb_24_81 bit_24_81 bit_24_82 R_bl
Rbb_24_81 bitb_24_81 bitb_24_82 R_bl
Cb_24_81 bit_24_81 gnd C_bl
Cbb_24_81 bitb_24_81 gnd C_bl
Rb_24_82 bit_24_82 bit_24_83 R_bl
Rbb_24_82 bitb_24_82 bitb_24_83 R_bl
Cb_24_82 bit_24_82 gnd C_bl
Cbb_24_82 bitb_24_82 gnd C_bl
Rb_24_83 bit_24_83 bit_24_84 R_bl
Rbb_24_83 bitb_24_83 bitb_24_84 R_bl
Cb_24_83 bit_24_83 gnd C_bl
Cbb_24_83 bitb_24_83 gnd C_bl
Rb_24_84 bit_24_84 bit_24_85 R_bl
Rbb_24_84 bitb_24_84 bitb_24_85 R_bl
Cb_24_84 bit_24_84 gnd C_bl
Cbb_24_84 bitb_24_84 gnd C_bl
Rb_24_85 bit_24_85 bit_24_86 R_bl
Rbb_24_85 bitb_24_85 bitb_24_86 R_bl
Cb_24_85 bit_24_85 gnd C_bl
Cbb_24_85 bitb_24_85 gnd C_bl
Rb_24_86 bit_24_86 bit_24_87 R_bl
Rbb_24_86 bitb_24_86 bitb_24_87 R_bl
Cb_24_86 bit_24_86 gnd C_bl
Cbb_24_86 bitb_24_86 gnd C_bl
Rb_24_87 bit_24_87 bit_24_88 R_bl
Rbb_24_87 bitb_24_87 bitb_24_88 R_bl
Cb_24_87 bit_24_87 gnd C_bl
Cbb_24_87 bitb_24_87 gnd C_bl
Rb_24_88 bit_24_88 bit_24_89 R_bl
Rbb_24_88 bitb_24_88 bitb_24_89 R_bl
Cb_24_88 bit_24_88 gnd C_bl
Cbb_24_88 bitb_24_88 gnd C_bl
Rb_24_89 bit_24_89 bit_24_90 R_bl
Rbb_24_89 bitb_24_89 bitb_24_90 R_bl
Cb_24_89 bit_24_89 gnd C_bl
Cbb_24_89 bitb_24_89 gnd C_bl
Rb_24_90 bit_24_90 bit_24_91 R_bl
Rbb_24_90 bitb_24_90 bitb_24_91 R_bl
Cb_24_90 bit_24_90 gnd C_bl
Cbb_24_90 bitb_24_90 gnd C_bl
Rb_24_91 bit_24_91 bit_24_92 R_bl
Rbb_24_91 bitb_24_91 bitb_24_92 R_bl
Cb_24_91 bit_24_91 gnd C_bl
Cbb_24_91 bitb_24_91 gnd C_bl
Rb_24_92 bit_24_92 bit_24_93 R_bl
Rbb_24_92 bitb_24_92 bitb_24_93 R_bl
Cb_24_92 bit_24_92 gnd C_bl
Cbb_24_92 bitb_24_92 gnd C_bl
Rb_24_93 bit_24_93 bit_24_94 R_bl
Rbb_24_93 bitb_24_93 bitb_24_94 R_bl
Cb_24_93 bit_24_93 gnd C_bl
Cbb_24_93 bitb_24_93 gnd C_bl
Rb_24_94 bit_24_94 bit_24_95 R_bl
Rbb_24_94 bitb_24_94 bitb_24_95 R_bl
Cb_24_94 bit_24_94 gnd C_bl
Cbb_24_94 bitb_24_94 gnd C_bl
Rb_24_95 bit_24_95 bit_24_96 R_bl
Rbb_24_95 bitb_24_95 bitb_24_96 R_bl
Cb_24_95 bit_24_95 gnd C_bl
Cbb_24_95 bitb_24_95 gnd C_bl
Rb_24_96 bit_24_96 bit_24_97 R_bl
Rbb_24_96 bitb_24_96 bitb_24_97 R_bl
Cb_24_96 bit_24_96 gnd C_bl
Cbb_24_96 bitb_24_96 gnd C_bl
Rb_24_97 bit_24_97 bit_24_98 R_bl
Rbb_24_97 bitb_24_97 bitb_24_98 R_bl
Cb_24_97 bit_24_97 gnd C_bl
Cbb_24_97 bitb_24_97 gnd C_bl
Rb_24_98 bit_24_98 bit_24_99 R_bl
Rbb_24_98 bitb_24_98 bitb_24_99 R_bl
Cb_24_98 bit_24_98 gnd C_bl
Cbb_24_98 bitb_24_98 gnd C_bl
Rb_24_99 bit_24_99 bit_24_100 R_bl
Rbb_24_99 bitb_24_99 bitb_24_100 R_bl
Cb_24_99 bit_24_99 gnd C_bl
Cbb_24_99 bitb_24_99 gnd C_bl
Rb_25_0 bit_25_0 bit_25_1 R_bl
Rbb_25_0 bitb_25_0 bitb_25_1 R_bl
Cb_25_0 bit_25_0 gnd C_bl
Cbb_25_0 bitb_25_0 gnd C_bl
Rb_25_1 bit_25_1 bit_25_2 R_bl
Rbb_25_1 bitb_25_1 bitb_25_2 R_bl
Cb_25_1 bit_25_1 gnd C_bl
Cbb_25_1 bitb_25_1 gnd C_bl
Rb_25_2 bit_25_2 bit_25_3 R_bl
Rbb_25_2 bitb_25_2 bitb_25_3 R_bl
Cb_25_2 bit_25_2 gnd C_bl
Cbb_25_2 bitb_25_2 gnd C_bl
Rb_25_3 bit_25_3 bit_25_4 R_bl
Rbb_25_3 bitb_25_3 bitb_25_4 R_bl
Cb_25_3 bit_25_3 gnd C_bl
Cbb_25_3 bitb_25_3 gnd C_bl
Rb_25_4 bit_25_4 bit_25_5 R_bl
Rbb_25_4 bitb_25_4 bitb_25_5 R_bl
Cb_25_4 bit_25_4 gnd C_bl
Cbb_25_4 bitb_25_4 gnd C_bl
Rb_25_5 bit_25_5 bit_25_6 R_bl
Rbb_25_5 bitb_25_5 bitb_25_6 R_bl
Cb_25_5 bit_25_5 gnd C_bl
Cbb_25_5 bitb_25_5 gnd C_bl
Rb_25_6 bit_25_6 bit_25_7 R_bl
Rbb_25_6 bitb_25_6 bitb_25_7 R_bl
Cb_25_6 bit_25_6 gnd C_bl
Cbb_25_6 bitb_25_6 gnd C_bl
Rb_25_7 bit_25_7 bit_25_8 R_bl
Rbb_25_7 bitb_25_7 bitb_25_8 R_bl
Cb_25_7 bit_25_7 gnd C_bl
Cbb_25_7 bitb_25_7 gnd C_bl
Rb_25_8 bit_25_8 bit_25_9 R_bl
Rbb_25_8 bitb_25_8 bitb_25_9 R_bl
Cb_25_8 bit_25_8 gnd C_bl
Cbb_25_8 bitb_25_8 gnd C_bl
Rb_25_9 bit_25_9 bit_25_10 R_bl
Rbb_25_9 bitb_25_9 bitb_25_10 R_bl
Cb_25_9 bit_25_9 gnd C_bl
Cbb_25_9 bitb_25_9 gnd C_bl
Rb_25_10 bit_25_10 bit_25_11 R_bl
Rbb_25_10 bitb_25_10 bitb_25_11 R_bl
Cb_25_10 bit_25_10 gnd C_bl
Cbb_25_10 bitb_25_10 gnd C_bl
Rb_25_11 bit_25_11 bit_25_12 R_bl
Rbb_25_11 bitb_25_11 bitb_25_12 R_bl
Cb_25_11 bit_25_11 gnd C_bl
Cbb_25_11 bitb_25_11 gnd C_bl
Rb_25_12 bit_25_12 bit_25_13 R_bl
Rbb_25_12 bitb_25_12 bitb_25_13 R_bl
Cb_25_12 bit_25_12 gnd C_bl
Cbb_25_12 bitb_25_12 gnd C_bl
Rb_25_13 bit_25_13 bit_25_14 R_bl
Rbb_25_13 bitb_25_13 bitb_25_14 R_bl
Cb_25_13 bit_25_13 gnd C_bl
Cbb_25_13 bitb_25_13 gnd C_bl
Rb_25_14 bit_25_14 bit_25_15 R_bl
Rbb_25_14 bitb_25_14 bitb_25_15 R_bl
Cb_25_14 bit_25_14 gnd C_bl
Cbb_25_14 bitb_25_14 gnd C_bl
Rb_25_15 bit_25_15 bit_25_16 R_bl
Rbb_25_15 bitb_25_15 bitb_25_16 R_bl
Cb_25_15 bit_25_15 gnd C_bl
Cbb_25_15 bitb_25_15 gnd C_bl
Rb_25_16 bit_25_16 bit_25_17 R_bl
Rbb_25_16 bitb_25_16 bitb_25_17 R_bl
Cb_25_16 bit_25_16 gnd C_bl
Cbb_25_16 bitb_25_16 gnd C_bl
Rb_25_17 bit_25_17 bit_25_18 R_bl
Rbb_25_17 bitb_25_17 bitb_25_18 R_bl
Cb_25_17 bit_25_17 gnd C_bl
Cbb_25_17 bitb_25_17 gnd C_bl
Rb_25_18 bit_25_18 bit_25_19 R_bl
Rbb_25_18 bitb_25_18 bitb_25_19 R_bl
Cb_25_18 bit_25_18 gnd C_bl
Cbb_25_18 bitb_25_18 gnd C_bl
Rb_25_19 bit_25_19 bit_25_20 R_bl
Rbb_25_19 bitb_25_19 bitb_25_20 R_bl
Cb_25_19 bit_25_19 gnd C_bl
Cbb_25_19 bitb_25_19 gnd C_bl
Rb_25_20 bit_25_20 bit_25_21 R_bl
Rbb_25_20 bitb_25_20 bitb_25_21 R_bl
Cb_25_20 bit_25_20 gnd C_bl
Cbb_25_20 bitb_25_20 gnd C_bl
Rb_25_21 bit_25_21 bit_25_22 R_bl
Rbb_25_21 bitb_25_21 bitb_25_22 R_bl
Cb_25_21 bit_25_21 gnd C_bl
Cbb_25_21 bitb_25_21 gnd C_bl
Rb_25_22 bit_25_22 bit_25_23 R_bl
Rbb_25_22 bitb_25_22 bitb_25_23 R_bl
Cb_25_22 bit_25_22 gnd C_bl
Cbb_25_22 bitb_25_22 gnd C_bl
Rb_25_23 bit_25_23 bit_25_24 R_bl
Rbb_25_23 bitb_25_23 bitb_25_24 R_bl
Cb_25_23 bit_25_23 gnd C_bl
Cbb_25_23 bitb_25_23 gnd C_bl
Rb_25_24 bit_25_24 bit_25_25 R_bl
Rbb_25_24 bitb_25_24 bitb_25_25 R_bl
Cb_25_24 bit_25_24 gnd C_bl
Cbb_25_24 bitb_25_24 gnd C_bl
Rb_25_25 bit_25_25 bit_25_26 R_bl
Rbb_25_25 bitb_25_25 bitb_25_26 R_bl
Cb_25_25 bit_25_25 gnd C_bl
Cbb_25_25 bitb_25_25 gnd C_bl
Rb_25_26 bit_25_26 bit_25_27 R_bl
Rbb_25_26 bitb_25_26 bitb_25_27 R_bl
Cb_25_26 bit_25_26 gnd C_bl
Cbb_25_26 bitb_25_26 gnd C_bl
Rb_25_27 bit_25_27 bit_25_28 R_bl
Rbb_25_27 bitb_25_27 bitb_25_28 R_bl
Cb_25_27 bit_25_27 gnd C_bl
Cbb_25_27 bitb_25_27 gnd C_bl
Rb_25_28 bit_25_28 bit_25_29 R_bl
Rbb_25_28 bitb_25_28 bitb_25_29 R_bl
Cb_25_28 bit_25_28 gnd C_bl
Cbb_25_28 bitb_25_28 gnd C_bl
Rb_25_29 bit_25_29 bit_25_30 R_bl
Rbb_25_29 bitb_25_29 bitb_25_30 R_bl
Cb_25_29 bit_25_29 gnd C_bl
Cbb_25_29 bitb_25_29 gnd C_bl
Rb_25_30 bit_25_30 bit_25_31 R_bl
Rbb_25_30 bitb_25_30 bitb_25_31 R_bl
Cb_25_30 bit_25_30 gnd C_bl
Cbb_25_30 bitb_25_30 gnd C_bl
Rb_25_31 bit_25_31 bit_25_32 R_bl
Rbb_25_31 bitb_25_31 bitb_25_32 R_bl
Cb_25_31 bit_25_31 gnd C_bl
Cbb_25_31 bitb_25_31 gnd C_bl
Rb_25_32 bit_25_32 bit_25_33 R_bl
Rbb_25_32 bitb_25_32 bitb_25_33 R_bl
Cb_25_32 bit_25_32 gnd C_bl
Cbb_25_32 bitb_25_32 gnd C_bl
Rb_25_33 bit_25_33 bit_25_34 R_bl
Rbb_25_33 bitb_25_33 bitb_25_34 R_bl
Cb_25_33 bit_25_33 gnd C_bl
Cbb_25_33 bitb_25_33 gnd C_bl
Rb_25_34 bit_25_34 bit_25_35 R_bl
Rbb_25_34 bitb_25_34 bitb_25_35 R_bl
Cb_25_34 bit_25_34 gnd C_bl
Cbb_25_34 bitb_25_34 gnd C_bl
Rb_25_35 bit_25_35 bit_25_36 R_bl
Rbb_25_35 bitb_25_35 bitb_25_36 R_bl
Cb_25_35 bit_25_35 gnd C_bl
Cbb_25_35 bitb_25_35 gnd C_bl
Rb_25_36 bit_25_36 bit_25_37 R_bl
Rbb_25_36 bitb_25_36 bitb_25_37 R_bl
Cb_25_36 bit_25_36 gnd C_bl
Cbb_25_36 bitb_25_36 gnd C_bl
Rb_25_37 bit_25_37 bit_25_38 R_bl
Rbb_25_37 bitb_25_37 bitb_25_38 R_bl
Cb_25_37 bit_25_37 gnd C_bl
Cbb_25_37 bitb_25_37 gnd C_bl
Rb_25_38 bit_25_38 bit_25_39 R_bl
Rbb_25_38 bitb_25_38 bitb_25_39 R_bl
Cb_25_38 bit_25_38 gnd C_bl
Cbb_25_38 bitb_25_38 gnd C_bl
Rb_25_39 bit_25_39 bit_25_40 R_bl
Rbb_25_39 bitb_25_39 bitb_25_40 R_bl
Cb_25_39 bit_25_39 gnd C_bl
Cbb_25_39 bitb_25_39 gnd C_bl
Rb_25_40 bit_25_40 bit_25_41 R_bl
Rbb_25_40 bitb_25_40 bitb_25_41 R_bl
Cb_25_40 bit_25_40 gnd C_bl
Cbb_25_40 bitb_25_40 gnd C_bl
Rb_25_41 bit_25_41 bit_25_42 R_bl
Rbb_25_41 bitb_25_41 bitb_25_42 R_bl
Cb_25_41 bit_25_41 gnd C_bl
Cbb_25_41 bitb_25_41 gnd C_bl
Rb_25_42 bit_25_42 bit_25_43 R_bl
Rbb_25_42 bitb_25_42 bitb_25_43 R_bl
Cb_25_42 bit_25_42 gnd C_bl
Cbb_25_42 bitb_25_42 gnd C_bl
Rb_25_43 bit_25_43 bit_25_44 R_bl
Rbb_25_43 bitb_25_43 bitb_25_44 R_bl
Cb_25_43 bit_25_43 gnd C_bl
Cbb_25_43 bitb_25_43 gnd C_bl
Rb_25_44 bit_25_44 bit_25_45 R_bl
Rbb_25_44 bitb_25_44 bitb_25_45 R_bl
Cb_25_44 bit_25_44 gnd C_bl
Cbb_25_44 bitb_25_44 gnd C_bl
Rb_25_45 bit_25_45 bit_25_46 R_bl
Rbb_25_45 bitb_25_45 bitb_25_46 R_bl
Cb_25_45 bit_25_45 gnd C_bl
Cbb_25_45 bitb_25_45 gnd C_bl
Rb_25_46 bit_25_46 bit_25_47 R_bl
Rbb_25_46 bitb_25_46 bitb_25_47 R_bl
Cb_25_46 bit_25_46 gnd C_bl
Cbb_25_46 bitb_25_46 gnd C_bl
Rb_25_47 bit_25_47 bit_25_48 R_bl
Rbb_25_47 bitb_25_47 bitb_25_48 R_bl
Cb_25_47 bit_25_47 gnd C_bl
Cbb_25_47 bitb_25_47 gnd C_bl
Rb_25_48 bit_25_48 bit_25_49 R_bl
Rbb_25_48 bitb_25_48 bitb_25_49 R_bl
Cb_25_48 bit_25_48 gnd C_bl
Cbb_25_48 bitb_25_48 gnd C_bl
Rb_25_49 bit_25_49 bit_25_50 R_bl
Rbb_25_49 bitb_25_49 bitb_25_50 R_bl
Cb_25_49 bit_25_49 gnd C_bl
Cbb_25_49 bitb_25_49 gnd C_bl
Rb_25_50 bit_25_50 bit_25_51 R_bl
Rbb_25_50 bitb_25_50 bitb_25_51 R_bl
Cb_25_50 bit_25_50 gnd C_bl
Cbb_25_50 bitb_25_50 gnd C_bl
Rb_25_51 bit_25_51 bit_25_52 R_bl
Rbb_25_51 bitb_25_51 bitb_25_52 R_bl
Cb_25_51 bit_25_51 gnd C_bl
Cbb_25_51 bitb_25_51 gnd C_bl
Rb_25_52 bit_25_52 bit_25_53 R_bl
Rbb_25_52 bitb_25_52 bitb_25_53 R_bl
Cb_25_52 bit_25_52 gnd C_bl
Cbb_25_52 bitb_25_52 gnd C_bl
Rb_25_53 bit_25_53 bit_25_54 R_bl
Rbb_25_53 bitb_25_53 bitb_25_54 R_bl
Cb_25_53 bit_25_53 gnd C_bl
Cbb_25_53 bitb_25_53 gnd C_bl
Rb_25_54 bit_25_54 bit_25_55 R_bl
Rbb_25_54 bitb_25_54 bitb_25_55 R_bl
Cb_25_54 bit_25_54 gnd C_bl
Cbb_25_54 bitb_25_54 gnd C_bl
Rb_25_55 bit_25_55 bit_25_56 R_bl
Rbb_25_55 bitb_25_55 bitb_25_56 R_bl
Cb_25_55 bit_25_55 gnd C_bl
Cbb_25_55 bitb_25_55 gnd C_bl
Rb_25_56 bit_25_56 bit_25_57 R_bl
Rbb_25_56 bitb_25_56 bitb_25_57 R_bl
Cb_25_56 bit_25_56 gnd C_bl
Cbb_25_56 bitb_25_56 gnd C_bl
Rb_25_57 bit_25_57 bit_25_58 R_bl
Rbb_25_57 bitb_25_57 bitb_25_58 R_bl
Cb_25_57 bit_25_57 gnd C_bl
Cbb_25_57 bitb_25_57 gnd C_bl
Rb_25_58 bit_25_58 bit_25_59 R_bl
Rbb_25_58 bitb_25_58 bitb_25_59 R_bl
Cb_25_58 bit_25_58 gnd C_bl
Cbb_25_58 bitb_25_58 gnd C_bl
Rb_25_59 bit_25_59 bit_25_60 R_bl
Rbb_25_59 bitb_25_59 bitb_25_60 R_bl
Cb_25_59 bit_25_59 gnd C_bl
Cbb_25_59 bitb_25_59 gnd C_bl
Rb_25_60 bit_25_60 bit_25_61 R_bl
Rbb_25_60 bitb_25_60 bitb_25_61 R_bl
Cb_25_60 bit_25_60 gnd C_bl
Cbb_25_60 bitb_25_60 gnd C_bl
Rb_25_61 bit_25_61 bit_25_62 R_bl
Rbb_25_61 bitb_25_61 bitb_25_62 R_bl
Cb_25_61 bit_25_61 gnd C_bl
Cbb_25_61 bitb_25_61 gnd C_bl
Rb_25_62 bit_25_62 bit_25_63 R_bl
Rbb_25_62 bitb_25_62 bitb_25_63 R_bl
Cb_25_62 bit_25_62 gnd C_bl
Cbb_25_62 bitb_25_62 gnd C_bl
Rb_25_63 bit_25_63 bit_25_64 R_bl
Rbb_25_63 bitb_25_63 bitb_25_64 R_bl
Cb_25_63 bit_25_63 gnd C_bl
Cbb_25_63 bitb_25_63 gnd C_bl
Rb_25_64 bit_25_64 bit_25_65 R_bl
Rbb_25_64 bitb_25_64 bitb_25_65 R_bl
Cb_25_64 bit_25_64 gnd C_bl
Cbb_25_64 bitb_25_64 gnd C_bl
Rb_25_65 bit_25_65 bit_25_66 R_bl
Rbb_25_65 bitb_25_65 bitb_25_66 R_bl
Cb_25_65 bit_25_65 gnd C_bl
Cbb_25_65 bitb_25_65 gnd C_bl
Rb_25_66 bit_25_66 bit_25_67 R_bl
Rbb_25_66 bitb_25_66 bitb_25_67 R_bl
Cb_25_66 bit_25_66 gnd C_bl
Cbb_25_66 bitb_25_66 gnd C_bl
Rb_25_67 bit_25_67 bit_25_68 R_bl
Rbb_25_67 bitb_25_67 bitb_25_68 R_bl
Cb_25_67 bit_25_67 gnd C_bl
Cbb_25_67 bitb_25_67 gnd C_bl
Rb_25_68 bit_25_68 bit_25_69 R_bl
Rbb_25_68 bitb_25_68 bitb_25_69 R_bl
Cb_25_68 bit_25_68 gnd C_bl
Cbb_25_68 bitb_25_68 gnd C_bl
Rb_25_69 bit_25_69 bit_25_70 R_bl
Rbb_25_69 bitb_25_69 bitb_25_70 R_bl
Cb_25_69 bit_25_69 gnd C_bl
Cbb_25_69 bitb_25_69 gnd C_bl
Rb_25_70 bit_25_70 bit_25_71 R_bl
Rbb_25_70 bitb_25_70 bitb_25_71 R_bl
Cb_25_70 bit_25_70 gnd C_bl
Cbb_25_70 bitb_25_70 gnd C_bl
Rb_25_71 bit_25_71 bit_25_72 R_bl
Rbb_25_71 bitb_25_71 bitb_25_72 R_bl
Cb_25_71 bit_25_71 gnd C_bl
Cbb_25_71 bitb_25_71 gnd C_bl
Rb_25_72 bit_25_72 bit_25_73 R_bl
Rbb_25_72 bitb_25_72 bitb_25_73 R_bl
Cb_25_72 bit_25_72 gnd C_bl
Cbb_25_72 bitb_25_72 gnd C_bl
Rb_25_73 bit_25_73 bit_25_74 R_bl
Rbb_25_73 bitb_25_73 bitb_25_74 R_bl
Cb_25_73 bit_25_73 gnd C_bl
Cbb_25_73 bitb_25_73 gnd C_bl
Rb_25_74 bit_25_74 bit_25_75 R_bl
Rbb_25_74 bitb_25_74 bitb_25_75 R_bl
Cb_25_74 bit_25_74 gnd C_bl
Cbb_25_74 bitb_25_74 gnd C_bl
Rb_25_75 bit_25_75 bit_25_76 R_bl
Rbb_25_75 bitb_25_75 bitb_25_76 R_bl
Cb_25_75 bit_25_75 gnd C_bl
Cbb_25_75 bitb_25_75 gnd C_bl
Rb_25_76 bit_25_76 bit_25_77 R_bl
Rbb_25_76 bitb_25_76 bitb_25_77 R_bl
Cb_25_76 bit_25_76 gnd C_bl
Cbb_25_76 bitb_25_76 gnd C_bl
Rb_25_77 bit_25_77 bit_25_78 R_bl
Rbb_25_77 bitb_25_77 bitb_25_78 R_bl
Cb_25_77 bit_25_77 gnd C_bl
Cbb_25_77 bitb_25_77 gnd C_bl
Rb_25_78 bit_25_78 bit_25_79 R_bl
Rbb_25_78 bitb_25_78 bitb_25_79 R_bl
Cb_25_78 bit_25_78 gnd C_bl
Cbb_25_78 bitb_25_78 gnd C_bl
Rb_25_79 bit_25_79 bit_25_80 R_bl
Rbb_25_79 bitb_25_79 bitb_25_80 R_bl
Cb_25_79 bit_25_79 gnd C_bl
Cbb_25_79 bitb_25_79 gnd C_bl
Rb_25_80 bit_25_80 bit_25_81 R_bl
Rbb_25_80 bitb_25_80 bitb_25_81 R_bl
Cb_25_80 bit_25_80 gnd C_bl
Cbb_25_80 bitb_25_80 gnd C_bl
Rb_25_81 bit_25_81 bit_25_82 R_bl
Rbb_25_81 bitb_25_81 bitb_25_82 R_bl
Cb_25_81 bit_25_81 gnd C_bl
Cbb_25_81 bitb_25_81 gnd C_bl
Rb_25_82 bit_25_82 bit_25_83 R_bl
Rbb_25_82 bitb_25_82 bitb_25_83 R_bl
Cb_25_82 bit_25_82 gnd C_bl
Cbb_25_82 bitb_25_82 gnd C_bl
Rb_25_83 bit_25_83 bit_25_84 R_bl
Rbb_25_83 bitb_25_83 bitb_25_84 R_bl
Cb_25_83 bit_25_83 gnd C_bl
Cbb_25_83 bitb_25_83 gnd C_bl
Rb_25_84 bit_25_84 bit_25_85 R_bl
Rbb_25_84 bitb_25_84 bitb_25_85 R_bl
Cb_25_84 bit_25_84 gnd C_bl
Cbb_25_84 bitb_25_84 gnd C_bl
Rb_25_85 bit_25_85 bit_25_86 R_bl
Rbb_25_85 bitb_25_85 bitb_25_86 R_bl
Cb_25_85 bit_25_85 gnd C_bl
Cbb_25_85 bitb_25_85 gnd C_bl
Rb_25_86 bit_25_86 bit_25_87 R_bl
Rbb_25_86 bitb_25_86 bitb_25_87 R_bl
Cb_25_86 bit_25_86 gnd C_bl
Cbb_25_86 bitb_25_86 gnd C_bl
Rb_25_87 bit_25_87 bit_25_88 R_bl
Rbb_25_87 bitb_25_87 bitb_25_88 R_bl
Cb_25_87 bit_25_87 gnd C_bl
Cbb_25_87 bitb_25_87 gnd C_bl
Rb_25_88 bit_25_88 bit_25_89 R_bl
Rbb_25_88 bitb_25_88 bitb_25_89 R_bl
Cb_25_88 bit_25_88 gnd C_bl
Cbb_25_88 bitb_25_88 gnd C_bl
Rb_25_89 bit_25_89 bit_25_90 R_bl
Rbb_25_89 bitb_25_89 bitb_25_90 R_bl
Cb_25_89 bit_25_89 gnd C_bl
Cbb_25_89 bitb_25_89 gnd C_bl
Rb_25_90 bit_25_90 bit_25_91 R_bl
Rbb_25_90 bitb_25_90 bitb_25_91 R_bl
Cb_25_90 bit_25_90 gnd C_bl
Cbb_25_90 bitb_25_90 gnd C_bl
Rb_25_91 bit_25_91 bit_25_92 R_bl
Rbb_25_91 bitb_25_91 bitb_25_92 R_bl
Cb_25_91 bit_25_91 gnd C_bl
Cbb_25_91 bitb_25_91 gnd C_bl
Rb_25_92 bit_25_92 bit_25_93 R_bl
Rbb_25_92 bitb_25_92 bitb_25_93 R_bl
Cb_25_92 bit_25_92 gnd C_bl
Cbb_25_92 bitb_25_92 gnd C_bl
Rb_25_93 bit_25_93 bit_25_94 R_bl
Rbb_25_93 bitb_25_93 bitb_25_94 R_bl
Cb_25_93 bit_25_93 gnd C_bl
Cbb_25_93 bitb_25_93 gnd C_bl
Rb_25_94 bit_25_94 bit_25_95 R_bl
Rbb_25_94 bitb_25_94 bitb_25_95 R_bl
Cb_25_94 bit_25_94 gnd C_bl
Cbb_25_94 bitb_25_94 gnd C_bl
Rb_25_95 bit_25_95 bit_25_96 R_bl
Rbb_25_95 bitb_25_95 bitb_25_96 R_bl
Cb_25_95 bit_25_95 gnd C_bl
Cbb_25_95 bitb_25_95 gnd C_bl
Rb_25_96 bit_25_96 bit_25_97 R_bl
Rbb_25_96 bitb_25_96 bitb_25_97 R_bl
Cb_25_96 bit_25_96 gnd C_bl
Cbb_25_96 bitb_25_96 gnd C_bl
Rb_25_97 bit_25_97 bit_25_98 R_bl
Rbb_25_97 bitb_25_97 bitb_25_98 R_bl
Cb_25_97 bit_25_97 gnd C_bl
Cbb_25_97 bitb_25_97 gnd C_bl
Rb_25_98 bit_25_98 bit_25_99 R_bl
Rbb_25_98 bitb_25_98 bitb_25_99 R_bl
Cb_25_98 bit_25_98 gnd C_bl
Cbb_25_98 bitb_25_98 gnd C_bl
Rb_25_99 bit_25_99 bit_25_100 R_bl
Rbb_25_99 bitb_25_99 bitb_25_100 R_bl
Cb_25_99 bit_25_99 gnd C_bl
Cbb_25_99 bitb_25_99 gnd C_bl
Rb_26_0 bit_26_0 bit_26_1 R_bl
Rbb_26_0 bitb_26_0 bitb_26_1 R_bl
Cb_26_0 bit_26_0 gnd C_bl
Cbb_26_0 bitb_26_0 gnd C_bl
Rb_26_1 bit_26_1 bit_26_2 R_bl
Rbb_26_1 bitb_26_1 bitb_26_2 R_bl
Cb_26_1 bit_26_1 gnd C_bl
Cbb_26_1 bitb_26_1 gnd C_bl
Rb_26_2 bit_26_2 bit_26_3 R_bl
Rbb_26_2 bitb_26_2 bitb_26_3 R_bl
Cb_26_2 bit_26_2 gnd C_bl
Cbb_26_2 bitb_26_2 gnd C_bl
Rb_26_3 bit_26_3 bit_26_4 R_bl
Rbb_26_3 bitb_26_3 bitb_26_4 R_bl
Cb_26_3 bit_26_3 gnd C_bl
Cbb_26_3 bitb_26_3 gnd C_bl
Rb_26_4 bit_26_4 bit_26_5 R_bl
Rbb_26_4 bitb_26_4 bitb_26_5 R_bl
Cb_26_4 bit_26_4 gnd C_bl
Cbb_26_4 bitb_26_4 gnd C_bl
Rb_26_5 bit_26_5 bit_26_6 R_bl
Rbb_26_5 bitb_26_5 bitb_26_6 R_bl
Cb_26_5 bit_26_5 gnd C_bl
Cbb_26_5 bitb_26_5 gnd C_bl
Rb_26_6 bit_26_6 bit_26_7 R_bl
Rbb_26_6 bitb_26_6 bitb_26_7 R_bl
Cb_26_6 bit_26_6 gnd C_bl
Cbb_26_6 bitb_26_6 gnd C_bl
Rb_26_7 bit_26_7 bit_26_8 R_bl
Rbb_26_7 bitb_26_7 bitb_26_8 R_bl
Cb_26_7 bit_26_7 gnd C_bl
Cbb_26_7 bitb_26_7 gnd C_bl
Rb_26_8 bit_26_8 bit_26_9 R_bl
Rbb_26_8 bitb_26_8 bitb_26_9 R_bl
Cb_26_8 bit_26_8 gnd C_bl
Cbb_26_8 bitb_26_8 gnd C_bl
Rb_26_9 bit_26_9 bit_26_10 R_bl
Rbb_26_9 bitb_26_9 bitb_26_10 R_bl
Cb_26_9 bit_26_9 gnd C_bl
Cbb_26_9 bitb_26_9 gnd C_bl
Rb_26_10 bit_26_10 bit_26_11 R_bl
Rbb_26_10 bitb_26_10 bitb_26_11 R_bl
Cb_26_10 bit_26_10 gnd C_bl
Cbb_26_10 bitb_26_10 gnd C_bl
Rb_26_11 bit_26_11 bit_26_12 R_bl
Rbb_26_11 bitb_26_11 bitb_26_12 R_bl
Cb_26_11 bit_26_11 gnd C_bl
Cbb_26_11 bitb_26_11 gnd C_bl
Rb_26_12 bit_26_12 bit_26_13 R_bl
Rbb_26_12 bitb_26_12 bitb_26_13 R_bl
Cb_26_12 bit_26_12 gnd C_bl
Cbb_26_12 bitb_26_12 gnd C_bl
Rb_26_13 bit_26_13 bit_26_14 R_bl
Rbb_26_13 bitb_26_13 bitb_26_14 R_bl
Cb_26_13 bit_26_13 gnd C_bl
Cbb_26_13 bitb_26_13 gnd C_bl
Rb_26_14 bit_26_14 bit_26_15 R_bl
Rbb_26_14 bitb_26_14 bitb_26_15 R_bl
Cb_26_14 bit_26_14 gnd C_bl
Cbb_26_14 bitb_26_14 gnd C_bl
Rb_26_15 bit_26_15 bit_26_16 R_bl
Rbb_26_15 bitb_26_15 bitb_26_16 R_bl
Cb_26_15 bit_26_15 gnd C_bl
Cbb_26_15 bitb_26_15 gnd C_bl
Rb_26_16 bit_26_16 bit_26_17 R_bl
Rbb_26_16 bitb_26_16 bitb_26_17 R_bl
Cb_26_16 bit_26_16 gnd C_bl
Cbb_26_16 bitb_26_16 gnd C_bl
Rb_26_17 bit_26_17 bit_26_18 R_bl
Rbb_26_17 bitb_26_17 bitb_26_18 R_bl
Cb_26_17 bit_26_17 gnd C_bl
Cbb_26_17 bitb_26_17 gnd C_bl
Rb_26_18 bit_26_18 bit_26_19 R_bl
Rbb_26_18 bitb_26_18 bitb_26_19 R_bl
Cb_26_18 bit_26_18 gnd C_bl
Cbb_26_18 bitb_26_18 gnd C_bl
Rb_26_19 bit_26_19 bit_26_20 R_bl
Rbb_26_19 bitb_26_19 bitb_26_20 R_bl
Cb_26_19 bit_26_19 gnd C_bl
Cbb_26_19 bitb_26_19 gnd C_bl
Rb_26_20 bit_26_20 bit_26_21 R_bl
Rbb_26_20 bitb_26_20 bitb_26_21 R_bl
Cb_26_20 bit_26_20 gnd C_bl
Cbb_26_20 bitb_26_20 gnd C_bl
Rb_26_21 bit_26_21 bit_26_22 R_bl
Rbb_26_21 bitb_26_21 bitb_26_22 R_bl
Cb_26_21 bit_26_21 gnd C_bl
Cbb_26_21 bitb_26_21 gnd C_bl
Rb_26_22 bit_26_22 bit_26_23 R_bl
Rbb_26_22 bitb_26_22 bitb_26_23 R_bl
Cb_26_22 bit_26_22 gnd C_bl
Cbb_26_22 bitb_26_22 gnd C_bl
Rb_26_23 bit_26_23 bit_26_24 R_bl
Rbb_26_23 bitb_26_23 bitb_26_24 R_bl
Cb_26_23 bit_26_23 gnd C_bl
Cbb_26_23 bitb_26_23 gnd C_bl
Rb_26_24 bit_26_24 bit_26_25 R_bl
Rbb_26_24 bitb_26_24 bitb_26_25 R_bl
Cb_26_24 bit_26_24 gnd C_bl
Cbb_26_24 bitb_26_24 gnd C_bl
Rb_26_25 bit_26_25 bit_26_26 R_bl
Rbb_26_25 bitb_26_25 bitb_26_26 R_bl
Cb_26_25 bit_26_25 gnd C_bl
Cbb_26_25 bitb_26_25 gnd C_bl
Rb_26_26 bit_26_26 bit_26_27 R_bl
Rbb_26_26 bitb_26_26 bitb_26_27 R_bl
Cb_26_26 bit_26_26 gnd C_bl
Cbb_26_26 bitb_26_26 gnd C_bl
Rb_26_27 bit_26_27 bit_26_28 R_bl
Rbb_26_27 bitb_26_27 bitb_26_28 R_bl
Cb_26_27 bit_26_27 gnd C_bl
Cbb_26_27 bitb_26_27 gnd C_bl
Rb_26_28 bit_26_28 bit_26_29 R_bl
Rbb_26_28 bitb_26_28 bitb_26_29 R_bl
Cb_26_28 bit_26_28 gnd C_bl
Cbb_26_28 bitb_26_28 gnd C_bl
Rb_26_29 bit_26_29 bit_26_30 R_bl
Rbb_26_29 bitb_26_29 bitb_26_30 R_bl
Cb_26_29 bit_26_29 gnd C_bl
Cbb_26_29 bitb_26_29 gnd C_bl
Rb_26_30 bit_26_30 bit_26_31 R_bl
Rbb_26_30 bitb_26_30 bitb_26_31 R_bl
Cb_26_30 bit_26_30 gnd C_bl
Cbb_26_30 bitb_26_30 gnd C_bl
Rb_26_31 bit_26_31 bit_26_32 R_bl
Rbb_26_31 bitb_26_31 bitb_26_32 R_bl
Cb_26_31 bit_26_31 gnd C_bl
Cbb_26_31 bitb_26_31 gnd C_bl
Rb_26_32 bit_26_32 bit_26_33 R_bl
Rbb_26_32 bitb_26_32 bitb_26_33 R_bl
Cb_26_32 bit_26_32 gnd C_bl
Cbb_26_32 bitb_26_32 gnd C_bl
Rb_26_33 bit_26_33 bit_26_34 R_bl
Rbb_26_33 bitb_26_33 bitb_26_34 R_bl
Cb_26_33 bit_26_33 gnd C_bl
Cbb_26_33 bitb_26_33 gnd C_bl
Rb_26_34 bit_26_34 bit_26_35 R_bl
Rbb_26_34 bitb_26_34 bitb_26_35 R_bl
Cb_26_34 bit_26_34 gnd C_bl
Cbb_26_34 bitb_26_34 gnd C_bl
Rb_26_35 bit_26_35 bit_26_36 R_bl
Rbb_26_35 bitb_26_35 bitb_26_36 R_bl
Cb_26_35 bit_26_35 gnd C_bl
Cbb_26_35 bitb_26_35 gnd C_bl
Rb_26_36 bit_26_36 bit_26_37 R_bl
Rbb_26_36 bitb_26_36 bitb_26_37 R_bl
Cb_26_36 bit_26_36 gnd C_bl
Cbb_26_36 bitb_26_36 gnd C_bl
Rb_26_37 bit_26_37 bit_26_38 R_bl
Rbb_26_37 bitb_26_37 bitb_26_38 R_bl
Cb_26_37 bit_26_37 gnd C_bl
Cbb_26_37 bitb_26_37 gnd C_bl
Rb_26_38 bit_26_38 bit_26_39 R_bl
Rbb_26_38 bitb_26_38 bitb_26_39 R_bl
Cb_26_38 bit_26_38 gnd C_bl
Cbb_26_38 bitb_26_38 gnd C_bl
Rb_26_39 bit_26_39 bit_26_40 R_bl
Rbb_26_39 bitb_26_39 bitb_26_40 R_bl
Cb_26_39 bit_26_39 gnd C_bl
Cbb_26_39 bitb_26_39 gnd C_bl
Rb_26_40 bit_26_40 bit_26_41 R_bl
Rbb_26_40 bitb_26_40 bitb_26_41 R_bl
Cb_26_40 bit_26_40 gnd C_bl
Cbb_26_40 bitb_26_40 gnd C_bl
Rb_26_41 bit_26_41 bit_26_42 R_bl
Rbb_26_41 bitb_26_41 bitb_26_42 R_bl
Cb_26_41 bit_26_41 gnd C_bl
Cbb_26_41 bitb_26_41 gnd C_bl
Rb_26_42 bit_26_42 bit_26_43 R_bl
Rbb_26_42 bitb_26_42 bitb_26_43 R_bl
Cb_26_42 bit_26_42 gnd C_bl
Cbb_26_42 bitb_26_42 gnd C_bl
Rb_26_43 bit_26_43 bit_26_44 R_bl
Rbb_26_43 bitb_26_43 bitb_26_44 R_bl
Cb_26_43 bit_26_43 gnd C_bl
Cbb_26_43 bitb_26_43 gnd C_bl
Rb_26_44 bit_26_44 bit_26_45 R_bl
Rbb_26_44 bitb_26_44 bitb_26_45 R_bl
Cb_26_44 bit_26_44 gnd C_bl
Cbb_26_44 bitb_26_44 gnd C_bl
Rb_26_45 bit_26_45 bit_26_46 R_bl
Rbb_26_45 bitb_26_45 bitb_26_46 R_bl
Cb_26_45 bit_26_45 gnd C_bl
Cbb_26_45 bitb_26_45 gnd C_bl
Rb_26_46 bit_26_46 bit_26_47 R_bl
Rbb_26_46 bitb_26_46 bitb_26_47 R_bl
Cb_26_46 bit_26_46 gnd C_bl
Cbb_26_46 bitb_26_46 gnd C_bl
Rb_26_47 bit_26_47 bit_26_48 R_bl
Rbb_26_47 bitb_26_47 bitb_26_48 R_bl
Cb_26_47 bit_26_47 gnd C_bl
Cbb_26_47 bitb_26_47 gnd C_bl
Rb_26_48 bit_26_48 bit_26_49 R_bl
Rbb_26_48 bitb_26_48 bitb_26_49 R_bl
Cb_26_48 bit_26_48 gnd C_bl
Cbb_26_48 bitb_26_48 gnd C_bl
Rb_26_49 bit_26_49 bit_26_50 R_bl
Rbb_26_49 bitb_26_49 bitb_26_50 R_bl
Cb_26_49 bit_26_49 gnd C_bl
Cbb_26_49 bitb_26_49 gnd C_bl
Rb_26_50 bit_26_50 bit_26_51 R_bl
Rbb_26_50 bitb_26_50 bitb_26_51 R_bl
Cb_26_50 bit_26_50 gnd C_bl
Cbb_26_50 bitb_26_50 gnd C_bl
Rb_26_51 bit_26_51 bit_26_52 R_bl
Rbb_26_51 bitb_26_51 bitb_26_52 R_bl
Cb_26_51 bit_26_51 gnd C_bl
Cbb_26_51 bitb_26_51 gnd C_bl
Rb_26_52 bit_26_52 bit_26_53 R_bl
Rbb_26_52 bitb_26_52 bitb_26_53 R_bl
Cb_26_52 bit_26_52 gnd C_bl
Cbb_26_52 bitb_26_52 gnd C_bl
Rb_26_53 bit_26_53 bit_26_54 R_bl
Rbb_26_53 bitb_26_53 bitb_26_54 R_bl
Cb_26_53 bit_26_53 gnd C_bl
Cbb_26_53 bitb_26_53 gnd C_bl
Rb_26_54 bit_26_54 bit_26_55 R_bl
Rbb_26_54 bitb_26_54 bitb_26_55 R_bl
Cb_26_54 bit_26_54 gnd C_bl
Cbb_26_54 bitb_26_54 gnd C_bl
Rb_26_55 bit_26_55 bit_26_56 R_bl
Rbb_26_55 bitb_26_55 bitb_26_56 R_bl
Cb_26_55 bit_26_55 gnd C_bl
Cbb_26_55 bitb_26_55 gnd C_bl
Rb_26_56 bit_26_56 bit_26_57 R_bl
Rbb_26_56 bitb_26_56 bitb_26_57 R_bl
Cb_26_56 bit_26_56 gnd C_bl
Cbb_26_56 bitb_26_56 gnd C_bl
Rb_26_57 bit_26_57 bit_26_58 R_bl
Rbb_26_57 bitb_26_57 bitb_26_58 R_bl
Cb_26_57 bit_26_57 gnd C_bl
Cbb_26_57 bitb_26_57 gnd C_bl
Rb_26_58 bit_26_58 bit_26_59 R_bl
Rbb_26_58 bitb_26_58 bitb_26_59 R_bl
Cb_26_58 bit_26_58 gnd C_bl
Cbb_26_58 bitb_26_58 gnd C_bl
Rb_26_59 bit_26_59 bit_26_60 R_bl
Rbb_26_59 bitb_26_59 bitb_26_60 R_bl
Cb_26_59 bit_26_59 gnd C_bl
Cbb_26_59 bitb_26_59 gnd C_bl
Rb_26_60 bit_26_60 bit_26_61 R_bl
Rbb_26_60 bitb_26_60 bitb_26_61 R_bl
Cb_26_60 bit_26_60 gnd C_bl
Cbb_26_60 bitb_26_60 gnd C_bl
Rb_26_61 bit_26_61 bit_26_62 R_bl
Rbb_26_61 bitb_26_61 bitb_26_62 R_bl
Cb_26_61 bit_26_61 gnd C_bl
Cbb_26_61 bitb_26_61 gnd C_bl
Rb_26_62 bit_26_62 bit_26_63 R_bl
Rbb_26_62 bitb_26_62 bitb_26_63 R_bl
Cb_26_62 bit_26_62 gnd C_bl
Cbb_26_62 bitb_26_62 gnd C_bl
Rb_26_63 bit_26_63 bit_26_64 R_bl
Rbb_26_63 bitb_26_63 bitb_26_64 R_bl
Cb_26_63 bit_26_63 gnd C_bl
Cbb_26_63 bitb_26_63 gnd C_bl
Rb_26_64 bit_26_64 bit_26_65 R_bl
Rbb_26_64 bitb_26_64 bitb_26_65 R_bl
Cb_26_64 bit_26_64 gnd C_bl
Cbb_26_64 bitb_26_64 gnd C_bl
Rb_26_65 bit_26_65 bit_26_66 R_bl
Rbb_26_65 bitb_26_65 bitb_26_66 R_bl
Cb_26_65 bit_26_65 gnd C_bl
Cbb_26_65 bitb_26_65 gnd C_bl
Rb_26_66 bit_26_66 bit_26_67 R_bl
Rbb_26_66 bitb_26_66 bitb_26_67 R_bl
Cb_26_66 bit_26_66 gnd C_bl
Cbb_26_66 bitb_26_66 gnd C_bl
Rb_26_67 bit_26_67 bit_26_68 R_bl
Rbb_26_67 bitb_26_67 bitb_26_68 R_bl
Cb_26_67 bit_26_67 gnd C_bl
Cbb_26_67 bitb_26_67 gnd C_bl
Rb_26_68 bit_26_68 bit_26_69 R_bl
Rbb_26_68 bitb_26_68 bitb_26_69 R_bl
Cb_26_68 bit_26_68 gnd C_bl
Cbb_26_68 bitb_26_68 gnd C_bl
Rb_26_69 bit_26_69 bit_26_70 R_bl
Rbb_26_69 bitb_26_69 bitb_26_70 R_bl
Cb_26_69 bit_26_69 gnd C_bl
Cbb_26_69 bitb_26_69 gnd C_bl
Rb_26_70 bit_26_70 bit_26_71 R_bl
Rbb_26_70 bitb_26_70 bitb_26_71 R_bl
Cb_26_70 bit_26_70 gnd C_bl
Cbb_26_70 bitb_26_70 gnd C_bl
Rb_26_71 bit_26_71 bit_26_72 R_bl
Rbb_26_71 bitb_26_71 bitb_26_72 R_bl
Cb_26_71 bit_26_71 gnd C_bl
Cbb_26_71 bitb_26_71 gnd C_bl
Rb_26_72 bit_26_72 bit_26_73 R_bl
Rbb_26_72 bitb_26_72 bitb_26_73 R_bl
Cb_26_72 bit_26_72 gnd C_bl
Cbb_26_72 bitb_26_72 gnd C_bl
Rb_26_73 bit_26_73 bit_26_74 R_bl
Rbb_26_73 bitb_26_73 bitb_26_74 R_bl
Cb_26_73 bit_26_73 gnd C_bl
Cbb_26_73 bitb_26_73 gnd C_bl
Rb_26_74 bit_26_74 bit_26_75 R_bl
Rbb_26_74 bitb_26_74 bitb_26_75 R_bl
Cb_26_74 bit_26_74 gnd C_bl
Cbb_26_74 bitb_26_74 gnd C_bl
Rb_26_75 bit_26_75 bit_26_76 R_bl
Rbb_26_75 bitb_26_75 bitb_26_76 R_bl
Cb_26_75 bit_26_75 gnd C_bl
Cbb_26_75 bitb_26_75 gnd C_bl
Rb_26_76 bit_26_76 bit_26_77 R_bl
Rbb_26_76 bitb_26_76 bitb_26_77 R_bl
Cb_26_76 bit_26_76 gnd C_bl
Cbb_26_76 bitb_26_76 gnd C_bl
Rb_26_77 bit_26_77 bit_26_78 R_bl
Rbb_26_77 bitb_26_77 bitb_26_78 R_bl
Cb_26_77 bit_26_77 gnd C_bl
Cbb_26_77 bitb_26_77 gnd C_bl
Rb_26_78 bit_26_78 bit_26_79 R_bl
Rbb_26_78 bitb_26_78 bitb_26_79 R_bl
Cb_26_78 bit_26_78 gnd C_bl
Cbb_26_78 bitb_26_78 gnd C_bl
Rb_26_79 bit_26_79 bit_26_80 R_bl
Rbb_26_79 bitb_26_79 bitb_26_80 R_bl
Cb_26_79 bit_26_79 gnd C_bl
Cbb_26_79 bitb_26_79 gnd C_bl
Rb_26_80 bit_26_80 bit_26_81 R_bl
Rbb_26_80 bitb_26_80 bitb_26_81 R_bl
Cb_26_80 bit_26_80 gnd C_bl
Cbb_26_80 bitb_26_80 gnd C_bl
Rb_26_81 bit_26_81 bit_26_82 R_bl
Rbb_26_81 bitb_26_81 bitb_26_82 R_bl
Cb_26_81 bit_26_81 gnd C_bl
Cbb_26_81 bitb_26_81 gnd C_bl
Rb_26_82 bit_26_82 bit_26_83 R_bl
Rbb_26_82 bitb_26_82 bitb_26_83 R_bl
Cb_26_82 bit_26_82 gnd C_bl
Cbb_26_82 bitb_26_82 gnd C_bl
Rb_26_83 bit_26_83 bit_26_84 R_bl
Rbb_26_83 bitb_26_83 bitb_26_84 R_bl
Cb_26_83 bit_26_83 gnd C_bl
Cbb_26_83 bitb_26_83 gnd C_bl
Rb_26_84 bit_26_84 bit_26_85 R_bl
Rbb_26_84 bitb_26_84 bitb_26_85 R_bl
Cb_26_84 bit_26_84 gnd C_bl
Cbb_26_84 bitb_26_84 gnd C_bl
Rb_26_85 bit_26_85 bit_26_86 R_bl
Rbb_26_85 bitb_26_85 bitb_26_86 R_bl
Cb_26_85 bit_26_85 gnd C_bl
Cbb_26_85 bitb_26_85 gnd C_bl
Rb_26_86 bit_26_86 bit_26_87 R_bl
Rbb_26_86 bitb_26_86 bitb_26_87 R_bl
Cb_26_86 bit_26_86 gnd C_bl
Cbb_26_86 bitb_26_86 gnd C_bl
Rb_26_87 bit_26_87 bit_26_88 R_bl
Rbb_26_87 bitb_26_87 bitb_26_88 R_bl
Cb_26_87 bit_26_87 gnd C_bl
Cbb_26_87 bitb_26_87 gnd C_bl
Rb_26_88 bit_26_88 bit_26_89 R_bl
Rbb_26_88 bitb_26_88 bitb_26_89 R_bl
Cb_26_88 bit_26_88 gnd C_bl
Cbb_26_88 bitb_26_88 gnd C_bl
Rb_26_89 bit_26_89 bit_26_90 R_bl
Rbb_26_89 bitb_26_89 bitb_26_90 R_bl
Cb_26_89 bit_26_89 gnd C_bl
Cbb_26_89 bitb_26_89 gnd C_bl
Rb_26_90 bit_26_90 bit_26_91 R_bl
Rbb_26_90 bitb_26_90 bitb_26_91 R_bl
Cb_26_90 bit_26_90 gnd C_bl
Cbb_26_90 bitb_26_90 gnd C_bl
Rb_26_91 bit_26_91 bit_26_92 R_bl
Rbb_26_91 bitb_26_91 bitb_26_92 R_bl
Cb_26_91 bit_26_91 gnd C_bl
Cbb_26_91 bitb_26_91 gnd C_bl
Rb_26_92 bit_26_92 bit_26_93 R_bl
Rbb_26_92 bitb_26_92 bitb_26_93 R_bl
Cb_26_92 bit_26_92 gnd C_bl
Cbb_26_92 bitb_26_92 gnd C_bl
Rb_26_93 bit_26_93 bit_26_94 R_bl
Rbb_26_93 bitb_26_93 bitb_26_94 R_bl
Cb_26_93 bit_26_93 gnd C_bl
Cbb_26_93 bitb_26_93 gnd C_bl
Rb_26_94 bit_26_94 bit_26_95 R_bl
Rbb_26_94 bitb_26_94 bitb_26_95 R_bl
Cb_26_94 bit_26_94 gnd C_bl
Cbb_26_94 bitb_26_94 gnd C_bl
Rb_26_95 bit_26_95 bit_26_96 R_bl
Rbb_26_95 bitb_26_95 bitb_26_96 R_bl
Cb_26_95 bit_26_95 gnd C_bl
Cbb_26_95 bitb_26_95 gnd C_bl
Rb_26_96 bit_26_96 bit_26_97 R_bl
Rbb_26_96 bitb_26_96 bitb_26_97 R_bl
Cb_26_96 bit_26_96 gnd C_bl
Cbb_26_96 bitb_26_96 gnd C_bl
Rb_26_97 bit_26_97 bit_26_98 R_bl
Rbb_26_97 bitb_26_97 bitb_26_98 R_bl
Cb_26_97 bit_26_97 gnd C_bl
Cbb_26_97 bitb_26_97 gnd C_bl
Rb_26_98 bit_26_98 bit_26_99 R_bl
Rbb_26_98 bitb_26_98 bitb_26_99 R_bl
Cb_26_98 bit_26_98 gnd C_bl
Cbb_26_98 bitb_26_98 gnd C_bl
Rb_26_99 bit_26_99 bit_26_100 R_bl
Rbb_26_99 bitb_26_99 bitb_26_100 R_bl
Cb_26_99 bit_26_99 gnd C_bl
Cbb_26_99 bitb_26_99 gnd C_bl
Rb_27_0 bit_27_0 bit_27_1 R_bl
Rbb_27_0 bitb_27_0 bitb_27_1 R_bl
Cb_27_0 bit_27_0 gnd C_bl
Cbb_27_0 bitb_27_0 gnd C_bl
Rb_27_1 bit_27_1 bit_27_2 R_bl
Rbb_27_1 bitb_27_1 bitb_27_2 R_bl
Cb_27_1 bit_27_1 gnd C_bl
Cbb_27_1 bitb_27_1 gnd C_bl
Rb_27_2 bit_27_2 bit_27_3 R_bl
Rbb_27_2 bitb_27_2 bitb_27_3 R_bl
Cb_27_2 bit_27_2 gnd C_bl
Cbb_27_2 bitb_27_2 gnd C_bl
Rb_27_3 bit_27_3 bit_27_4 R_bl
Rbb_27_3 bitb_27_3 bitb_27_4 R_bl
Cb_27_3 bit_27_3 gnd C_bl
Cbb_27_3 bitb_27_3 gnd C_bl
Rb_27_4 bit_27_4 bit_27_5 R_bl
Rbb_27_4 bitb_27_4 bitb_27_5 R_bl
Cb_27_4 bit_27_4 gnd C_bl
Cbb_27_4 bitb_27_4 gnd C_bl
Rb_27_5 bit_27_5 bit_27_6 R_bl
Rbb_27_5 bitb_27_5 bitb_27_6 R_bl
Cb_27_5 bit_27_5 gnd C_bl
Cbb_27_5 bitb_27_5 gnd C_bl
Rb_27_6 bit_27_6 bit_27_7 R_bl
Rbb_27_6 bitb_27_6 bitb_27_7 R_bl
Cb_27_6 bit_27_6 gnd C_bl
Cbb_27_6 bitb_27_6 gnd C_bl
Rb_27_7 bit_27_7 bit_27_8 R_bl
Rbb_27_7 bitb_27_7 bitb_27_8 R_bl
Cb_27_7 bit_27_7 gnd C_bl
Cbb_27_7 bitb_27_7 gnd C_bl
Rb_27_8 bit_27_8 bit_27_9 R_bl
Rbb_27_8 bitb_27_8 bitb_27_9 R_bl
Cb_27_8 bit_27_8 gnd C_bl
Cbb_27_8 bitb_27_8 gnd C_bl
Rb_27_9 bit_27_9 bit_27_10 R_bl
Rbb_27_9 bitb_27_9 bitb_27_10 R_bl
Cb_27_9 bit_27_9 gnd C_bl
Cbb_27_9 bitb_27_9 gnd C_bl
Rb_27_10 bit_27_10 bit_27_11 R_bl
Rbb_27_10 bitb_27_10 bitb_27_11 R_bl
Cb_27_10 bit_27_10 gnd C_bl
Cbb_27_10 bitb_27_10 gnd C_bl
Rb_27_11 bit_27_11 bit_27_12 R_bl
Rbb_27_11 bitb_27_11 bitb_27_12 R_bl
Cb_27_11 bit_27_11 gnd C_bl
Cbb_27_11 bitb_27_11 gnd C_bl
Rb_27_12 bit_27_12 bit_27_13 R_bl
Rbb_27_12 bitb_27_12 bitb_27_13 R_bl
Cb_27_12 bit_27_12 gnd C_bl
Cbb_27_12 bitb_27_12 gnd C_bl
Rb_27_13 bit_27_13 bit_27_14 R_bl
Rbb_27_13 bitb_27_13 bitb_27_14 R_bl
Cb_27_13 bit_27_13 gnd C_bl
Cbb_27_13 bitb_27_13 gnd C_bl
Rb_27_14 bit_27_14 bit_27_15 R_bl
Rbb_27_14 bitb_27_14 bitb_27_15 R_bl
Cb_27_14 bit_27_14 gnd C_bl
Cbb_27_14 bitb_27_14 gnd C_bl
Rb_27_15 bit_27_15 bit_27_16 R_bl
Rbb_27_15 bitb_27_15 bitb_27_16 R_bl
Cb_27_15 bit_27_15 gnd C_bl
Cbb_27_15 bitb_27_15 gnd C_bl
Rb_27_16 bit_27_16 bit_27_17 R_bl
Rbb_27_16 bitb_27_16 bitb_27_17 R_bl
Cb_27_16 bit_27_16 gnd C_bl
Cbb_27_16 bitb_27_16 gnd C_bl
Rb_27_17 bit_27_17 bit_27_18 R_bl
Rbb_27_17 bitb_27_17 bitb_27_18 R_bl
Cb_27_17 bit_27_17 gnd C_bl
Cbb_27_17 bitb_27_17 gnd C_bl
Rb_27_18 bit_27_18 bit_27_19 R_bl
Rbb_27_18 bitb_27_18 bitb_27_19 R_bl
Cb_27_18 bit_27_18 gnd C_bl
Cbb_27_18 bitb_27_18 gnd C_bl
Rb_27_19 bit_27_19 bit_27_20 R_bl
Rbb_27_19 bitb_27_19 bitb_27_20 R_bl
Cb_27_19 bit_27_19 gnd C_bl
Cbb_27_19 bitb_27_19 gnd C_bl
Rb_27_20 bit_27_20 bit_27_21 R_bl
Rbb_27_20 bitb_27_20 bitb_27_21 R_bl
Cb_27_20 bit_27_20 gnd C_bl
Cbb_27_20 bitb_27_20 gnd C_bl
Rb_27_21 bit_27_21 bit_27_22 R_bl
Rbb_27_21 bitb_27_21 bitb_27_22 R_bl
Cb_27_21 bit_27_21 gnd C_bl
Cbb_27_21 bitb_27_21 gnd C_bl
Rb_27_22 bit_27_22 bit_27_23 R_bl
Rbb_27_22 bitb_27_22 bitb_27_23 R_bl
Cb_27_22 bit_27_22 gnd C_bl
Cbb_27_22 bitb_27_22 gnd C_bl
Rb_27_23 bit_27_23 bit_27_24 R_bl
Rbb_27_23 bitb_27_23 bitb_27_24 R_bl
Cb_27_23 bit_27_23 gnd C_bl
Cbb_27_23 bitb_27_23 gnd C_bl
Rb_27_24 bit_27_24 bit_27_25 R_bl
Rbb_27_24 bitb_27_24 bitb_27_25 R_bl
Cb_27_24 bit_27_24 gnd C_bl
Cbb_27_24 bitb_27_24 gnd C_bl
Rb_27_25 bit_27_25 bit_27_26 R_bl
Rbb_27_25 bitb_27_25 bitb_27_26 R_bl
Cb_27_25 bit_27_25 gnd C_bl
Cbb_27_25 bitb_27_25 gnd C_bl
Rb_27_26 bit_27_26 bit_27_27 R_bl
Rbb_27_26 bitb_27_26 bitb_27_27 R_bl
Cb_27_26 bit_27_26 gnd C_bl
Cbb_27_26 bitb_27_26 gnd C_bl
Rb_27_27 bit_27_27 bit_27_28 R_bl
Rbb_27_27 bitb_27_27 bitb_27_28 R_bl
Cb_27_27 bit_27_27 gnd C_bl
Cbb_27_27 bitb_27_27 gnd C_bl
Rb_27_28 bit_27_28 bit_27_29 R_bl
Rbb_27_28 bitb_27_28 bitb_27_29 R_bl
Cb_27_28 bit_27_28 gnd C_bl
Cbb_27_28 bitb_27_28 gnd C_bl
Rb_27_29 bit_27_29 bit_27_30 R_bl
Rbb_27_29 bitb_27_29 bitb_27_30 R_bl
Cb_27_29 bit_27_29 gnd C_bl
Cbb_27_29 bitb_27_29 gnd C_bl
Rb_27_30 bit_27_30 bit_27_31 R_bl
Rbb_27_30 bitb_27_30 bitb_27_31 R_bl
Cb_27_30 bit_27_30 gnd C_bl
Cbb_27_30 bitb_27_30 gnd C_bl
Rb_27_31 bit_27_31 bit_27_32 R_bl
Rbb_27_31 bitb_27_31 bitb_27_32 R_bl
Cb_27_31 bit_27_31 gnd C_bl
Cbb_27_31 bitb_27_31 gnd C_bl
Rb_27_32 bit_27_32 bit_27_33 R_bl
Rbb_27_32 bitb_27_32 bitb_27_33 R_bl
Cb_27_32 bit_27_32 gnd C_bl
Cbb_27_32 bitb_27_32 gnd C_bl
Rb_27_33 bit_27_33 bit_27_34 R_bl
Rbb_27_33 bitb_27_33 bitb_27_34 R_bl
Cb_27_33 bit_27_33 gnd C_bl
Cbb_27_33 bitb_27_33 gnd C_bl
Rb_27_34 bit_27_34 bit_27_35 R_bl
Rbb_27_34 bitb_27_34 bitb_27_35 R_bl
Cb_27_34 bit_27_34 gnd C_bl
Cbb_27_34 bitb_27_34 gnd C_bl
Rb_27_35 bit_27_35 bit_27_36 R_bl
Rbb_27_35 bitb_27_35 bitb_27_36 R_bl
Cb_27_35 bit_27_35 gnd C_bl
Cbb_27_35 bitb_27_35 gnd C_bl
Rb_27_36 bit_27_36 bit_27_37 R_bl
Rbb_27_36 bitb_27_36 bitb_27_37 R_bl
Cb_27_36 bit_27_36 gnd C_bl
Cbb_27_36 bitb_27_36 gnd C_bl
Rb_27_37 bit_27_37 bit_27_38 R_bl
Rbb_27_37 bitb_27_37 bitb_27_38 R_bl
Cb_27_37 bit_27_37 gnd C_bl
Cbb_27_37 bitb_27_37 gnd C_bl
Rb_27_38 bit_27_38 bit_27_39 R_bl
Rbb_27_38 bitb_27_38 bitb_27_39 R_bl
Cb_27_38 bit_27_38 gnd C_bl
Cbb_27_38 bitb_27_38 gnd C_bl
Rb_27_39 bit_27_39 bit_27_40 R_bl
Rbb_27_39 bitb_27_39 bitb_27_40 R_bl
Cb_27_39 bit_27_39 gnd C_bl
Cbb_27_39 bitb_27_39 gnd C_bl
Rb_27_40 bit_27_40 bit_27_41 R_bl
Rbb_27_40 bitb_27_40 bitb_27_41 R_bl
Cb_27_40 bit_27_40 gnd C_bl
Cbb_27_40 bitb_27_40 gnd C_bl
Rb_27_41 bit_27_41 bit_27_42 R_bl
Rbb_27_41 bitb_27_41 bitb_27_42 R_bl
Cb_27_41 bit_27_41 gnd C_bl
Cbb_27_41 bitb_27_41 gnd C_bl
Rb_27_42 bit_27_42 bit_27_43 R_bl
Rbb_27_42 bitb_27_42 bitb_27_43 R_bl
Cb_27_42 bit_27_42 gnd C_bl
Cbb_27_42 bitb_27_42 gnd C_bl
Rb_27_43 bit_27_43 bit_27_44 R_bl
Rbb_27_43 bitb_27_43 bitb_27_44 R_bl
Cb_27_43 bit_27_43 gnd C_bl
Cbb_27_43 bitb_27_43 gnd C_bl
Rb_27_44 bit_27_44 bit_27_45 R_bl
Rbb_27_44 bitb_27_44 bitb_27_45 R_bl
Cb_27_44 bit_27_44 gnd C_bl
Cbb_27_44 bitb_27_44 gnd C_bl
Rb_27_45 bit_27_45 bit_27_46 R_bl
Rbb_27_45 bitb_27_45 bitb_27_46 R_bl
Cb_27_45 bit_27_45 gnd C_bl
Cbb_27_45 bitb_27_45 gnd C_bl
Rb_27_46 bit_27_46 bit_27_47 R_bl
Rbb_27_46 bitb_27_46 bitb_27_47 R_bl
Cb_27_46 bit_27_46 gnd C_bl
Cbb_27_46 bitb_27_46 gnd C_bl
Rb_27_47 bit_27_47 bit_27_48 R_bl
Rbb_27_47 bitb_27_47 bitb_27_48 R_bl
Cb_27_47 bit_27_47 gnd C_bl
Cbb_27_47 bitb_27_47 gnd C_bl
Rb_27_48 bit_27_48 bit_27_49 R_bl
Rbb_27_48 bitb_27_48 bitb_27_49 R_bl
Cb_27_48 bit_27_48 gnd C_bl
Cbb_27_48 bitb_27_48 gnd C_bl
Rb_27_49 bit_27_49 bit_27_50 R_bl
Rbb_27_49 bitb_27_49 bitb_27_50 R_bl
Cb_27_49 bit_27_49 gnd C_bl
Cbb_27_49 bitb_27_49 gnd C_bl
Rb_27_50 bit_27_50 bit_27_51 R_bl
Rbb_27_50 bitb_27_50 bitb_27_51 R_bl
Cb_27_50 bit_27_50 gnd C_bl
Cbb_27_50 bitb_27_50 gnd C_bl
Rb_27_51 bit_27_51 bit_27_52 R_bl
Rbb_27_51 bitb_27_51 bitb_27_52 R_bl
Cb_27_51 bit_27_51 gnd C_bl
Cbb_27_51 bitb_27_51 gnd C_bl
Rb_27_52 bit_27_52 bit_27_53 R_bl
Rbb_27_52 bitb_27_52 bitb_27_53 R_bl
Cb_27_52 bit_27_52 gnd C_bl
Cbb_27_52 bitb_27_52 gnd C_bl
Rb_27_53 bit_27_53 bit_27_54 R_bl
Rbb_27_53 bitb_27_53 bitb_27_54 R_bl
Cb_27_53 bit_27_53 gnd C_bl
Cbb_27_53 bitb_27_53 gnd C_bl
Rb_27_54 bit_27_54 bit_27_55 R_bl
Rbb_27_54 bitb_27_54 bitb_27_55 R_bl
Cb_27_54 bit_27_54 gnd C_bl
Cbb_27_54 bitb_27_54 gnd C_bl
Rb_27_55 bit_27_55 bit_27_56 R_bl
Rbb_27_55 bitb_27_55 bitb_27_56 R_bl
Cb_27_55 bit_27_55 gnd C_bl
Cbb_27_55 bitb_27_55 gnd C_bl
Rb_27_56 bit_27_56 bit_27_57 R_bl
Rbb_27_56 bitb_27_56 bitb_27_57 R_bl
Cb_27_56 bit_27_56 gnd C_bl
Cbb_27_56 bitb_27_56 gnd C_bl
Rb_27_57 bit_27_57 bit_27_58 R_bl
Rbb_27_57 bitb_27_57 bitb_27_58 R_bl
Cb_27_57 bit_27_57 gnd C_bl
Cbb_27_57 bitb_27_57 gnd C_bl
Rb_27_58 bit_27_58 bit_27_59 R_bl
Rbb_27_58 bitb_27_58 bitb_27_59 R_bl
Cb_27_58 bit_27_58 gnd C_bl
Cbb_27_58 bitb_27_58 gnd C_bl
Rb_27_59 bit_27_59 bit_27_60 R_bl
Rbb_27_59 bitb_27_59 bitb_27_60 R_bl
Cb_27_59 bit_27_59 gnd C_bl
Cbb_27_59 bitb_27_59 gnd C_bl
Rb_27_60 bit_27_60 bit_27_61 R_bl
Rbb_27_60 bitb_27_60 bitb_27_61 R_bl
Cb_27_60 bit_27_60 gnd C_bl
Cbb_27_60 bitb_27_60 gnd C_bl
Rb_27_61 bit_27_61 bit_27_62 R_bl
Rbb_27_61 bitb_27_61 bitb_27_62 R_bl
Cb_27_61 bit_27_61 gnd C_bl
Cbb_27_61 bitb_27_61 gnd C_bl
Rb_27_62 bit_27_62 bit_27_63 R_bl
Rbb_27_62 bitb_27_62 bitb_27_63 R_bl
Cb_27_62 bit_27_62 gnd C_bl
Cbb_27_62 bitb_27_62 gnd C_bl
Rb_27_63 bit_27_63 bit_27_64 R_bl
Rbb_27_63 bitb_27_63 bitb_27_64 R_bl
Cb_27_63 bit_27_63 gnd C_bl
Cbb_27_63 bitb_27_63 gnd C_bl
Rb_27_64 bit_27_64 bit_27_65 R_bl
Rbb_27_64 bitb_27_64 bitb_27_65 R_bl
Cb_27_64 bit_27_64 gnd C_bl
Cbb_27_64 bitb_27_64 gnd C_bl
Rb_27_65 bit_27_65 bit_27_66 R_bl
Rbb_27_65 bitb_27_65 bitb_27_66 R_bl
Cb_27_65 bit_27_65 gnd C_bl
Cbb_27_65 bitb_27_65 gnd C_bl
Rb_27_66 bit_27_66 bit_27_67 R_bl
Rbb_27_66 bitb_27_66 bitb_27_67 R_bl
Cb_27_66 bit_27_66 gnd C_bl
Cbb_27_66 bitb_27_66 gnd C_bl
Rb_27_67 bit_27_67 bit_27_68 R_bl
Rbb_27_67 bitb_27_67 bitb_27_68 R_bl
Cb_27_67 bit_27_67 gnd C_bl
Cbb_27_67 bitb_27_67 gnd C_bl
Rb_27_68 bit_27_68 bit_27_69 R_bl
Rbb_27_68 bitb_27_68 bitb_27_69 R_bl
Cb_27_68 bit_27_68 gnd C_bl
Cbb_27_68 bitb_27_68 gnd C_bl
Rb_27_69 bit_27_69 bit_27_70 R_bl
Rbb_27_69 bitb_27_69 bitb_27_70 R_bl
Cb_27_69 bit_27_69 gnd C_bl
Cbb_27_69 bitb_27_69 gnd C_bl
Rb_27_70 bit_27_70 bit_27_71 R_bl
Rbb_27_70 bitb_27_70 bitb_27_71 R_bl
Cb_27_70 bit_27_70 gnd C_bl
Cbb_27_70 bitb_27_70 gnd C_bl
Rb_27_71 bit_27_71 bit_27_72 R_bl
Rbb_27_71 bitb_27_71 bitb_27_72 R_bl
Cb_27_71 bit_27_71 gnd C_bl
Cbb_27_71 bitb_27_71 gnd C_bl
Rb_27_72 bit_27_72 bit_27_73 R_bl
Rbb_27_72 bitb_27_72 bitb_27_73 R_bl
Cb_27_72 bit_27_72 gnd C_bl
Cbb_27_72 bitb_27_72 gnd C_bl
Rb_27_73 bit_27_73 bit_27_74 R_bl
Rbb_27_73 bitb_27_73 bitb_27_74 R_bl
Cb_27_73 bit_27_73 gnd C_bl
Cbb_27_73 bitb_27_73 gnd C_bl
Rb_27_74 bit_27_74 bit_27_75 R_bl
Rbb_27_74 bitb_27_74 bitb_27_75 R_bl
Cb_27_74 bit_27_74 gnd C_bl
Cbb_27_74 bitb_27_74 gnd C_bl
Rb_27_75 bit_27_75 bit_27_76 R_bl
Rbb_27_75 bitb_27_75 bitb_27_76 R_bl
Cb_27_75 bit_27_75 gnd C_bl
Cbb_27_75 bitb_27_75 gnd C_bl
Rb_27_76 bit_27_76 bit_27_77 R_bl
Rbb_27_76 bitb_27_76 bitb_27_77 R_bl
Cb_27_76 bit_27_76 gnd C_bl
Cbb_27_76 bitb_27_76 gnd C_bl
Rb_27_77 bit_27_77 bit_27_78 R_bl
Rbb_27_77 bitb_27_77 bitb_27_78 R_bl
Cb_27_77 bit_27_77 gnd C_bl
Cbb_27_77 bitb_27_77 gnd C_bl
Rb_27_78 bit_27_78 bit_27_79 R_bl
Rbb_27_78 bitb_27_78 bitb_27_79 R_bl
Cb_27_78 bit_27_78 gnd C_bl
Cbb_27_78 bitb_27_78 gnd C_bl
Rb_27_79 bit_27_79 bit_27_80 R_bl
Rbb_27_79 bitb_27_79 bitb_27_80 R_bl
Cb_27_79 bit_27_79 gnd C_bl
Cbb_27_79 bitb_27_79 gnd C_bl
Rb_27_80 bit_27_80 bit_27_81 R_bl
Rbb_27_80 bitb_27_80 bitb_27_81 R_bl
Cb_27_80 bit_27_80 gnd C_bl
Cbb_27_80 bitb_27_80 gnd C_bl
Rb_27_81 bit_27_81 bit_27_82 R_bl
Rbb_27_81 bitb_27_81 bitb_27_82 R_bl
Cb_27_81 bit_27_81 gnd C_bl
Cbb_27_81 bitb_27_81 gnd C_bl
Rb_27_82 bit_27_82 bit_27_83 R_bl
Rbb_27_82 bitb_27_82 bitb_27_83 R_bl
Cb_27_82 bit_27_82 gnd C_bl
Cbb_27_82 bitb_27_82 gnd C_bl
Rb_27_83 bit_27_83 bit_27_84 R_bl
Rbb_27_83 bitb_27_83 bitb_27_84 R_bl
Cb_27_83 bit_27_83 gnd C_bl
Cbb_27_83 bitb_27_83 gnd C_bl
Rb_27_84 bit_27_84 bit_27_85 R_bl
Rbb_27_84 bitb_27_84 bitb_27_85 R_bl
Cb_27_84 bit_27_84 gnd C_bl
Cbb_27_84 bitb_27_84 gnd C_bl
Rb_27_85 bit_27_85 bit_27_86 R_bl
Rbb_27_85 bitb_27_85 bitb_27_86 R_bl
Cb_27_85 bit_27_85 gnd C_bl
Cbb_27_85 bitb_27_85 gnd C_bl
Rb_27_86 bit_27_86 bit_27_87 R_bl
Rbb_27_86 bitb_27_86 bitb_27_87 R_bl
Cb_27_86 bit_27_86 gnd C_bl
Cbb_27_86 bitb_27_86 gnd C_bl
Rb_27_87 bit_27_87 bit_27_88 R_bl
Rbb_27_87 bitb_27_87 bitb_27_88 R_bl
Cb_27_87 bit_27_87 gnd C_bl
Cbb_27_87 bitb_27_87 gnd C_bl
Rb_27_88 bit_27_88 bit_27_89 R_bl
Rbb_27_88 bitb_27_88 bitb_27_89 R_bl
Cb_27_88 bit_27_88 gnd C_bl
Cbb_27_88 bitb_27_88 gnd C_bl
Rb_27_89 bit_27_89 bit_27_90 R_bl
Rbb_27_89 bitb_27_89 bitb_27_90 R_bl
Cb_27_89 bit_27_89 gnd C_bl
Cbb_27_89 bitb_27_89 gnd C_bl
Rb_27_90 bit_27_90 bit_27_91 R_bl
Rbb_27_90 bitb_27_90 bitb_27_91 R_bl
Cb_27_90 bit_27_90 gnd C_bl
Cbb_27_90 bitb_27_90 gnd C_bl
Rb_27_91 bit_27_91 bit_27_92 R_bl
Rbb_27_91 bitb_27_91 bitb_27_92 R_bl
Cb_27_91 bit_27_91 gnd C_bl
Cbb_27_91 bitb_27_91 gnd C_bl
Rb_27_92 bit_27_92 bit_27_93 R_bl
Rbb_27_92 bitb_27_92 bitb_27_93 R_bl
Cb_27_92 bit_27_92 gnd C_bl
Cbb_27_92 bitb_27_92 gnd C_bl
Rb_27_93 bit_27_93 bit_27_94 R_bl
Rbb_27_93 bitb_27_93 bitb_27_94 R_bl
Cb_27_93 bit_27_93 gnd C_bl
Cbb_27_93 bitb_27_93 gnd C_bl
Rb_27_94 bit_27_94 bit_27_95 R_bl
Rbb_27_94 bitb_27_94 bitb_27_95 R_bl
Cb_27_94 bit_27_94 gnd C_bl
Cbb_27_94 bitb_27_94 gnd C_bl
Rb_27_95 bit_27_95 bit_27_96 R_bl
Rbb_27_95 bitb_27_95 bitb_27_96 R_bl
Cb_27_95 bit_27_95 gnd C_bl
Cbb_27_95 bitb_27_95 gnd C_bl
Rb_27_96 bit_27_96 bit_27_97 R_bl
Rbb_27_96 bitb_27_96 bitb_27_97 R_bl
Cb_27_96 bit_27_96 gnd C_bl
Cbb_27_96 bitb_27_96 gnd C_bl
Rb_27_97 bit_27_97 bit_27_98 R_bl
Rbb_27_97 bitb_27_97 bitb_27_98 R_bl
Cb_27_97 bit_27_97 gnd C_bl
Cbb_27_97 bitb_27_97 gnd C_bl
Rb_27_98 bit_27_98 bit_27_99 R_bl
Rbb_27_98 bitb_27_98 bitb_27_99 R_bl
Cb_27_98 bit_27_98 gnd C_bl
Cbb_27_98 bitb_27_98 gnd C_bl
Rb_27_99 bit_27_99 bit_27_100 R_bl
Rbb_27_99 bitb_27_99 bitb_27_100 R_bl
Cb_27_99 bit_27_99 gnd C_bl
Cbb_27_99 bitb_27_99 gnd C_bl
Rb_28_0 bit_28_0 bit_28_1 R_bl
Rbb_28_0 bitb_28_0 bitb_28_1 R_bl
Cb_28_0 bit_28_0 gnd C_bl
Cbb_28_0 bitb_28_0 gnd C_bl
Rb_28_1 bit_28_1 bit_28_2 R_bl
Rbb_28_1 bitb_28_1 bitb_28_2 R_bl
Cb_28_1 bit_28_1 gnd C_bl
Cbb_28_1 bitb_28_1 gnd C_bl
Rb_28_2 bit_28_2 bit_28_3 R_bl
Rbb_28_2 bitb_28_2 bitb_28_3 R_bl
Cb_28_2 bit_28_2 gnd C_bl
Cbb_28_2 bitb_28_2 gnd C_bl
Rb_28_3 bit_28_3 bit_28_4 R_bl
Rbb_28_3 bitb_28_3 bitb_28_4 R_bl
Cb_28_3 bit_28_3 gnd C_bl
Cbb_28_3 bitb_28_3 gnd C_bl
Rb_28_4 bit_28_4 bit_28_5 R_bl
Rbb_28_4 bitb_28_4 bitb_28_5 R_bl
Cb_28_4 bit_28_4 gnd C_bl
Cbb_28_4 bitb_28_4 gnd C_bl
Rb_28_5 bit_28_5 bit_28_6 R_bl
Rbb_28_5 bitb_28_5 bitb_28_6 R_bl
Cb_28_5 bit_28_5 gnd C_bl
Cbb_28_5 bitb_28_5 gnd C_bl
Rb_28_6 bit_28_6 bit_28_7 R_bl
Rbb_28_6 bitb_28_6 bitb_28_7 R_bl
Cb_28_6 bit_28_6 gnd C_bl
Cbb_28_6 bitb_28_6 gnd C_bl
Rb_28_7 bit_28_7 bit_28_8 R_bl
Rbb_28_7 bitb_28_7 bitb_28_8 R_bl
Cb_28_7 bit_28_7 gnd C_bl
Cbb_28_7 bitb_28_7 gnd C_bl
Rb_28_8 bit_28_8 bit_28_9 R_bl
Rbb_28_8 bitb_28_8 bitb_28_9 R_bl
Cb_28_8 bit_28_8 gnd C_bl
Cbb_28_8 bitb_28_8 gnd C_bl
Rb_28_9 bit_28_9 bit_28_10 R_bl
Rbb_28_9 bitb_28_9 bitb_28_10 R_bl
Cb_28_9 bit_28_9 gnd C_bl
Cbb_28_9 bitb_28_9 gnd C_bl
Rb_28_10 bit_28_10 bit_28_11 R_bl
Rbb_28_10 bitb_28_10 bitb_28_11 R_bl
Cb_28_10 bit_28_10 gnd C_bl
Cbb_28_10 bitb_28_10 gnd C_bl
Rb_28_11 bit_28_11 bit_28_12 R_bl
Rbb_28_11 bitb_28_11 bitb_28_12 R_bl
Cb_28_11 bit_28_11 gnd C_bl
Cbb_28_11 bitb_28_11 gnd C_bl
Rb_28_12 bit_28_12 bit_28_13 R_bl
Rbb_28_12 bitb_28_12 bitb_28_13 R_bl
Cb_28_12 bit_28_12 gnd C_bl
Cbb_28_12 bitb_28_12 gnd C_bl
Rb_28_13 bit_28_13 bit_28_14 R_bl
Rbb_28_13 bitb_28_13 bitb_28_14 R_bl
Cb_28_13 bit_28_13 gnd C_bl
Cbb_28_13 bitb_28_13 gnd C_bl
Rb_28_14 bit_28_14 bit_28_15 R_bl
Rbb_28_14 bitb_28_14 bitb_28_15 R_bl
Cb_28_14 bit_28_14 gnd C_bl
Cbb_28_14 bitb_28_14 gnd C_bl
Rb_28_15 bit_28_15 bit_28_16 R_bl
Rbb_28_15 bitb_28_15 bitb_28_16 R_bl
Cb_28_15 bit_28_15 gnd C_bl
Cbb_28_15 bitb_28_15 gnd C_bl
Rb_28_16 bit_28_16 bit_28_17 R_bl
Rbb_28_16 bitb_28_16 bitb_28_17 R_bl
Cb_28_16 bit_28_16 gnd C_bl
Cbb_28_16 bitb_28_16 gnd C_bl
Rb_28_17 bit_28_17 bit_28_18 R_bl
Rbb_28_17 bitb_28_17 bitb_28_18 R_bl
Cb_28_17 bit_28_17 gnd C_bl
Cbb_28_17 bitb_28_17 gnd C_bl
Rb_28_18 bit_28_18 bit_28_19 R_bl
Rbb_28_18 bitb_28_18 bitb_28_19 R_bl
Cb_28_18 bit_28_18 gnd C_bl
Cbb_28_18 bitb_28_18 gnd C_bl
Rb_28_19 bit_28_19 bit_28_20 R_bl
Rbb_28_19 bitb_28_19 bitb_28_20 R_bl
Cb_28_19 bit_28_19 gnd C_bl
Cbb_28_19 bitb_28_19 gnd C_bl
Rb_28_20 bit_28_20 bit_28_21 R_bl
Rbb_28_20 bitb_28_20 bitb_28_21 R_bl
Cb_28_20 bit_28_20 gnd C_bl
Cbb_28_20 bitb_28_20 gnd C_bl
Rb_28_21 bit_28_21 bit_28_22 R_bl
Rbb_28_21 bitb_28_21 bitb_28_22 R_bl
Cb_28_21 bit_28_21 gnd C_bl
Cbb_28_21 bitb_28_21 gnd C_bl
Rb_28_22 bit_28_22 bit_28_23 R_bl
Rbb_28_22 bitb_28_22 bitb_28_23 R_bl
Cb_28_22 bit_28_22 gnd C_bl
Cbb_28_22 bitb_28_22 gnd C_bl
Rb_28_23 bit_28_23 bit_28_24 R_bl
Rbb_28_23 bitb_28_23 bitb_28_24 R_bl
Cb_28_23 bit_28_23 gnd C_bl
Cbb_28_23 bitb_28_23 gnd C_bl
Rb_28_24 bit_28_24 bit_28_25 R_bl
Rbb_28_24 bitb_28_24 bitb_28_25 R_bl
Cb_28_24 bit_28_24 gnd C_bl
Cbb_28_24 bitb_28_24 gnd C_bl
Rb_28_25 bit_28_25 bit_28_26 R_bl
Rbb_28_25 bitb_28_25 bitb_28_26 R_bl
Cb_28_25 bit_28_25 gnd C_bl
Cbb_28_25 bitb_28_25 gnd C_bl
Rb_28_26 bit_28_26 bit_28_27 R_bl
Rbb_28_26 bitb_28_26 bitb_28_27 R_bl
Cb_28_26 bit_28_26 gnd C_bl
Cbb_28_26 bitb_28_26 gnd C_bl
Rb_28_27 bit_28_27 bit_28_28 R_bl
Rbb_28_27 bitb_28_27 bitb_28_28 R_bl
Cb_28_27 bit_28_27 gnd C_bl
Cbb_28_27 bitb_28_27 gnd C_bl
Rb_28_28 bit_28_28 bit_28_29 R_bl
Rbb_28_28 bitb_28_28 bitb_28_29 R_bl
Cb_28_28 bit_28_28 gnd C_bl
Cbb_28_28 bitb_28_28 gnd C_bl
Rb_28_29 bit_28_29 bit_28_30 R_bl
Rbb_28_29 bitb_28_29 bitb_28_30 R_bl
Cb_28_29 bit_28_29 gnd C_bl
Cbb_28_29 bitb_28_29 gnd C_bl
Rb_28_30 bit_28_30 bit_28_31 R_bl
Rbb_28_30 bitb_28_30 bitb_28_31 R_bl
Cb_28_30 bit_28_30 gnd C_bl
Cbb_28_30 bitb_28_30 gnd C_bl
Rb_28_31 bit_28_31 bit_28_32 R_bl
Rbb_28_31 bitb_28_31 bitb_28_32 R_bl
Cb_28_31 bit_28_31 gnd C_bl
Cbb_28_31 bitb_28_31 gnd C_bl
Rb_28_32 bit_28_32 bit_28_33 R_bl
Rbb_28_32 bitb_28_32 bitb_28_33 R_bl
Cb_28_32 bit_28_32 gnd C_bl
Cbb_28_32 bitb_28_32 gnd C_bl
Rb_28_33 bit_28_33 bit_28_34 R_bl
Rbb_28_33 bitb_28_33 bitb_28_34 R_bl
Cb_28_33 bit_28_33 gnd C_bl
Cbb_28_33 bitb_28_33 gnd C_bl
Rb_28_34 bit_28_34 bit_28_35 R_bl
Rbb_28_34 bitb_28_34 bitb_28_35 R_bl
Cb_28_34 bit_28_34 gnd C_bl
Cbb_28_34 bitb_28_34 gnd C_bl
Rb_28_35 bit_28_35 bit_28_36 R_bl
Rbb_28_35 bitb_28_35 bitb_28_36 R_bl
Cb_28_35 bit_28_35 gnd C_bl
Cbb_28_35 bitb_28_35 gnd C_bl
Rb_28_36 bit_28_36 bit_28_37 R_bl
Rbb_28_36 bitb_28_36 bitb_28_37 R_bl
Cb_28_36 bit_28_36 gnd C_bl
Cbb_28_36 bitb_28_36 gnd C_bl
Rb_28_37 bit_28_37 bit_28_38 R_bl
Rbb_28_37 bitb_28_37 bitb_28_38 R_bl
Cb_28_37 bit_28_37 gnd C_bl
Cbb_28_37 bitb_28_37 gnd C_bl
Rb_28_38 bit_28_38 bit_28_39 R_bl
Rbb_28_38 bitb_28_38 bitb_28_39 R_bl
Cb_28_38 bit_28_38 gnd C_bl
Cbb_28_38 bitb_28_38 gnd C_bl
Rb_28_39 bit_28_39 bit_28_40 R_bl
Rbb_28_39 bitb_28_39 bitb_28_40 R_bl
Cb_28_39 bit_28_39 gnd C_bl
Cbb_28_39 bitb_28_39 gnd C_bl
Rb_28_40 bit_28_40 bit_28_41 R_bl
Rbb_28_40 bitb_28_40 bitb_28_41 R_bl
Cb_28_40 bit_28_40 gnd C_bl
Cbb_28_40 bitb_28_40 gnd C_bl
Rb_28_41 bit_28_41 bit_28_42 R_bl
Rbb_28_41 bitb_28_41 bitb_28_42 R_bl
Cb_28_41 bit_28_41 gnd C_bl
Cbb_28_41 bitb_28_41 gnd C_bl
Rb_28_42 bit_28_42 bit_28_43 R_bl
Rbb_28_42 bitb_28_42 bitb_28_43 R_bl
Cb_28_42 bit_28_42 gnd C_bl
Cbb_28_42 bitb_28_42 gnd C_bl
Rb_28_43 bit_28_43 bit_28_44 R_bl
Rbb_28_43 bitb_28_43 bitb_28_44 R_bl
Cb_28_43 bit_28_43 gnd C_bl
Cbb_28_43 bitb_28_43 gnd C_bl
Rb_28_44 bit_28_44 bit_28_45 R_bl
Rbb_28_44 bitb_28_44 bitb_28_45 R_bl
Cb_28_44 bit_28_44 gnd C_bl
Cbb_28_44 bitb_28_44 gnd C_bl
Rb_28_45 bit_28_45 bit_28_46 R_bl
Rbb_28_45 bitb_28_45 bitb_28_46 R_bl
Cb_28_45 bit_28_45 gnd C_bl
Cbb_28_45 bitb_28_45 gnd C_bl
Rb_28_46 bit_28_46 bit_28_47 R_bl
Rbb_28_46 bitb_28_46 bitb_28_47 R_bl
Cb_28_46 bit_28_46 gnd C_bl
Cbb_28_46 bitb_28_46 gnd C_bl
Rb_28_47 bit_28_47 bit_28_48 R_bl
Rbb_28_47 bitb_28_47 bitb_28_48 R_bl
Cb_28_47 bit_28_47 gnd C_bl
Cbb_28_47 bitb_28_47 gnd C_bl
Rb_28_48 bit_28_48 bit_28_49 R_bl
Rbb_28_48 bitb_28_48 bitb_28_49 R_bl
Cb_28_48 bit_28_48 gnd C_bl
Cbb_28_48 bitb_28_48 gnd C_bl
Rb_28_49 bit_28_49 bit_28_50 R_bl
Rbb_28_49 bitb_28_49 bitb_28_50 R_bl
Cb_28_49 bit_28_49 gnd C_bl
Cbb_28_49 bitb_28_49 gnd C_bl
Rb_28_50 bit_28_50 bit_28_51 R_bl
Rbb_28_50 bitb_28_50 bitb_28_51 R_bl
Cb_28_50 bit_28_50 gnd C_bl
Cbb_28_50 bitb_28_50 gnd C_bl
Rb_28_51 bit_28_51 bit_28_52 R_bl
Rbb_28_51 bitb_28_51 bitb_28_52 R_bl
Cb_28_51 bit_28_51 gnd C_bl
Cbb_28_51 bitb_28_51 gnd C_bl
Rb_28_52 bit_28_52 bit_28_53 R_bl
Rbb_28_52 bitb_28_52 bitb_28_53 R_bl
Cb_28_52 bit_28_52 gnd C_bl
Cbb_28_52 bitb_28_52 gnd C_bl
Rb_28_53 bit_28_53 bit_28_54 R_bl
Rbb_28_53 bitb_28_53 bitb_28_54 R_bl
Cb_28_53 bit_28_53 gnd C_bl
Cbb_28_53 bitb_28_53 gnd C_bl
Rb_28_54 bit_28_54 bit_28_55 R_bl
Rbb_28_54 bitb_28_54 bitb_28_55 R_bl
Cb_28_54 bit_28_54 gnd C_bl
Cbb_28_54 bitb_28_54 gnd C_bl
Rb_28_55 bit_28_55 bit_28_56 R_bl
Rbb_28_55 bitb_28_55 bitb_28_56 R_bl
Cb_28_55 bit_28_55 gnd C_bl
Cbb_28_55 bitb_28_55 gnd C_bl
Rb_28_56 bit_28_56 bit_28_57 R_bl
Rbb_28_56 bitb_28_56 bitb_28_57 R_bl
Cb_28_56 bit_28_56 gnd C_bl
Cbb_28_56 bitb_28_56 gnd C_bl
Rb_28_57 bit_28_57 bit_28_58 R_bl
Rbb_28_57 bitb_28_57 bitb_28_58 R_bl
Cb_28_57 bit_28_57 gnd C_bl
Cbb_28_57 bitb_28_57 gnd C_bl
Rb_28_58 bit_28_58 bit_28_59 R_bl
Rbb_28_58 bitb_28_58 bitb_28_59 R_bl
Cb_28_58 bit_28_58 gnd C_bl
Cbb_28_58 bitb_28_58 gnd C_bl
Rb_28_59 bit_28_59 bit_28_60 R_bl
Rbb_28_59 bitb_28_59 bitb_28_60 R_bl
Cb_28_59 bit_28_59 gnd C_bl
Cbb_28_59 bitb_28_59 gnd C_bl
Rb_28_60 bit_28_60 bit_28_61 R_bl
Rbb_28_60 bitb_28_60 bitb_28_61 R_bl
Cb_28_60 bit_28_60 gnd C_bl
Cbb_28_60 bitb_28_60 gnd C_bl
Rb_28_61 bit_28_61 bit_28_62 R_bl
Rbb_28_61 bitb_28_61 bitb_28_62 R_bl
Cb_28_61 bit_28_61 gnd C_bl
Cbb_28_61 bitb_28_61 gnd C_bl
Rb_28_62 bit_28_62 bit_28_63 R_bl
Rbb_28_62 bitb_28_62 bitb_28_63 R_bl
Cb_28_62 bit_28_62 gnd C_bl
Cbb_28_62 bitb_28_62 gnd C_bl
Rb_28_63 bit_28_63 bit_28_64 R_bl
Rbb_28_63 bitb_28_63 bitb_28_64 R_bl
Cb_28_63 bit_28_63 gnd C_bl
Cbb_28_63 bitb_28_63 gnd C_bl
Rb_28_64 bit_28_64 bit_28_65 R_bl
Rbb_28_64 bitb_28_64 bitb_28_65 R_bl
Cb_28_64 bit_28_64 gnd C_bl
Cbb_28_64 bitb_28_64 gnd C_bl
Rb_28_65 bit_28_65 bit_28_66 R_bl
Rbb_28_65 bitb_28_65 bitb_28_66 R_bl
Cb_28_65 bit_28_65 gnd C_bl
Cbb_28_65 bitb_28_65 gnd C_bl
Rb_28_66 bit_28_66 bit_28_67 R_bl
Rbb_28_66 bitb_28_66 bitb_28_67 R_bl
Cb_28_66 bit_28_66 gnd C_bl
Cbb_28_66 bitb_28_66 gnd C_bl
Rb_28_67 bit_28_67 bit_28_68 R_bl
Rbb_28_67 bitb_28_67 bitb_28_68 R_bl
Cb_28_67 bit_28_67 gnd C_bl
Cbb_28_67 bitb_28_67 gnd C_bl
Rb_28_68 bit_28_68 bit_28_69 R_bl
Rbb_28_68 bitb_28_68 bitb_28_69 R_bl
Cb_28_68 bit_28_68 gnd C_bl
Cbb_28_68 bitb_28_68 gnd C_bl
Rb_28_69 bit_28_69 bit_28_70 R_bl
Rbb_28_69 bitb_28_69 bitb_28_70 R_bl
Cb_28_69 bit_28_69 gnd C_bl
Cbb_28_69 bitb_28_69 gnd C_bl
Rb_28_70 bit_28_70 bit_28_71 R_bl
Rbb_28_70 bitb_28_70 bitb_28_71 R_bl
Cb_28_70 bit_28_70 gnd C_bl
Cbb_28_70 bitb_28_70 gnd C_bl
Rb_28_71 bit_28_71 bit_28_72 R_bl
Rbb_28_71 bitb_28_71 bitb_28_72 R_bl
Cb_28_71 bit_28_71 gnd C_bl
Cbb_28_71 bitb_28_71 gnd C_bl
Rb_28_72 bit_28_72 bit_28_73 R_bl
Rbb_28_72 bitb_28_72 bitb_28_73 R_bl
Cb_28_72 bit_28_72 gnd C_bl
Cbb_28_72 bitb_28_72 gnd C_bl
Rb_28_73 bit_28_73 bit_28_74 R_bl
Rbb_28_73 bitb_28_73 bitb_28_74 R_bl
Cb_28_73 bit_28_73 gnd C_bl
Cbb_28_73 bitb_28_73 gnd C_bl
Rb_28_74 bit_28_74 bit_28_75 R_bl
Rbb_28_74 bitb_28_74 bitb_28_75 R_bl
Cb_28_74 bit_28_74 gnd C_bl
Cbb_28_74 bitb_28_74 gnd C_bl
Rb_28_75 bit_28_75 bit_28_76 R_bl
Rbb_28_75 bitb_28_75 bitb_28_76 R_bl
Cb_28_75 bit_28_75 gnd C_bl
Cbb_28_75 bitb_28_75 gnd C_bl
Rb_28_76 bit_28_76 bit_28_77 R_bl
Rbb_28_76 bitb_28_76 bitb_28_77 R_bl
Cb_28_76 bit_28_76 gnd C_bl
Cbb_28_76 bitb_28_76 gnd C_bl
Rb_28_77 bit_28_77 bit_28_78 R_bl
Rbb_28_77 bitb_28_77 bitb_28_78 R_bl
Cb_28_77 bit_28_77 gnd C_bl
Cbb_28_77 bitb_28_77 gnd C_bl
Rb_28_78 bit_28_78 bit_28_79 R_bl
Rbb_28_78 bitb_28_78 bitb_28_79 R_bl
Cb_28_78 bit_28_78 gnd C_bl
Cbb_28_78 bitb_28_78 gnd C_bl
Rb_28_79 bit_28_79 bit_28_80 R_bl
Rbb_28_79 bitb_28_79 bitb_28_80 R_bl
Cb_28_79 bit_28_79 gnd C_bl
Cbb_28_79 bitb_28_79 gnd C_bl
Rb_28_80 bit_28_80 bit_28_81 R_bl
Rbb_28_80 bitb_28_80 bitb_28_81 R_bl
Cb_28_80 bit_28_80 gnd C_bl
Cbb_28_80 bitb_28_80 gnd C_bl
Rb_28_81 bit_28_81 bit_28_82 R_bl
Rbb_28_81 bitb_28_81 bitb_28_82 R_bl
Cb_28_81 bit_28_81 gnd C_bl
Cbb_28_81 bitb_28_81 gnd C_bl
Rb_28_82 bit_28_82 bit_28_83 R_bl
Rbb_28_82 bitb_28_82 bitb_28_83 R_bl
Cb_28_82 bit_28_82 gnd C_bl
Cbb_28_82 bitb_28_82 gnd C_bl
Rb_28_83 bit_28_83 bit_28_84 R_bl
Rbb_28_83 bitb_28_83 bitb_28_84 R_bl
Cb_28_83 bit_28_83 gnd C_bl
Cbb_28_83 bitb_28_83 gnd C_bl
Rb_28_84 bit_28_84 bit_28_85 R_bl
Rbb_28_84 bitb_28_84 bitb_28_85 R_bl
Cb_28_84 bit_28_84 gnd C_bl
Cbb_28_84 bitb_28_84 gnd C_bl
Rb_28_85 bit_28_85 bit_28_86 R_bl
Rbb_28_85 bitb_28_85 bitb_28_86 R_bl
Cb_28_85 bit_28_85 gnd C_bl
Cbb_28_85 bitb_28_85 gnd C_bl
Rb_28_86 bit_28_86 bit_28_87 R_bl
Rbb_28_86 bitb_28_86 bitb_28_87 R_bl
Cb_28_86 bit_28_86 gnd C_bl
Cbb_28_86 bitb_28_86 gnd C_bl
Rb_28_87 bit_28_87 bit_28_88 R_bl
Rbb_28_87 bitb_28_87 bitb_28_88 R_bl
Cb_28_87 bit_28_87 gnd C_bl
Cbb_28_87 bitb_28_87 gnd C_bl
Rb_28_88 bit_28_88 bit_28_89 R_bl
Rbb_28_88 bitb_28_88 bitb_28_89 R_bl
Cb_28_88 bit_28_88 gnd C_bl
Cbb_28_88 bitb_28_88 gnd C_bl
Rb_28_89 bit_28_89 bit_28_90 R_bl
Rbb_28_89 bitb_28_89 bitb_28_90 R_bl
Cb_28_89 bit_28_89 gnd C_bl
Cbb_28_89 bitb_28_89 gnd C_bl
Rb_28_90 bit_28_90 bit_28_91 R_bl
Rbb_28_90 bitb_28_90 bitb_28_91 R_bl
Cb_28_90 bit_28_90 gnd C_bl
Cbb_28_90 bitb_28_90 gnd C_bl
Rb_28_91 bit_28_91 bit_28_92 R_bl
Rbb_28_91 bitb_28_91 bitb_28_92 R_bl
Cb_28_91 bit_28_91 gnd C_bl
Cbb_28_91 bitb_28_91 gnd C_bl
Rb_28_92 bit_28_92 bit_28_93 R_bl
Rbb_28_92 bitb_28_92 bitb_28_93 R_bl
Cb_28_92 bit_28_92 gnd C_bl
Cbb_28_92 bitb_28_92 gnd C_bl
Rb_28_93 bit_28_93 bit_28_94 R_bl
Rbb_28_93 bitb_28_93 bitb_28_94 R_bl
Cb_28_93 bit_28_93 gnd C_bl
Cbb_28_93 bitb_28_93 gnd C_bl
Rb_28_94 bit_28_94 bit_28_95 R_bl
Rbb_28_94 bitb_28_94 bitb_28_95 R_bl
Cb_28_94 bit_28_94 gnd C_bl
Cbb_28_94 bitb_28_94 gnd C_bl
Rb_28_95 bit_28_95 bit_28_96 R_bl
Rbb_28_95 bitb_28_95 bitb_28_96 R_bl
Cb_28_95 bit_28_95 gnd C_bl
Cbb_28_95 bitb_28_95 gnd C_bl
Rb_28_96 bit_28_96 bit_28_97 R_bl
Rbb_28_96 bitb_28_96 bitb_28_97 R_bl
Cb_28_96 bit_28_96 gnd C_bl
Cbb_28_96 bitb_28_96 gnd C_bl
Rb_28_97 bit_28_97 bit_28_98 R_bl
Rbb_28_97 bitb_28_97 bitb_28_98 R_bl
Cb_28_97 bit_28_97 gnd C_bl
Cbb_28_97 bitb_28_97 gnd C_bl
Rb_28_98 bit_28_98 bit_28_99 R_bl
Rbb_28_98 bitb_28_98 bitb_28_99 R_bl
Cb_28_98 bit_28_98 gnd C_bl
Cbb_28_98 bitb_28_98 gnd C_bl
Rb_28_99 bit_28_99 bit_28_100 R_bl
Rbb_28_99 bitb_28_99 bitb_28_100 R_bl
Cb_28_99 bit_28_99 gnd C_bl
Cbb_28_99 bitb_28_99 gnd C_bl
Rb_29_0 bit_29_0 bit_29_1 R_bl
Rbb_29_0 bitb_29_0 bitb_29_1 R_bl
Cb_29_0 bit_29_0 gnd C_bl
Cbb_29_0 bitb_29_0 gnd C_bl
Rb_29_1 bit_29_1 bit_29_2 R_bl
Rbb_29_1 bitb_29_1 bitb_29_2 R_bl
Cb_29_1 bit_29_1 gnd C_bl
Cbb_29_1 bitb_29_1 gnd C_bl
Rb_29_2 bit_29_2 bit_29_3 R_bl
Rbb_29_2 bitb_29_2 bitb_29_3 R_bl
Cb_29_2 bit_29_2 gnd C_bl
Cbb_29_2 bitb_29_2 gnd C_bl
Rb_29_3 bit_29_3 bit_29_4 R_bl
Rbb_29_3 bitb_29_3 bitb_29_4 R_bl
Cb_29_3 bit_29_3 gnd C_bl
Cbb_29_3 bitb_29_3 gnd C_bl
Rb_29_4 bit_29_4 bit_29_5 R_bl
Rbb_29_4 bitb_29_4 bitb_29_5 R_bl
Cb_29_4 bit_29_4 gnd C_bl
Cbb_29_4 bitb_29_4 gnd C_bl
Rb_29_5 bit_29_5 bit_29_6 R_bl
Rbb_29_5 bitb_29_5 bitb_29_6 R_bl
Cb_29_5 bit_29_5 gnd C_bl
Cbb_29_5 bitb_29_5 gnd C_bl
Rb_29_6 bit_29_6 bit_29_7 R_bl
Rbb_29_6 bitb_29_6 bitb_29_7 R_bl
Cb_29_6 bit_29_6 gnd C_bl
Cbb_29_6 bitb_29_6 gnd C_bl
Rb_29_7 bit_29_7 bit_29_8 R_bl
Rbb_29_7 bitb_29_7 bitb_29_8 R_bl
Cb_29_7 bit_29_7 gnd C_bl
Cbb_29_7 bitb_29_7 gnd C_bl
Rb_29_8 bit_29_8 bit_29_9 R_bl
Rbb_29_8 bitb_29_8 bitb_29_9 R_bl
Cb_29_8 bit_29_8 gnd C_bl
Cbb_29_8 bitb_29_8 gnd C_bl
Rb_29_9 bit_29_9 bit_29_10 R_bl
Rbb_29_9 bitb_29_9 bitb_29_10 R_bl
Cb_29_9 bit_29_9 gnd C_bl
Cbb_29_9 bitb_29_9 gnd C_bl
Rb_29_10 bit_29_10 bit_29_11 R_bl
Rbb_29_10 bitb_29_10 bitb_29_11 R_bl
Cb_29_10 bit_29_10 gnd C_bl
Cbb_29_10 bitb_29_10 gnd C_bl
Rb_29_11 bit_29_11 bit_29_12 R_bl
Rbb_29_11 bitb_29_11 bitb_29_12 R_bl
Cb_29_11 bit_29_11 gnd C_bl
Cbb_29_11 bitb_29_11 gnd C_bl
Rb_29_12 bit_29_12 bit_29_13 R_bl
Rbb_29_12 bitb_29_12 bitb_29_13 R_bl
Cb_29_12 bit_29_12 gnd C_bl
Cbb_29_12 bitb_29_12 gnd C_bl
Rb_29_13 bit_29_13 bit_29_14 R_bl
Rbb_29_13 bitb_29_13 bitb_29_14 R_bl
Cb_29_13 bit_29_13 gnd C_bl
Cbb_29_13 bitb_29_13 gnd C_bl
Rb_29_14 bit_29_14 bit_29_15 R_bl
Rbb_29_14 bitb_29_14 bitb_29_15 R_bl
Cb_29_14 bit_29_14 gnd C_bl
Cbb_29_14 bitb_29_14 gnd C_bl
Rb_29_15 bit_29_15 bit_29_16 R_bl
Rbb_29_15 bitb_29_15 bitb_29_16 R_bl
Cb_29_15 bit_29_15 gnd C_bl
Cbb_29_15 bitb_29_15 gnd C_bl
Rb_29_16 bit_29_16 bit_29_17 R_bl
Rbb_29_16 bitb_29_16 bitb_29_17 R_bl
Cb_29_16 bit_29_16 gnd C_bl
Cbb_29_16 bitb_29_16 gnd C_bl
Rb_29_17 bit_29_17 bit_29_18 R_bl
Rbb_29_17 bitb_29_17 bitb_29_18 R_bl
Cb_29_17 bit_29_17 gnd C_bl
Cbb_29_17 bitb_29_17 gnd C_bl
Rb_29_18 bit_29_18 bit_29_19 R_bl
Rbb_29_18 bitb_29_18 bitb_29_19 R_bl
Cb_29_18 bit_29_18 gnd C_bl
Cbb_29_18 bitb_29_18 gnd C_bl
Rb_29_19 bit_29_19 bit_29_20 R_bl
Rbb_29_19 bitb_29_19 bitb_29_20 R_bl
Cb_29_19 bit_29_19 gnd C_bl
Cbb_29_19 bitb_29_19 gnd C_bl
Rb_29_20 bit_29_20 bit_29_21 R_bl
Rbb_29_20 bitb_29_20 bitb_29_21 R_bl
Cb_29_20 bit_29_20 gnd C_bl
Cbb_29_20 bitb_29_20 gnd C_bl
Rb_29_21 bit_29_21 bit_29_22 R_bl
Rbb_29_21 bitb_29_21 bitb_29_22 R_bl
Cb_29_21 bit_29_21 gnd C_bl
Cbb_29_21 bitb_29_21 gnd C_bl
Rb_29_22 bit_29_22 bit_29_23 R_bl
Rbb_29_22 bitb_29_22 bitb_29_23 R_bl
Cb_29_22 bit_29_22 gnd C_bl
Cbb_29_22 bitb_29_22 gnd C_bl
Rb_29_23 bit_29_23 bit_29_24 R_bl
Rbb_29_23 bitb_29_23 bitb_29_24 R_bl
Cb_29_23 bit_29_23 gnd C_bl
Cbb_29_23 bitb_29_23 gnd C_bl
Rb_29_24 bit_29_24 bit_29_25 R_bl
Rbb_29_24 bitb_29_24 bitb_29_25 R_bl
Cb_29_24 bit_29_24 gnd C_bl
Cbb_29_24 bitb_29_24 gnd C_bl
Rb_29_25 bit_29_25 bit_29_26 R_bl
Rbb_29_25 bitb_29_25 bitb_29_26 R_bl
Cb_29_25 bit_29_25 gnd C_bl
Cbb_29_25 bitb_29_25 gnd C_bl
Rb_29_26 bit_29_26 bit_29_27 R_bl
Rbb_29_26 bitb_29_26 bitb_29_27 R_bl
Cb_29_26 bit_29_26 gnd C_bl
Cbb_29_26 bitb_29_26 gnd C_bl
Rb_29_27 bit_29_27 bit_29_28 R_bl
Rbb_29_27 bitb_29_27 bitb_29_28 R_bl
Cb_29_27 bit_29_27 gnd C_bl
Cbb_29_27 bitb_29_27 gnd C_bl
Rb_29_28 bit_29_28 bit_29_29 R_bl
Rbb_29_28 bitb_29_28 bitb_29_29 R_bl
Cb_29_28 bit_29_28 gnd C_bl
Cbb_29_28 bitb_29_28 gnd C_bl
Rb_29_29 bit_29_29 bit_29_30 R_bl
Rbb_29_29 bitb_29_29 bitb_29_30 R_bl
Cb_29_29 bit_29_29 gnd C_bl
Cbb_29_29 bitb_29_29 gnd C_bl
Rb_29_30 bit_29_30 bit_29_31 R_bl
Rbb_29_30 bitb_29_30 bitb_29_31 R_bl
Cb_29_30 bit_29_30 gnd C_bl
Cbb_29_30 bitb_29_30 gnd C_bl
Rb_29_31 bit_29_31 bit_29_32 R_bl
Rbb_29_31 bitb_29_31 bitb_29_32 R_bl
Cb_29_31 bit_29_31 gnd C_bl
Cbb_29_31 bitb_29_31 gnd C_bl
Rb_29_32 bit_29_32 bit_29_33 R_bl
Rbb_29_32 bitb_29_32 bitb_29_33 R_bl
Cb_29_32 bit_29_32 gnd C_bl
Cbb_29_32 bitb_29_32 gnd C_bl
Rb_29_33 bit_29_33 bit_29_34 R_bl
Rbb_29_33 bitb_29_33 bitb_29_34 R_bl
Cb_29_33 bit_29_33 gnd C_bl
Cbb_29_33 bitb_29_33 gnd C_bl
Rb_29_34 bit_29_34 bit_29_35 R_bl
Rbb_29_34 bitb_29_34 bitb_29_35 R_bl
Cb_29_34 bit_29_34 gnd C_bl
Cbb_29_34 bitb_29_34 gnd C_bl
Rb_29_35 bit_29_35 bit_29_36 R_bl
Rbb_29_35 bitb_29_35 bitb_29_36 R_bl
Cb_29_35 bit_29_35 gnd C_bl
Cbb_29_35 bitb_29_35 gnd C_bl
Rb_29_36 bit_29_36 bit_29_37 R_bl
Rbb_29_36 bitb_29_36 bitb_29_37 R_bl
Cb_29_36 bit_29_36 gnd C_bl
Cbb_29_36 bitb_29_36 gnd C_bl
Rb_29_37 bit_29_37 bit_29_38 R_bl
Rbb_29_37 bitb_29_37 bitb_29_38 R_bl
Cb_29_37 bit_29_37 gnd C_bl
Cbb_29_37 bitb_29_37 gnd C_bl
Rb_29_38 bit_29_38 bit_29_39 R_bl
Rbb_29_38 bitb_29_38 bitb_29_39 R_bl
Cb_29_38 bit_29_38 gnd C_bl
Cbb_29_38 bitb_29_38 gnd C_bl
Rb_29_39 bit_29_39 bit_29_40 R_bl
Rbb_29_39 bitb_29_39 bitb_29_40 R_bl
Cb_29_39 bit_29_39 gnd C_bl
Cbb_29_39 bitb_29_39 gnd C_bl
Rb_29_40 bit_29_40 bit_29_41 R_bl
Rbb_29_40 bitb_29_40 bitb_29_41 R_bl
Cb_29_40 bit_29_40 gnd C_bl
Cbb_29_40 bitb_29_40 gnd C_bl
Rb_29_41 bit_29_41 bit_29_42 R_bl
Rbb_29_41 bitb_29_41 bitb_29_42 R_bl
Cb_29_41 bit_29_41 gnd C_bl
Cbb_29_41 bitb_29_41 gnd C_bl
Rb_29_42 bit_29_42 bit_29_43 R_bl
Rbb_29_42 bitb_29_42 bitb_29_43 R_bl
Cb_29_42 bit_29_42 gnd C_bl
Cbb_29_42 bitb_29_42 gnd C_bl
Rb_29_43 bit_29_43 bit_29_44 R_bl
Rbb_29_43 bitb_29_43 bitb_29_44 R_bl
Cb_29_43 bit_29_43 gnd C_bl
Cbb_29_43 bitb_29_43 gnd C_bl
Rb_29_44 bit_29_44 bit_29_45 R_bl
Rbb_29_44 bitb_29_44 bitb_29_45 R_bl
Cb_29_44 bit_29_44 gnd C_bl
Cbb_29_44 bitb_29_44 gnd C_bl
Rb_29_45 bit_29_45 bit_29_46 R_bl
Rbb_29_45 bitb_29_45 bitb_29_46 R_bl
Cb_29_45 bit_29_45 gnd C_bl
Cbb_29_45 bitb_29_45 gnd C_bl
Rb_29_46 bit_29_46 bit_29_47 R_bl
Rbb_29_46 bitb_29_46 bitb_29_47 R_bl
Cb_29_46 bit_29_46 gnd C_bl
Cbb_29_46 bitb_29_46 gnd C_bl
Rb_29_47 bit_29_47 bit_29_48 R_bl
Rbb_29_47 bitb_29_47 bitb_29_48 R_bl
Cb_29_47 bit_29_47 gnd C_bl
Cbb_29_47 bitb_29_47 gnd C_bl
Rb_29_48 bit_29_48 bit_29_49 R_bl
Rbb_29_48 bitb_29_48 bitb_29_49 R_bl
Cb_29_48 bit_29_48 gnd C_bl
Cbb_29_48 bitb_29_48 gnd C_bl
Rb_29_49 bit_29_49 bit_29_50 R_bl
Rbb_29_49 bitb_29_49 bitb_29_50 R_bl
Cb_29_49 bit_29_49 gnd C_bl
Cbb_29_49 bitb_29_49 gnd C_bl
Rb_29_50 bit_29_50 bit_29_51 R_bl
Rbb_29_50 bitb_29_50 bitb_29_51 R_bl
Cb_29_50 bit_29_50 gnd C_bl
Cbb_29_50 bitb_29_50 gnd C_bl
Rb_29_51 bit_29_51 bit_29_52 R_bl
Rbb_29_51 bitb_29_51 bitb_29_52 R_bl
Cb_29_51 bit_29_51 gnd C_bl
Cbb_29_51 bitb_29_51 gnd C_bl
Rb_29_52 bit_29_52 bit_29_53 R_bl
Rbb_29_52 bitb_29_52 bitb_29_53 R_bl
Cb_29_52 bit_29_52 gnd C_bl
Cbb_29_52 bitb_29_52 gnd C_bl
Rb_29_53 bit_29_53 bit_29_54 R_bl
Rbb_29_53 bitb_29_53 bitb_29_54 R_bl
Cb_29_53 bit_29_53 gnd C_bl
Cbb_29_53 bitb_29_53 gnd C_bl
Rb_29_54 bit_29_54 bit_29_55 R_bl
Rbb_29_54 bitb_29_54 bitb_29_55 R_bl
Cb_29_54 bit_29_54 gnd C_bl
Cbb_29_54 bitb_29_54 gnd C_bl
Rb_29_55 bit_29_55 bit_29_56 R_bl
Rbb_29_55 bitb_29_55 bitb_29_56 R_bl
Cb_29_55 bit_29_55 gnd C_bl
Cbb_29_55 bitb_29_55 gnd C_bl
Rb_29_56 bit_29_56 bit_29_57 R_bl
Rbb_29_56 bitb_29_56 bitb_29_57 R_bl
Cb_29_56 bit_29_56 gnd C_bl
Cbb_29_56 bitb_29_56 gnd C_bl
Rb_29_57 bit_29_57 bit_29_58 R_bl
Rbb_29_57 bitb_29_57 bitb_29_58 R_bl
Cb_29_57 bit_29_57 gnd C_bl
Cbb_29_57 bitb_29_57 gnd C_bl
Rb_29_58 bit_29_58 bit_29_59 R_bl
Rbb_29_58 bitb_29_58 bitb_29_59 R_bl
Cb_29_58 bit_29_58 gnd C_bl
Cbb_29_58 bitb_29_58 gnd C_bl
Rb_29_59 bit_29_59 bit_29_60 R_bl
Rbb_29_59 bitb_29_59 bitb_29_60 R_bl
Cb_29_59 bit_29_59 gnd C_bl
Cbb_29_59 bitb_29_59 gnd C_bl
Rb_29_60 bit_29_60 bit_29_61 R_bl
Rbb_29_60 bitb_29_60 bitb_29_61 R_bl
Cb_29_60 bit_29_60 gnd C_bl
Cbb_29_60 bitb_29_60 gnd C_bl
Rb_29_61 bit_29_61 bit_29_62 R_bl
Rbb_29_61 bitb_29_61 bitb_29_62 R_bl
Cb_29_61 bit_29_61 gnd C_bl
Cbb_29_61 bitb_29_61 gnd C_bl
Rb_29_62 bit_29_62 bit_29_63 R_bl
Rbb_29_62 bitb_29_62 bitb_29_63 R_bl
Cb_29_62 bit_29_62 gnd C_bl
Cbb_29_62 bitb_29_62 gnd C_bl
Rb_29_63 bit_29_63 bit_29_64 R_bl
Rbb_29_63 bitb_29_63 bitb_29_64 R_bl
Cb_29_63 bit_29_63 gnd C_bl
Cbb_29_63 bitb_29_63 gnd C_bl
Rb_29_64 bit_29_64 bit_29_65 R_bl
Rbb_29_64 bitb_29_64 bitb_29_65 R_bl
Cb_29_64 bit_29_64 gnd C_bl
Cbb_29_64 bitb_29_64 gnd C_bl
Rb_29_65 bit_29_65 bit_29_66 R_bl
Rbb_29_65 bitb_29_65 bitb_29_66 R_bl
Cb_29_65 bit_29_65 gnd C_bl
Cbb_29_65 bitb_29_65 gnd C_bl
Rb_29_66 bit_29_66 bit_29_67 R_bl
Rbb_29_66 bitb_29_66 bitb_29_67 R_bl
Cb_29_66 bit_29_66 gnd C_bl
Cbb_29_66 bitb_29_66 gnd C_bl
Rb_29_67 bit_29_67 bit_29_68 R_bl
Rbb_29_67 bitb_29_67 bitb_29_68 R_bl
Cb_29_67 bit_29_67 gnd C_bl
Cbb_29_67 bitb_29_67 gnd C_bl
Rb_29_68 bit_29_68 bit_29_69 R_bl
Rbb_29_68 bitb_29_68 bitb_29_69 R_bl
Cb_29_68 bit_29_68 gnd C_bl
Cbb_29_68 bitb_29_68 gnd C_bl
Rb_29_69 bit_29_69 bit_29_70 R_bl
Rbb_29_69 bitb_29_69 bitb_29_70 R_bl
Cb_29_69 bit_29_69 gnd C_bl
Cbb_29_69 bitb_29_69 gnd C_bl
Rb_29_70 bit_29_70 bit_29_71 R_bl
Rbb_29_70 bitb_29_70 bitb_29_71 R_bl
Cb_29_70 bit_29_70 gnd C_bl
Cbb_29_70 bitb_29_70 gnd C_bl
Rb_29_71 bit_29_71 bit_29_72 R_bl
Rbb_29_71 bitb_29_71 bitb_29_72 R_bl
Cb_29_71 bit_29_71 gnd C_bl
Cbb_29_71 bitb_29_71 gnd C_bl
Rb_29_72 bit_29_72 bit_29_73 R_bl
Rbb_29_72 bitb_29_72 bitb_29_73 R_bl
Cb_29_72 bit_29_72 gnd C_bl
Cbb_29_72 bitb_29_72 gnd C_bl
Rb_29_73 bit_29_73 bit_29_74 R_bl
Rbb_29_73 bitb_29_73 bitb_29_74 R_bl
Cb_29_73 bit_29_73 gnd C_bl
Cbb_29_73 bitb_29_73 gnd C_bl
Rb_29_74 bit_29_74 bit_29_75 R_bl
Rbb_29_74 bitb_29_74 bitb_29_75 R_bl
Cb_29_74 bit_29_74 gnd C_bl
Cbb_29_74 bitb_29_74 gnd C_bl
Rb_29_75 bit_29_75 bit_29_76 R_bl
Rbb_29_75 bitb_29_75 bitb_29_76 R_bl
Cb_29_75 bit_29_75 gnd C_bl
Cbb_29_75 bitb_29_75 gnd C_bl
Rb_29_76 bit_29_76 bit_29_77 R_bl
Rbb_29_76 bitb_29_76 bitb_29_77 R_bl
Cb_29_76 bit_29_76 gnd C_bl
Cbb_29_76 bitb_29_76 gnd C_bl
Rb_29_77 bit_29_77 bit_29_78 R_bl
Rbb_29_77 bitb_29_77 bitb_29_78 R_bl
Cb_29_77 bit_29_77 gnd C_bl
Cbb_29_77 bitb_29_77 gnd C_bl
Rb_29_78 bit_29_78 bit_29_79 R_bl
Rbb_29_78 bitb_29_78 bitb_29_79 R_bl
Cb_29_78 bit_29_78 gnd C_bl
Cbb_29_78 bitb_29_78 gnd C_bl
Rb_29_79 bit_29_79 bit_29_80 R_bl
Rbb_29_79 bitb_29_79 bitb_29_80 R_bl
Cb_29_79 bit_29_79 gnd C_bl
Cbb_29_79 bitb_29_79 gnd C_bl
Rb_29_80 bit_29_80 bit_29_81 R_bl
Rbb_29_80 bitb_29_80 bitb_29_81 R_bl
Cb_29_80 bit_29_80 gnd C_bl
Cbb_29_80 bitb_29_80 gnd C_bl
Rb_29_81 bit_29_81 bit_29_82 R_bl
Rbb_29_81 bitb_29_81 bitb_29_82 R_bl
Cb_29_81 bit_29_81 gnd C_bl
Cbb_29_81 bitb_29_81 gnd C_bl
Rb_29_82 bit_29_82 bit_29_83 R_bl
Rbb_29_82 bitb_29_82 bitb_29_83 R_bl
Cb_29_82 bit_29_82 gnd C_bl
Cbb_29_82 bitb_29_82 gnd C_bl
Rb_29_83 bit_29_83 bit_29_84 R_bl
Rbb_29_83 bitb_29_83 bitb_29_84 R_bl
Cb_29_83 bit_29_83 gnd C_bl
Cbb_29_83 bitb_29_83 gnd C_bl
Rb_29_84 bit_29_84 bit_29_85 R_bl
Rbb_29_84 bitb_29_84 bitb_29_85 R_bl
Cb_29_84 bit_29_84 gnd C_bl
Cbb_29_84 bitb_29_84 gnd C_bl
Rb_29_85 bit_29_85 bit_29_86 R_bl
Rbb_29_85 bitb_29_85 bitb_29_86 R_bl
Cb_29_85 bit_29_85 gnd C_bl
Cbb_29_85 bitb_29_85 gnd C_bl
Rb_29_86 bit_29_86 bit_29_87 R_bl
Rbb_29_86 bitb_29_86 bitb_29_87 R_bl
Cb_29_86 bit_29_86 gnd C_bl
Cbb_29_86 bitb_29_86 gnd C_bl
Rb_29_87 bit_29_87 bit_29_88 R_bl
Rbb_29_87 bitb_29_87 bitb_29_88 R_bl
Cb_29_87 bit_29_87 gnd C_bl
Cbb_29_87 bitb_29_87 gnd C_bl
Rb_29_88 bit_29_88 bit_29_89 R_bl
Rbb_29_88 bitb_29_88 bitb_29_89 R_bl
Cb_29_88 bit_29_88 gnd C_bl
Cbb_29_88 bitb_29_88 gnd C_bl
Rb_29_89 bit_29_89 bit_29_90 R_bl
Rbb_29_89 bitb_29_89 bitb_29_90 R_bl
Cb_29_89 bit_29_89 gnd C_bl
Cbb_29_89 bitb_29_89 gnd C_bl
Rb_29_90 bit_29_90 bit_29_91 R_bl
Rbb_29_90 bitb_29_90 bitb_29_91 R_bl
Cb_29_90 bit_29_90 gnd C_bl
Cbb_29_90 bitb_29_90 gnd C_bl
Rb_29_91 bit_29_91 bit_29_92 R_bl
Rbb_29_91 bitb_29_91 bitb_29_92 R_bl
Cb_29_91 bit_29_91 gnd C_bl
Cbb_29_91 bitb_29_91 gnd C_bl
Rb_29_92 bit_29_92 bit_29_93 R_bl
Rbb_29_92 bitb_29_92 bitb_29_93 R_bl
Cb_29_92 bit_29_92 gnd C_bl
Cbb_29_92 bitb_29_92 gnd C_bl
Rb_29_93 bit_29_93 bit_29_94 R_bl
Rbb_29_93 bitb_29_93 bitb_29_94 R_bl
Cb_29_93 bit_29_93 gnd C_bl
Cbb_29_93 bitb_29_93 gnd C_bl
Rb_29_94 bit_29_94 bit_29_95 R_bl
Rbb_29_94 bitb_29_94 bitb_29_95 R_bl
Cb_29_94 bit_29_94 gnd C_bl
Cbb_29_94 bitb_29_94 gnd C_bl
Rb_29_95 bit_29_95 bit_29_96 R_bl
Rbb_29_95 bitb_29_95 bitb_29_96 R_bl
Cb_29_95 bit_29_95 gnd C_bl
Cbb_29_95 bitb_29_95 gnd C_bl
Rb_29_96 bit_29_96 bit_29_97 R_bl
Rbb_29_96 bitb_29_96 bitb_29_97 R_bl
Cb_29_96 bit_29_96 gnd C_bl
Cbb_29_96 bitb_29_96 gnd C_bl
Rb_29_97 bit_29_97 bit_29_98 R_bl
Rbb_29_97 bitb_29_97 bitb_29_98 R_bl
Cb_29_97 bit_29_97 gnd C_bl
Cbb_29_97 bitb_29_97 gnd C_bl
Rb_29_98 bit_29_98 bit_29_99 R_bl
Rbb_29_98 bitb_29_98 bitb_29_99 R_bl
Cb_29_98 bit_29_98 gnd C_bl
Cbb_29_98 bitb_29_98 gnd C_bl
Rb_29_99 bit_29_99 bit_29_100 R_bl
Rbb_29_99 bitb_29_99 bitb_29_100 R_bl
Cb_29_99 bit_29_99 gnd C_bl
Cbb_29_99 bitb_29_99 gnd C_bl
Rb_30_0 bit_30_0 bit_30_1 R_bl
Rbb_30_0 bitb_30_0 bitb_30_1 R_bl
Cb_30_0 bit_30_0 gnd C_bl
Cbb_30_0 bitb_30_0 gnd C_bl
Rb_30_1 bit_30_1 bit_30_2 R_bl
Rbb_30_1 bitb_30_1 bitb_30_2 R_bl
Cb_30_1 bit_30_1 gnd C_bl
Cbb_30_1 bitb_30_1 gnd C_bl
Rb_30_2 bit_30_2 bit_30_3 R_bl
Rbb_30_2 bitb_30_2 bitb_30_3 R_bl
Cb_30_2 bit_30_2 gnd C_bl
Cbb_30_2 bitb_30_2 gnd C_bl
Rb_30_3 bit_30_3 bit_30_4 R_bl
Rbb_30_3 bitb_30_3 bitb_30_4 R_bl
Cb_30_3 bit_30_3 gnd C_bl
Cbb_30_3 bitb_30_3 gnd C_bl
Rb_30_4 bit_30_4 bit_30_5 R_bl
Rbb_30_4 bitb_30_4 bitb_30_5 R_bl
Cb_30_4 bit_30_4 gnd C_bl
Cbb_30_4 bitb_30_4 gnd C_bl
Rb_30_5 bit_30_5 bit_30_6 R_bl
Rbb_30_5 bitb_30_5 bitb_30_6 R_bl
Cb_30_5 bit_30_5 gnd C_bl
Cbb_30_5 bitb_30_5 gnd C_bl
Rb_30_6 bit_30_6 bit_30_7 R_bl
Rbb_30_6 bitb_30_6 bitb_30_7 R_bl
Cb_30_6 bit_30_6 gnd C_bl
Cbb_30_6 bitb_30_6 gnd C_bl
Rb_30_7 bit_30_7 bit_30_8 R_bl
Rbb_30_7 bitb_30_7 bitb_30_8 R_bl
Cb_30_7 bit_30_7 gnd C_bl
Cbb_30_7 bitb_30_7 gnd C_bl
Rb_30_8 bit_30_8 bit_30_9 R_bl
Rbb_30_8 bitb_30_8 bitb_30_9 R_bl
Cb_30_8 bit_30_8 gnd C_bl
Cbb_30_8 bitb_30_8 gnd C_bl
Rb_30_9 bit_30_9 bit_30_10 R_bl
Rbb_30_9 bitb_30_9 bitb_30_10 R_bl
Cb_30_9 bit_30_9 gnd C_bl
Cbb_30_9 bitb_30_9 gnd C_bl
Rb_30_10 bit_30_10 bit_30_11 R_bl
Rbb_30_10 bitb_30_10 bitb_30_11 R_bl
Cb_30_10 bit_30_10 gnd C_bl
Cbb_30_10 bitb_30_10 gnd C_bl
Rb_30_11 bit_30_11 bit_30_12 R_bl
Rbb_30_11 bitb_30_11 bitb_30_12 R_bl
Cb_30_11 bit_30_11 gnd C_bl
Cbb_30_11 bitb_30_11 gnd C_bl
Rb_30_12 bit_30_12 bit_30_13 R_bl
Rbb_30_12 bitb_30_12 bitb_30_13 R_bl
Cb_30_12 bit_30_12 gnd C_bl
Cbb_30_12 bitb_30_12 gnd C_bl
Rb_30_13 bit_30_13 bit_30_14 R_bl
Rbb_30_13 bitb_30_13 bitb_30_14 R_bl
Cb_30_13 bit_30_13 gnd C_bl
Cbb_30_13 bitb_30_13 gnd C_bl
Rb_30_14 bit_30_14 bit_30_15 R_bl
Rbb_30_14 bitb_30_14 bitb_30_15 R_bl
Cb_30_14 bit_30_14 gnd C_bl
Cbb_30_14 bitb_30_14 gnd C_bl
Rb_30_15 bit_30_15 bit_30_16 R_bl
Rbb_30_15 bitb_30_15 bitb_30_16 R_bl
Cb_30_15 bit_30_15 gnd C_bl
Cbb_30_15 bitb_30_15 gnd C_bl
Rb_30_16 bit_30_16 bit_30_17 R_bl
Rbb_30_16 bitb_30_16 bitb_30_17 R_bl
Cb_30_16 bit_30_16 gnd C_bl
Cbb_30_16 bitb_30_16 gnd C_bl
Rb_30_17 bit_30_17 bit_30_18 R_bl
Rbb_30_17 bitb_30_17 bitb_30_18 R_bl
Cb_30_17 bit_30_17 gnd C_bl
Cbb_30_17 bitb_30_17 gnd C_bl
Rb_30_18 bit_30_18 bit_30_19 R_bl
Rbb_30_18 bitb_30_18 bitb_30_19 R_bl
Cb_30_18 bit_30_18 gnd C_bl
Cbb_30_18 bitb_30_18 gnd C_bl
Rb_30_19 bit_30_19 bit_30_20 R_bl
Rbb_30_19 bitb_30_19 bitb_30_20 R_bl
Cb_30_19 bit_30_19 gnd C_bl
Cbb_30_19 bitb_30_19 gnd C_bl
Rb_30_20 bit_30_20 bit_30_21 R_bl
Rbb_30_20 bitb_30_20 bitb_30_21 R_bl
Cb_30_20 bit_30_20 gnd C_bl
Cbb_30_20 bitb_30_20 gnd C_bl
Rb_30_21 bit_30_21 bit_30_22 R_bl
Rbb_30_21 bitb_30_21 bitb_30_22 R_bl
Cb_30_21 bit_30_21 gnd C_bl
Cbb_30_21 bitb_30_21 gnd C_bl
Rb_30_22 bit_30_22 bit_30_23 R_bl
Rbb_30_22 bitb_30_22 bitb_30_23 R_bl
Cb_30_22 bit_30_22 gnd C_bl
Cbb_30_22 bitb_30_22 gnd C_bl
Rb_30_23 bit_30_23 bit_30_24 R_bl
Rbb_30_23 bitb_30_23 bitb_30_24 R_bl
Cb_30_23 bit_30_23 gnd C_bl
Cbb_30_23 bitb_30_23 gnd C_bl
Rb_30_24 bit_30_24 bit_30_25 R_bl
Rbb_30_24 bitb_30_24 bitb_30_25 R_bl
Cb_30_24 bit_30_24 gnd C_bl
Cbb_30_24 bitb_30_24 gnd C_bl
Rb_30_25 bit_30_25 bit_30_26 R_bl
Rbb_30_25 bitb_30_25 bitb_30_26 R_bl
Cb_30_25 bit_30_25 gnd C_bl
Cbb_30_25 bitb_30_25 gnd C_bl
Rb_30_26 bit_30_26 bit_30_27 R_bl
Rbb_30_26 bitb_30_26 bitb_30_27 R_bl
Cb_30_26 bit_30_26 gnd C_bl
Cbb_30_26 bitb_30_26 gnd C_bl
Rb_30_27 bit_30_27 bit_30_28 R_bl
Rbb_30_27 bitb_30_27 bitb_30_28 R_bl
Cb_30_27 bit_30_27 gnd C_bl
Cbb_30_27 bitb_30_27 gnd C_bl
Rb_30_28 bit_30_28 bit_30_29 R_bl
Rbb_30_28 bitb_30_28 bitb_30_29 R_bl
Cb_30_28 bit_30_28 gnd C_bl
Cbb_30_28 bitb_30_28 gnd C_bl
Rb_30_29 bit_30_29 bit_30_30 R_bl
Rbb_30_29 bitb_30_29 bitb_30_30 R_bl
Cb_30_29 bit_30_29 gnd C_bl
Cbb_30_29 bitb_30_29 gnd C_bl
Rb_30_30 bit_30_30 bit_30_31 R_bl
Rbb_30_30 bitb_30_30 bitb_30_31 R_bl
Cb_30_30 bit_30_30 gnd C_bl
Cbb_30_30 bitb_30_30 gnd C_bl
Rb_30_31 bit_30_31 bit_30_32 R_bl
Rbb_30_31 bitb_30_31 bitb_30_32 R_bl
Cb_30_31 bit_30_31 gnd C_bl
Cbb_30_31 bitb_30_31 gnd C_bl
Rb_30_32 bit_30_32 bit_30_33 R_bl
Rbb_30_32 bitb_30_32 bitb_30_33 R_bl
Cb_30_32 bit_30_32 gnd C_bl
Cbb_30_32 bitb_30_32 gnd C_bl
Rb_30_33 bit_30_33 bit_30_34 R_bl
Rbb_30_33 bitb_30_33 bitb_30_34 R_bl
Cb_30_33 bit_30_33 gnd C_bl
Cbb_30_33 bitb_30_33 gnd C_bl
Rb_30_34 bit_30_34 bit_30_35 R_bl
Rbb_30_34 bitb_30_34 bitb_30_35 R_bl
Cb_30_34 bit_30_34 gnd C_bl
Cbb_30_34 bitb_30_34 gnd C_bl
Rb_30_35 bit_30_35 bit_30_36 R_bl
Rbb_30_35 bitb_30_35 bitb_30_36 R_bl
Cb_30_35 bit_30_35 gnd C_bl
Cbb_30_35 bitb_30_35 gnd C_bl
Rb_30_36 bit_30_36 bit_30_37 R_bl
Rbb_30_36 bitb_30_36 bitb_30_37 R_bl
Cb_30_36 bit_30_36 gnd C_bl
Cbb_30_36 bitb_30_36 gnd C_bl
Rb_30_37 bit_30_37 bit_30_38 R_bl
Rbb_30_37 bitb_30_37 bitb_30_38 R_bl
Cb_30_37 bit_30_37 gnd C_bl
Cbb_30_37 bitb_30_37 gnd C_bl
Rb_30_38 bit_30_38 bit_30_39 R_bl
Rbb_30_38 bitb_30_38 bitb_30_39 R_bl
Cb_30_38 bit_30_38 gnd C_bl
Cbb_30_38 bitb_30_38 gnd C_bl
Rb_30_39 bit_30_39 bit_30_40 R_bl
Rbb_30_39 bitb_30_39 bitb_30_40 R_bl
Cb_30_39 bit_30_39 gnd C_bl
Cbb_30_39 bitb_30_39 gnd C_bl
Rb_30_40 bit_30_40 bit_30_41 R_bl
Rbb_30_40 bitb_30_40 bitb_30_41 R_bl
Cb_30_40 bit_30_40 gnd C_bl
Cbb_30_40 bitb_30_40 gnd C_bl
Rb_30_41 bit_30_41 bit_30_42 R_bl
Rbb_30_41 bitb_30_41 bitb_30_42 R_bl
Cb_30_41 bit_30_41 gnd C_bl
Cbb_30_41 bitb_30_41 gnd C_bl
Rb_30_42 bit_30_42 bit_30_43 R_bl
Rbb_30_42 bitb_30_42 bitb_30_43 R_bl
Cb_30_42 bit_30_42 gnd C_bl
Cbb_30_42 bitb_30_42 gnd C_bl
Rb_30_43 bit_30_43 bit_30_44 R_bl
Rbb_30_43 bitb_30_43 bitb_30_44 R_bl
Cb_30_43 bit_30_43 gnd C_bl
Cbb_30_43 bitb_30_43 gnd C_bl
Rb_30_44 bit_30_44 bit_30_45 R_bl
Rbb_30_44 bitb_30_44 bitb_30_45 R_bl
Cb_30_44 bit_30_44 gnd C_bl
Cbb_30_44 bitb_30_44 gnd C_bl
Rb_30_45 bit_30_45 bit_30_46 R_bl
Rbb_30_45 bitb_30_45 bitb_30_46 R_bl
Cb_30_45 bit_30_45 gnd C_bl
Cbb_30_45 bitb_30_45 gnd C_bl
Rb_30_46 bit_30_46 bit_30_47 R_bl
Rbb_30_46 bitb_30_46 bitb_30_47 R_bl
Cb_30_46 bit_30_46 gnd C_bl
Cbb_30_46 bitb_30_46 gnd C_bl
Rb_30_47 bit_30_47 bit_30_48 R_bl
Rbb_30_47 bitb_30_47 bitb_30_48 R_bl
Cb_30_47 bit_30_47 gnd C_bl
Cbb_30_47 bitb_30_47 gnd C_bl
Rb_30_48 bit_30_48 bit_30_49 R_bl
Rbb_30_48 bitb_30_48 bitb_30_49 R_bl
Cb_30_48 bit_30_48 gnd C_bl
Cbb_30_48 bitb_30_48 gnd C_bl
Rb_30_49 bit_30_49 bit_30_50 R_bl
Rbb_30_49 bitb_30_49 bitb_30_50 R_bl
Cb_30_49 bit_30_49 gnd C_bl
Cbb_30_49 bitb_30_49 gnd C_bl
Rb_30_50 bit_30_50 bit_30_51 R_bl
Rbb_30_50 bitb_30_50 bitb_30_51 R_bl
Cb_30_50 bit_30_50 gnd C_bl
Cbb_30_50 bitb_30_50 gnd C_bl
Rb_30_51 bit_30_51 bit_30_52 R_bl
Rbb_30_51 bitb_30_51 bitb_30_52 R_bl
Cb_30_51 bit_30_51 gnd C_bl
Cbb_30_51 bitb_30_51 gnd C_bl
Rb_30_52 bit_30_52 bit_30_53 R_bl
Rbb_30_52 bitb_30_52 bitb_30_53 R_bl
Cb_30_52 bit_30_52 gnd C_bl
Cbb_30_52 bitb_30_52 gnd C_bl
Rb_30_53 bit_30_53 bit_30_54 R_bl
Rbb_30_53 bitb_30_53 bitb_30_54 R_bl
Cb_30_53 bit_30_53 gnd C_bl
Cbb_30_53 bitb_30_53 gnd C_bl
Rb_30_54 bit_30_54 bit_30_55 R_bl
Rbb_30_54 bitb_30_54 bitb_30_55 R_bl
Cb_30_54 bit_30_54 gnd C_bl
Cbb_30_54 bitb_30_54 gnd C_bl
Rb_30_55 bit_30_55 bit_30_56 R_bl
Rbb_30_55 bitb_30_55 bitb_30_56 R_bl
Cb_30_55 bit_30_55 gnd C_bl
Cbb_30_55 bitb_30_55 gnd C_bl
Rb_30_56 bit_30_56 bit_30_57 R_bl
Rbb_30_56 bitb_30_56 bitb_30_57 R_bl
Cb_30_56 bit_30_56 gnd C_bl
Cbb_30_56 bitb_30_56 gnd C_bl
Rb_30_57 bit_30_57 bit_30_58 R_bl
Rbb_30_57 bitb_30_57 bitb_30_58 R_bl
Cb_30_57 bit_30_57 gnd C_bl
Cbb_30_57 bitb_30_57 gnd C_bl
Rb_30_58 bit_30_58 bit_30_59 R_bl
Rbb_30_58 bitb_30_58 bitb_30_59 R_bl
Cb_30_58 bit_30_58 gnd C_bl
Cbb_30_58 bitb_30_58 gnd C_bl
Rb_30_59 bit_30_59 bit_30_60 R_bl
Rbb_30_59 bitb_30_59 bitb_30_60 R_bl
Cb_30_59 bit_30_59 gnd C_bl
Cbb_30_59 bitb_30_59 gnd C_bl
Rb_30_60 bit_30_60 bit_30_61 R_bl
Rbb_30_60 bitb_30_60 bitb_30_61 R_bl
Cb_30_60 bit_30_60 gnd C_bl
Cbb_30_60 bitb_30_60 gnd C_bl
Rb_30_61 bit_30_61 bit_30_62 R_bl
Rbb_30_61 bitb_30_61 bitb_30_62 R_bl
Cb_30_61 bit_30_61 gnd C_bl
Cbb_30_61 bitb_30_61 gnd C_bl
Rb_30_62 bit_30_62 bit_30_63 R_bl
Rbb_30_62 bitb_30_62 bitb_30_63 R_bl
Cb_30_62 bit_30_62 gnd C_bl
Cbb_30_62 bitb_30_62 gnd C_bl
Rb_30_63 bit_30_63 bit_30_64 R_bl
Rbb_30_63 bitb_30_63 bitb_30_64 R_bl
Cb_30_63 bit_30_63 gnd C_bl
Cbb_30_63 bitb_30_63 gnd C_bl
Rb_30_64 bit_30_64 bit_30_65 R_bl
Rbb_30_64 bitb_30_64 bitb_30_65 R_bl
Cb_30_64 bit_30_64 gnd C_bl
Cbb_30_64 bitb_30_64 gnd C_bl
Rb_30_65 bit_30_65 bit_30_66 R_bl
Rbb_30_65 bitb_30_65 bitb_30_66 R_bl
Cb_30_65 bit_30_65 gnd C_bl
Cbb_30_65 bitb_30_65 gnd C_bl
Rb_30_66 bit_30_66 bit_30_67 R_bl
Rbb_30_66 bitb_30_66 bitb_30_67 R_bl
Cb_30_66 bit_30_66 gnd C_bl
Cbb_30_66 bitb_30_66 gnd C_bl
Rb_30_67 bit_30_67 bit_30_68 R_bl
Rbb_30_67 bitb_30_67 bitb_30_68 R_bl
Cb_30_67 bit_30_67 gnd C_bl
Cbb_30_67 bitb_30_67 gnd C_bl
Rb_30_68 bit_30_68 bit_30_69 R_bl
Rbb_30_68 bitb_30_68 bitb_30_69 R_bl
Cb_30_68 bit_30_68 gnd C_bl
Cbb_30_68 bitb_30_68 gnd C_bl
Rb_30_69 bit_30_69 bit_30_70 R_bl
Rbb_30_69 bitb_30_69 bitb_30_70 R_bl
Cb_30_69 bit_30_69 gnd C_bl
Cbb_30_69 bitb_30_69 gnd C_bl
Rb_30_70 bit_30_70 bit_30_71 R_bl
Rbb_30_70 bitb_30_70 bitb_30_71 R_bl
Cb_30_70 bit_30_70 gnd C_bl
Cbb_30_70 bitb_30_70 gnd C_bl
Rb_30_71 bit_30_71 bit_30_72 R_bl
Rbb_30_71 bitb_30_71 bitb_30_72 R_bl
Cb_30_71 bit_30_71 gnd C_bl
Cbb_30_71 bitb_30_71 gnd C_bl
Rb_30_72 bit_30_72 bit_30_73 R_bl
Rbb_30_72 bitb_30_72 bitb_30_73 R_bl
Cb_30_72 bit_30_72 gnd C_bl
Cbb_30_72 bitb_30_72 gnd C_bl
Rb_30_73 bit_30_73 bit_30_74 R_bl
Rbb_30_73 bitb_30_73 bitb_30_74 R_bl
Cb_30_73 bit_30_73 gnd C_bl
Cbb_30_73 bitb_30_73 gnd C_bl
Rb_30_74 bit_30_74 bit_30_75 R_bl
Rbb_30_74 bitb_30_74 bitb_30_75 R_bl
Cb_30_74 bit_30_74 gnd C_bl
Cbb_30_74 bitb_30_74 gnd C_bl
Rb_30_75 bit_30_75 bit_30_76 R_bl
Rbb_30_75 bitb_30_75 bitb_30_76 R_bl
Cb_30_75 bit_30_75 gnd C_bl
Cbb_30_75 bitb_30_75 gnd C_bl
Rb_30_76 bit_30_76 bit_30_77 R_bl
Rbb_30_76 bitb_30_76 bitb_30_77 R_bl
Cb_30_76 bit_30_76 gnd C_bl
Cbb_30_76 bitb_30_76 gnd C_bl
Rb_30_77 bit_30_77 bit_30_78 R_bl
Rbb_30_77 bitb_30_77 bitb_30_78 R_bl
Cb_30_77 bit_30_77 gnd C_bl
Cbb_30_77 bitb_30_77 gnd C_bl
Rb_30_78 bit_30_78 bit_30_79 R_bl
Rbb_30_78 bitb_30_78 bitb_30_79 R_bl
Cb_30_78 bit_30_78 gnd C_bl
Cbb_30_78 bitb_30_78 gnd C_bl
Rb_30_79 bit_30_79 bit_30_80 R_bl
Rbb_30_79 bitb_30_79 bitb_30_80 R_bl
Cb_30_79 bit_30_79 gnd C_bl
Cbb_30_79 bitb_30_79 gnd C_bl
Rb_30_80 bit_30_80 bit_30_81 R_bl
Rbb_30_80 bitb_30_80 bitb_30_81 R_bl
Cb_30_80 bit_30_80 gnd C_bl
Cbb_30_80 bitb_30_80 gnd C_bl
Rb_30_81 bit_30_81 bit_30_82 R_bl
Rbb_30_81 bitb_30_81 bitb_30_82 R_bl
Cb_30_81 bit_30_81 gnd C_bl
Cbb_30_81 bitb_30_81 gnd C_bl
Rb_30_82 bit_30_82 bit_30_83 R_bl
Rbb_30_82 bitb_30_82 bitb_30_83 R_bl
Cb_30_82 bit_30_82 gnd C_bl
Cbb_30_82 bitb_30_82 gnd C_bl
Rb_30_83 bit_30_83 bit_30_84 R_bl
Rbb_30_83 bitb_30_83 bitb_30_84 R_bl
Cb_30_83 bit_30_83 gnd C_bl
Cbb_30_83 bitb_30_83 gnd C_bl
Rb_30_84 bit_30_84 bit_30_85 R_bl
Rbb_30_84 bitb_30_84 bitb_30_85 R_bl
Cb_30_84 bit_30_84 gnd C_bl
Cbb_30_84 bitb_30_84 gnd C_bl
Rb_30_85 bit_30_85 bit_30_86 R_bl
Rbb_30_85 bitb_30_85 bitb_30_86 R_bl
Cb_30_85 bit_30_85 gnd C_bl
Cbb_30_85 bitb_30_85 gnd C_bl
Rb_30_86 bit_30_86 bit_30_87 R_bl
Rbb_30_86 bitb_30_86 bitb_30_87 R_bl
Cb_30_86 bit_30_86 gnd C_bl
Cbb_30_86 bitb_30_86 gnd C_bl
Rb_30_87 bit_30_87 bit_30_88 R_bl
Rbb_30_87 bitb_30_87 bitb_30_88 R_bl
Cb_30_87 bit_30_87 gnd C_bl
Cbb_30_87 bitb_30_87 gnd C_bl
Rb_30_88 bit_30_88 bit_30_89 R_bl
Rbb_30_88 bitb_30_88 bitb_30_89 R_bl
Cb_30_88 bit_30_88 gnd C_bl
Cbb_30_88 bitb_30_88 gnd C_bl
Rb_30_89 bit_30_89 bit_30_90 R_bl
Rbb_30_89 bitb_30_89 bitb_30_90 R_bl
Cb_30_89 bit_30_89 gnd C_bl
Cbb_30_89 bitb_30_89 gnd C_bl
Rb_30_90 bit_30_90 bit_30_91 R_bl
Rbb_30_90 bitb_30_90 bitb_30_91 R_bl
Cb_30_90 bit_30_90 gnd C_bl
Cbb_30_90 bitb_30_90 gnd C_bl
Rb_30_91 bit_30_91 bit_30_92 R_bl
Rbb_30_91 bitb_30_91 bitb_30_92 R_bl
Cb_30_91 bit_30_91 gnd C_bl
Cbb_30_91 bitb_30_91 gnd C_bl
Rb_30_92 bit_30_92 bit_30_93 R_bl
Rbb_30_92 bitb_30_92 bitb_30_93 R_bl
Cb_30_92 bit_30_92 gnd C_bl
Cbb_30_92 bitb_30_92 gnd C_bl
Rb_30_93 bit_30_93 bit_30_94 R_bl
Rbb_30_93 bitb_30_93 bitb_30_94 R_bl
Cb_30_93 bit_30_93 gnd C_bl
Cbb_30_93 bitb_30_93 gnd C_bl
Rb_30_94 bit_30_94 bit_30_95 R_bl
Rbb_30_94 bitb_30_94 bitb_30_95 R_bl
Cb_30_94 bit_30_94 gnd C_bl
Cbb_30_94 bitb_30_94 gnd C_bl
Rb_30_95 bit_30_95 bit_30_96 R_bl
Rbb_30_95 bitb_30_95 bitb_30_96 R_bl
Cb_30_95 bit_30_95 gnd C_bl
Cbb_30_95 bitb_30_95 gnd C_bl
Rb_30_96 bit_30_96 bit_30_97 R_bl
Rbb_30_96 bitb_30_96 bitb_30_97 R_bl
Cb_30_96 bit_30_96 gnd C_bl
Cbb_30_96 bitb_30_96 gnd C_bl
Rb_30_97 bit_30_97 bit_30_98 R_bl
Rbb_30_97 bitb_30_97 bitb_30_98 R_bl
Cb_30_97 bit_30_97 gnd C_bl
Cbb_30_97 bitb_30_97 gnd C_bl
Rb_30_98 bit_30_98 bit_30_99 R_bl
Rbb_30_98 bitb_30_98 bitb_30_99 R_bl
Cb_30_98 bit_30_98 gnd C_bl
Cbb_30_98 bitb_30_98 gnd C_bl
Rb_30_99 bit_30_99 bit_30_100 R_bl
Rbb_30_99 bitb_30_99 bitb_30_100 R_bl
Cb_30_99 bit_30_99 gnd C_bl
Cbb_30_99 bitb_30_99 gnd C_bl
Rb_31_0 bit_31_0 bit_31_1 R_bl
Rbb_31_0 bitb_31_0 bitb_31_1 R_bl
Cb_31_0 bit_31_0 gnd C_bl
Cbb_31_0 bitb_31_0 gnd C_bl
Rb_31_1 bit_31_1 bit_31_2 R_bl
Rbb_31_1 bitb_31_1 bitb_31_2 R_bl
Cb_31_1 bit_31_1 gnd C_bl
Cbb_31_1 bitb_31_1 gnd C_bl
Rb_31_2 bit_31_2 bit_31_3 R_bl
Rbb_31_2 bitb_31_2 bitb_31_3 R_bl
Cb_31_2 bit_31_2 gnd C_bl
Cbb_31_2 bitb_31_2 gnd C_bl
Rb_31_3 bit_31_3 bit_31_4 R_bl
Rbb_31_3 bitb_31_3 bitb_31_4 R_bl
Cb_31_3 bit_31_3 gnd C_bl
Cbb_31_3 bitb_31_3 gnd C_bl
Rb_31_4 bit_31_4 bit_31_5 R_bl
Rbb_31_4 bitb_31_4 bitb_31_5 R_bl
Cb_31_4 bit_31_4 gnd C_bl
Cbb_31_4 bitb_31_4 gnd C_bl
Rb_31_5 bit_31_5 bit_31_6 R_bl
Rbb_31_5 bitb_31_5 bitb_31_6 R_bl
Cb_31_5 bit_31_5 gnd C_bl
Cbb_31_5 bitb_31_5 gnd C_bl
Rb_31_6 bit_31_6 bit_31_7 R_bl
Rbb_31_6 bitb_31_6 bitb_31_7 R_bl
Cb_31_6 bit_31_6 gnd C_bl
Cbb_31_6 bitb_31_6 gnd C_bl
Rb_31_7 bit_31_7 bit_31_8 R_bl
Rbb_31_7 bitb_31_7 bitb_31_8 R_bl
Cb_31_7 bit_31_7 gnd C_bl
Cbb_31_7 bitb_31_7 gnd C_bl
Rb_31_8 bit_31_8 bit_31_9 R_bl
Rbb_31_8 bitb_31_8 bitb_31_9 R_bl
Cb_31_8 bit_31_8 gnd C_bl
Cbb_31_8 bitb_31_8 gnd C_bl
Rb_31_9 bit_31_9 bit_31_10 R_bl
Rbb_31_9 bitb_31_9 bitb_31_10 R_bl
Cb_31_9 bit_31_9 gnd C_bl
Cbb_31_9 bitb_31_9 gnd C_bl
Rb_31_10 bit_31_10 bit_31_11 R_bl
Rbb_31_10 bitb_31_10 bitb_31_11 R_bl
Cb_31_10 bit_31_10 gnd C_bl
Cbb_31_10 bitb_31_10 gnd C_bl
Rb_31_11 bit_31_11 bit_31_12 R_bl
Rbb_31_11 bitb_31_11 bitb_31_12 R_bl
Cb_31_11 bit_31_11 gnd C_bl
Cbb_31_11 bitb_31_11 gnd C_bl
Rb_31_12 bit_31_12 bit_31_13 R_bl
Rbb_31_12 bitb_31_12 bitb_31_13 R_bl
Cb_31_12 bit_31_12 gnd C_bl
Cbb_31_12 bitb_31_12 gnd C_bl
Rb_31_13 bit_31_13 bit_31_14 R_bl
Rbb_31_13 bitb_31_13 bitb_31_14 R_bl
Cb_31_13 bit_31_13 gnd C_bl
Cbb_31_13 bitb_31_13 gnd C_bl
Rb_31_14 bit_31_14 bit_31_15 R_bl
Rbb_31_14 bitb_31_14 bitb_31_15 R_bl
Cb_31_14 bit_31_14 gnd C_bl
Cbb_31_14 bitb_31_14 gnd C_bl
Rb_31_15 bit_31_15 bit_31_16 R_bl
Rbb_31_15 bitb_31_15 bitb_31_16 R_bl
Cb_31_15 bit_31_15 gnd C_bl
Cbb_31_15 bitb_31_15 gnd C_bl
Rb_31_16 bit_31_16 bit_31_17 R_bl
Rbb_31_16 bitb_31_16 bitb_31_17 R_bl
Cb_31_16 bit_31_16 gnd C_bl
Cbb_31_16 bitb_31_16 gnd C_bl
Rb_31_17 bit_31_17 bit_31_18 R_bl
Rbb_31_17 bitb_31_17 bitb_31_18 R_bl
Cb_31_17 bit_31_17 gnd C_bl
Cbb_31_17 bitb_31_17 gnd C_bl
Rb_31_18 bit_31_18 bit_31_19 R_bl
Rbb_31_18 bitb_31_18 bitb_31_19 R_bl
Cb_31_18 bit_31_18 gnd C_bl
Cbb_31_18 bitb_31_18 gnd C_bl
Rb_31_19 bit_31_19 bit_31_20 R_bl
Rbb_31_19 bitb_31_19 bitb_31_20 R_bl
Cb_31_19 bit_31_19 gnd C_bl
Cbb_31_19 bitb_31_19 gnd C_bl
Rb_31_20 bit_31_20 bit_31_21 R_bl
Rbb_31_20 bitb_31_20 bitb_31_21 R_bl
Cb_31_20 bit_31_20 gnd C_bl
Cbb_31_20 bitb_31_20 gnd C_bl
Rb_31_21 bit_31_21 bit_31_22 R_bl
Rbb_31_21 bitb_31_21 bitb_31_22 R_bl
Cb_31_21 bit_31_21 gnd C_bl
Cbb_31_21 bitb_31_21 gnd C_bl
Rb_31_22 bit_31_22 bit_31_23 R_bl
Rbb_31_22 bitb_31_22 bitb_31_23 R_bl
Cb_31_22 bit_31_22 gnd C_bl
Cbb_31_22 bitb_31_22 gnd C_bl
Rb_31_23 bit_31_23 bit_31_24 R_bl
Rbb_31_23 bitb_31_23 bitb_31_24 R_bl
Cb_31_23 bit_31_23 gnd C_bl
Cbb_31_23 bitb_31_23 gnd C_bl
Rb_31_24 bit_31_24 bit_31_25 R_bl
Rbb_31_24 bitb_31_24 bitb_31_25 R_bl
Cb_31_24 bit_31_24 gnd C_bl
Cbb_31_24 bitb_31_24 gnd C_bl
Rb_31_25 bit_31_25 bit_31_26 R_bl
Rbb_31_25 bitb_31_25 bitb_31_26 R_bl
Cb_31_25 bit_31_25 gnd C_bl
Cbb_31_25 bitb_31_25 gnd C_bl
Rb_31_26 bit_31_26 bit_31_27 R_bl
Rbb_31_26 bitb_31_26 bitb_31_27 R_bl
Cb_31_26 bit_31_26 gnd C_bl
Cbb_31_26 bitb_31_26 gnd C_bl
Rb_31_27 bit_31_27 bit_31_28 R_bl
Rbb_31_27 bitb_31_27 bitb_31_28 R_bl
Cb_31_27 bit_31_27 gnd C_bl
Cbb_31_27 bitb_31_27 gnd C_bl
Rb_31_28 bit_31_28 bit_31_29 R_bl
Rbb_31_28 bitb_31_28 bitb_31_29 R_bl
Cb_31_28 bit_31_28 gnd C_bl
Cbb_31_28 bitb_31_28 gnd C_bl
Rb_31_29 bit_31_29 bit_31_30 R_bl
Rbb_31_29 bitb_31_29 bitb_31_30 R_bl
Cb_31_29 bit_31_29 gnd C_bl
Cbb_31_29 bitb_31_29 gnd C_bl
Rb_31_30 bit_31_30 bit_31_31 R_bl
Rbb_31_30 bitb_31_30 bitb_31_31 R_bl
Cb_31_30 bit_31_30 gnd C_bl
Cbb_31_30 bitb_31_30 gnd C_bl
Rb_31_31 bit_31_31 bit_31_32 R_bl
Rbb_31_31 bitb_31_31 bitb_31_32 R_bl
Cb_31_31 bit_31_31 gnd C_bl
Cbb_31_31 bitb_31_31 gnd C_bl
Rb_31_32 bit_31_32 bit_31_33 R_bl
Rbb_31_32 bitb_31_32 bitb_31_33 R_bl
Cb_31_32 bit_31_32 gnd C_bl
Cbb_31_32 bitb_31_32 gnd C_bl
Rb_31_33 bit_31_33 bit_31_34 R_bl
Rbb_31_33 bitb_31_33 bitb_31_34 R_bl
Cb_31_33 bit_31_33 gnd C_bl
Cbb_31_33 bitb_31_33 gnd C_bl
Rb_31_34 bit_31_34 bit_31_35 R_bl
Rbb_31_34 bitb_31_34 bitb_31_35 R_bl
Cb_31_34 bit_31_34 gnd C_bl
Cbb_31_34 bitb_31_34 gnd C_bl
Rb_31_35 bit_31_35 bit_31_36 R_bl
Rbb_31_35 bitb_31_35 bitb_31_36 R_bl
Cb_31_35 bit_31_35 gnd C_bl
Cbb_31_35 bitb_31_35 gnd C_bl
Rb_31_36 bit_31_36 bit_31_37 R_bl
Rbb_31_36 bitb_31_36 bitb_31_37 R_bl
Cb_31_36 bit_31_36 gnd C_bl
Cbb_31_36 bitb_31_36 gnd C_bl
Rb_31_37 bit_31_37 bit_31_38 R_bl
Rbb_31_37 bitb_31_37 bitb_31_38 R_bl
Cb_31_37 bit_31_37 gnd C_bl
Cbb_31_37 bitb_31_37 gnd C_bl
Rb_31_38 bit_31_38 bit_31_39 R_bl
Rbb_31_38 bitb_31_38 bitb_31_39 R_bl
Cb_31_38 bit_31_38 gnd C_bl
Cbb_31_38 bitb_31_38 gnd C_bl
Rb_31_39 bit_31_39 bit_31_40 R_bl
Rbb_31_39 bitb_31_39 bitb_31_40 R_bl
Cb_31_39 bit_31_39 gnd C_bl
Cbb_31_39 bitb_31_39 gnd C_bl
Rb_31_40 bit_31_40 bit_31_41 R_bl
Rbb_31_40 bitb_31_40 bitb_31_41 R_bl
Cb_31_40 bit_31_40 gnd C_bl
Cbb_31_40 bitb_31_40 gnd C_bl
Rb_31_41 bit_31_41 bit_31_42 R_bl
Rbb_31_41 bitb_31_41 bitb_31_42 R_bl
Cb_31_41 bit_31_41 gnd C_bl
Cbb_31_41 bitb_31_41 gnd C_bl
Rb_31_42 bit_31_42 bit_31_43 R_bl
Rbb_31_42 bitb_31_42 bitb_31_43 R_bl
Cb_31_42 bit_31_42 gnd C_bl
Cbb_31_42 bitb_31_42 gnd C_bl
Rb_31_43 bit_31_43 bit_31_44 R_bl
Rbb_31_43 bitb_31_43 bitb_31_44 R_bl
Cb_31_43 bit_31_43 gnd C_bl
Cbb_31_43 bitb_31_43 gnd C_bl
Rb_31_44 bit_31_44 bit_31_45 R_bl
Rbb_31_44 bitb_31_44 bitb_31_45 R_bl
Cb_31_44 bit_31_44 gnd C_bl
Cbb_31_44 bitb_31_44 gnd C_bl
Rb_31_45 bit_31_45 bit_31_46 R_bl
Rbb_31_45 bitb_31_45 bitb_31_46 R_bl
Cb_31_45 bit_31_45 gnd C_bl
Cbb_31_45 bitb_31_45 gnd C_bl
Rb_31_46 bit_31_46 bit_31_47 R_bl
Rbb_31_46 bitb_31_46 bitb_31_47 R_bl
Cb_31_46 bit_31_46 gnd C_bl
Cbb_31_46 bitb_31_46 gnd C_bl
Rb_31_47 bit_31_47 bit_31_48 R_bl
Rbb_31_47 bitb_31_47 bitb_31_48 R_bl
Cb_31_47 bit_31_47 gnd C_bl
Cbb_31_47 bitb_31_47 gnd C_bl
Rb_31_48 bit_31_48 bit_31_49 R_bl
Rbb_31_48 bitb_31_48 bitb_31_49 R_bl
Cb_31_48 bit_31_48 gnd C_bl
Cbb_31_48 bitb_31_48 gnd C_bl
Rb_31_49 bit_31_49 bit_31_50 R_bl
Rbb_31_49 bitb_31_49 bitb_31_50 R_bl
Cb_31_49 bit_31_49 gnd C_bl
Cbb_31_49 bitb_31_49 gnd C_bl
Rb_31_50 bit_31_50 bit_31_51 R_bl
Rbb_31_50 bitb_31_50 bitb_31_51 R_bl
Cb_31_50 bit_31_50 gnd C_bl
Cbb_31_50 bitb_31_50 gnd C_bl
Rb_31_51 bit_31_51 bit_31_52 R_bl
Rbb_31_51 bitb_31_51 bitb_31_52 R_bl
Cb_31_51 bit_31_51 gnd C_bl
Cbb_31_51 bitb_31_51 gnd C_bl
Rb_31_52 bit_31_52 bit_31_53 R_bl
Rbb_31_52 bitb_31_52 bitb_31_53 R_bl
Cb_31_52 bit_31_52 gnd C_bl
Cbb_31_52 bitb_31_52 gnd C_bl
Rb_31_53 bit_31_53 bit_31_54 R_bl
Rbb_31_53 bitb_31_53 bitb_31_54 R_bl
Cb_31_53 bit_31_53 gnd C_bl
Cbb_31_53 bitb_31_53 gnd C_bl
Rb_31_54 bit_31_54 bit_31_55 R_bl
Rbb_31_54 bitb_31_54 bitb_31_55 R_bl
Cb_31_54 bit_31_54 gnd C_bl
Cbb_31_54 bitb_31_54 gnd C_bl
Rb_31_55 bit_31_55 bit_31_56 R_bl
Rbb_31_55 bitb_31_55 bitb_31_56 R_bl
Cb_31_55 bit_31_55 gnd C_bl
Cbb_31_55 bitb_31_55 gnd C_bl
Rb_31_56 bit_31_56 bit_31_57 R_bl
Rbb_31_56 bitb_31_56 bitb_31_57 R_bl
Cb_31_56 bit_31_56 gnd C_bl
Cbb_31_56 bitb_31_56 gnd C_bl
Rb_31_57 bit_31_57 bit_31_58 R_bl
Rbb_31_57 bitb_31_57 bitb_31_58 R_bl
Cb_31_57 bit_31_57 gnd C_bl
Cbb_31_57 bitb_31_57 gnd C_bl
Rb_31_58 bit_31_58 bit_31_59 R_bl
Rbb_31_58 bitb_31_58 bitb_31_59 R_bl
Cb_31_58 bit_31_58 gnd C_bl
Cbb_31_58 bitb_31_58 gnd C_bl
Rb_31_59 bit_31_59 bit_31_60 R_bl
Rbb_31_59 bitb_31_59 bitb_31_60 R_bl
Cb_31_59 bit_31_59 gnd C_bl
Cbb_31_59 bitb_31_59 gnd C_bl
Rb_31_60 bit_31_60 bit_31_61 R_bl
Rbb_31_60 bitb_31_60 bitb_31_61 R_bl
Cb_31_60 bit_31_60 gnd C_bl
Cbb_31_60 bitb_31_60 gnd C_bl
Rb_31_61 bit_31_61 bit_31_62 R_bl
Rbb_31_61 bitb_31_61 bitb_31_62 R_bl
Cb_31_61 bit_31_61 gnd C_bl
Cbb_31_61 bitb_31_61 gnd C_bl
Rb_31_62 bit_31_62 bit_31_63 R_bl
Rbb_31_62 bitb_31_62 bitb_31_63 R_bl
Cb_31_62 bit_31_62 gnd C_bl
Cbb_31_62 bitb_31_62 gnd C_bl
Rb_31_63 bit_31_63 bit_31_64 R_bl
Rbb_31_63 bitb_31_63 bitb_31_64 R_bl
Cb_31_63 bit_31_63 gnd C_bl
Cbb_31_63 bitb_31_63 gnd C_bl
Rb_31_64 bit_31_64 bit_31_65 R_bl
Rbb_31_64 bitb_31_64 bitb_31_65 R_bl
Cb_31_64 bit_31_64 gnd C_bl
Cbb_31_64 bitb_31_64 gnd C_bl
Rb_31_65 bit_31_65 bit_31_66 R_bl
Rbb_31_65 bitb_31_65 bitb_31_66 R_bl
Cb_31_65 bit_31_65 gnd C_bl
Cbb_31_65 bitb_31_65 gnd C_bl
Rb_31_66 bit_31_66 bit_31_67 R_bl
Rbb_31_66 bitb_31_66 bitb_31_67 R_bl
Cb_31_66 bit_31_66 gnd C_bl
Cbb_31_66 bitb_31_66 gnd C_bl
Rb_31_67 bit_31_67 bit_31_68 R_bl
Rbb_31_67 bitb_31_67 bitb_31_68 R_bl
Cb_31_67 bit_31_67 gnd C_bl
Cbb_31_67 bitb_31_67 gnd C_bl
Rb_31_68 bit_31_68 bit_31_69 R_bl
Rbb_31_68 bitb_31_68 bitb_31_69 R_bl
Cb_31_68 bit_31_68 gnd C_bl
Cbb_31_68 bitb_31_68 gnd C_bl
Rb_31_69 bit_31_69 bit_31_70 R_bl
Rbb_31_69 bitb_31_69 bitb_31_70 R_bl
Cb_31_69 bit_31_69 gnd C_bl
Cbb_31_69 bitb_31_69 gnd C_bl
Rb_31_70 bit_31_70 bit_31_71 R_bl
Rbb_31_70 bitb_31_70 bitb_31_71 R_bl
Cb_31_70 bit_31_70 gnd C_bl
Cbb_31_70 bitb_31_70 gnd C_bl
Rb_31_71 bit_31_71 bit_31_72 R_bl
Rbb_31_71 bitb_31_71 bitb_31_72 R_bl
Cb_31_71 bit_31_71 gnd C_bl
Cbb_31_71 bitb_31_71 gnd C_bl
Rb_31_72 bit_31_72 bit_31_73 R_bl
Rbb_31_72 bitb_31_72 bitb_31_73 R_bl
Cb_31_72 bit_31_72 gnd C_bl
Cbb_31_72 bitb_31_72 gnd C_bl
Rb_31_73 bit_31_73 bit_31_74 R_bl
Rbb_31_73 bitb_31_73 bitb_31_74 R_bl
Cb_31_73 bit_31_73 gnd C_bl
Cbb_31_73 bitb_31_73 gnd C_bl
Rb_31_74 bit_31_74 bit_31_75 R_bl
Rbb_31_74 bitb_31_74 bitb_31_75 R_bl
Cb_31_74 bit_31_74 gnd C_bl
Cbb_31_74 bitb_31_74 gnd C_bl
Rb_31_75 bit_31_75 bit_31_76 R_bl
Rbb_31_75 bitb_31_75 bitb_31_76 R_bl
Cb_31_75 bit_31_75 gnd C_bl
Cbb_31_75 bitb_31_75 gnd C_bl
Rb_31_76 bit_31_76 bit_31_77 R_bl
Rbb_31_76 bitb_31_76 bitb_31_77 R_bl
Cb_31_76 bit_31_76 gnd C_bl
Cbb_31_76 bitb_31_76 gnd C_bl
Rb_31_77 bit_31_77 bit_31_78 R_bl
Rbb_31_77 bitb_31_77 bitb_31_78 R_bl
Cb_31_77 bit_31_77 gnd C_bl
Cbb_31_77 bitb_31_77 gnd C_bl
Rb_31_78 bit_31_78 bit_31_79 R_bl
Rbb_31_78 bitb_31_78 bitb_31_79 R_bl
Cb_31_78 bit_31_78 gnd C_bl
Cbb_31_78 bitb_31_78 gnd C_bl
Rb_31_79 bit_31_79 bit_31_80 R_bl
Rbb_31_79 bitb_31_79 bitb_31_80 R_bl
Cb_31_79 bit_31_79 gnd C_bl
Cbb_31_79 bitb_31_79 gnd C_bl
Rb_31_80 bit_31_80 bit_31_81 R_bl
Rbb_31_80 bitb_31_80 bitb_31_81 R_bl
Cb_31_80 bit_31_80 gnd C_bl
Cbb_31_80 bitb_31_80 gnd C_bl
Rb_31_81 bit_31_81 bit_31_82 R_bl
Rbb_31_81 bitb_31_81 bitb_31_82 R_bl
Cb_31_81 bit_31_81 gnd C_bl
Cbb_31_81 bitb_31_81 gnd C_bl
Rb_31_82 bit_31_82 bit_31_83 R_bl
Rbb_31_82 bitb_31_82 bitb_31_83 R_bl
Cb_31_82 bit_31_82 gnd C_bl
Cbb_31_82 bitb_31_82 gnd C_bl
Rb_31_83 bit_31_83 bit_31_84 R_bl
Rbb_31_83 bitb_31_83 bitb_31_84 R_bl
Cb_31_83 bit_31_83 gnd C_bl
Cbb_31_83 bitb_31_83 gnd C_bl
Rb_31_84 bit_31_84 bit_31_85 R_bl
Rbb_31_84 bitb_31_84 bitb_31_85 R_bl
Cb_31_84 bit_31_84 gnd C_bl
Cbb_31_84 bitb_31_84 gnd C_bl
Rb_31_85 bit_31_85 bit_31_86 R_bl
Rbb_31_85 bitb_31_85 bitb_31_86 R_bl
Cb_31_85 bit_31_85 gnd C_bl
Cbb_31_85 bitb_31_85 gnd C_bl
Rb_31_86 bit_31_86 bit_31_87 R_bl
Rbb_31_86 bitb_31_86 bitb_31_87 R_bl
Cb_31_86 bit_31_86 gnd C_bl
Cbb_31_86 bitb_31_86 gnd C_bl
Rb_31_87 bit_31_87 bit_31_88 R_bl
Rbb_31_87 bitb_31_87 bitb_31_88 R_bl
Cb_31_87 bit_31_87 gnd C_bl
Cbb_31_87 bitb_31_87 gnd C_bl
Rb_31_88 bit_31_88 bit_31_89 R_bl
Rbb_31_88 bitb_31_88 bitb_31_89 R_bl
Cb_31_88 bit_31_88 gnd C_bl
Cbb_31_88 bitb_31_88 gnd C_bl
Rb_31_89 bit_31_89 bit_31_90 R_bl
Rbb_31_89 bitb_31_89 bitb_31_90 R_bl
Cb_31_89 bit_31_89 gnd C_bl
Cbb_31_89 bitb_31_89 gnd C_bl
Rb_31_90 bit_31_90 bit_31_91 R_bl
Rbb_31_90 bitb_31_90 bitb_31_91 R_bl
Cb_31_90 bit_31_90 gnd C_bl
Cbb_31_90 bitb_31_90 gnd C_bl
Rb_31_91 bit_31_91 bit_31_92 R_bl
Rbb_31_91 bitb_31_91 bitb_31_92 R_bl
Cb_31_91 bit_31_91 gnd C_bl
Cbb_31_91 bitb_31_91 gnd C_bl
Rb_31_92 bit_31_92 bit_31_93 R_bl
Rbb_31_92 bitb_31_92 bitb_31_93 R_bl
Cb_31_92 bit_31_92 gnd C_bl
Cbb_31_92 bitb_31_92 gnd C_bl
Rb_31_93 bit_31_93 bit_31_94 R_bl
Rbb_31_93 bitb_31_93 bitb_31_94 R_bl
Cb_31_93 bit_31_93 gnd C_bl
Cbb_31_93 bitb_31_93 gnd C_bl
Rb_31_94 bit_31_94 bit_31_95 R_bl
Rbb_31_94 bitb_31_94 bitb_31_95 R_bl
Cb_31_94 bit_31_94 gnd C_bl
Cbb_31_94 bitb_31_94 gnd C_bl
Rb_31_95 bit_31_95 bit_31_96 R_bl
Rbb_31_95 bitb_31_95 bitb_31_96 R_bl
Cb_31_95 bit_31_95 gnd C_bl
Cbb_31_95 bitb_31_95 gnd C_bl
Rb_31_96 bit_31_96 bit_31_97 R_bl
Rbb_31_96 bitb_31_96 bitb_31_97 R_bl
Cb_31_96 bit_31_96 gnd C_bl
Cbb_31_96 bitb_31_96 gnd C_bl
Rb_31_97 bit_31_97 bit_31_98 R_bl
Rbb_31_97 bitb_31_97 bitb_31_98 R_bl
Cb_31_97 bit_31_97 gnd C_bl
Cbb_31_97 bitb_31_97 gnd C_bl
Rb_31_98 bit_31_98 bit_31_99 R_bl
Rbb_31_98 bitb_31_98 bitb_31_99 R_bl
Cb_31_98 bit_31_98 gnd C_bl
Cbb_31_98 bitb_31_98 gnd C_bl
Rb_31_99 bit_31_99 bit_31_100 R_bl
Rbb_31_99 bitb_31_99 bitb_31_100 R_bl
Cb_31_99 bit_31_99 gnd C_bl
Cbb_31_99 bitb_31_99 gnd C_bl
Rb_32_0 bit_32_0 bit_32_1 R_bl
Rbb_32_0 bitb_32_0 bitb_32_1 R_bl
Cb_32_0 bit_32_0 gnd C_bl
Cbb_32_0 bitb_32_0 gnd C_bl
Rb_32_1 bit_32_1 bit_32_2 R_bl
Rbb_32_1 bitb_32_1 bitb_32_2 R_bl
Cb_32_1 bit_32_1 gnd C_bl
Cbb_32_1 bitb_32_1 gnd C_bl
Rb_32_2 bit_32_2 bit_32_3 R_bl
Rbb_32_2 bitb_32_2 bitb_32_3 R_bl
Cb_32_2 bit_32_2 gnd C_bl
Cbb_32_2 bitb_32_2 gnd C_bl
Rb_32_3 bit_32_3 bit_32_4 R_bl
Rbb_32_3 bitb_32_3 bitb_32_4 R_bl
Cb_32_3 bit_32_3 gnd C_bl
Cbb_32_3 bitb_32_3 gnd C_bl
Rb_32_4 bit_32_4 bit_32_5 R_bl
Rbb_32_4 bitb_32_4 bitb_32_5 R_bl
Cb_32_4 bit_32_4 gnd C_bl
Cbb_32_4 bitb_32_4 gnd C_bl
Rb_32_5 bit_32_5 bit_32_6 R_bl
Rbb_32_5 bitb_32_5 bitb_32_6 R_bl
Cb_32_5 bit_32_5 gnd C_bl
Cbb_32_5 bitb_32_5 gnd C_bl
Rb_32_6 bit_32_6 bit_32_7 R_bl
Rbb_32_6 bitb_32_6 bitb_32_7 R_bl
Cb_32_6 bit_32_6 gnd C_bl
Cbb_32_6 bitb_32_6 gnd C_bl
Rb_32_7 bit_32_7 bit_32_8 R_bl
Rbb_32_7 bitb_32_7 bitb_32_8 R_bl
Cb_32_7 bit_32_7 gnd C_bl
Cbb_32_7 bitb_32_7 gnd C_bl
Rb_32_8 bit_32_8 bit_32_9 R_bl
Rbb_32_8 bitb_32_8 bitb_32_9 R_bl
Cb_32_8 bit_32_8 gnd C_bl
Cbb_32_8 bitb_32_8 gnd C_bl
Rb_32_9 bit_32_9 bit_32_10 R_bl
Rbb_32_9 bitb_32_9 bitb_32_10 R_bl
Cb_32_9 bit_32_9 gnd C_bl
Cbb_32_9 bitb_32_9 gnd C_bl
Rb_32_10 bit_32_10 bit_32_11 R_bl
Rbb_32_10 bitb_32_10 bitb_32_11 R_bl
Cb_32_10 bit_32_10 gnd C_bl
Cbb_32_10 bitb_32_10 gnd C_bl
Rb_32_11 bit_32_11 bit_32_12 R_bl
Rbb_32_11 bitb_32_11 bitb_32_12 R_bl
Cb_32_11 bit_32_11 gnd C_bl
Cbb_32_11 bitb_32_11 gnd C_bl
Rb_32_12 bit_32_12 bit_32_13 R_bl
Rbb_32_12 bitb_32_12 bitb_32_13 R_bl
Cb_32_12 bit_32_12 gnd C_bl
Cbb_32_12 bitb_32_12 gnd C_bl
Rb_32_13 bit_32_13 bit_32_14 R_bl
Rbb_32_13 bitb_32_13 bitb_32_14 R_bl
Cb_32_13 bit_32_13 gnd C_bl
Cbb_32_13 bitb_32_13 gnd C_bl
Rb_32_14 bit_32_14 bit_32_15 R_bl
Rbb_32_14 bitb_32_14 bitb_32_15 R_bl
Cb_32_14 bit_32_14 gnd C_bl
Cbb_32_14 bitb_32_14 gnd C_bl
Rb_32_15 bit_32_15 bit_32_16 R_bl
Rbb_32_15 bitb_32_15 bitb_32_16 R_bl
Cb_32_15 bit_32_15 gnd C_bl
Cbb_32_15 bitb_32_15 gnd C_bl
Rb_32_16 bit_32_16 bit_32_17 R_bl
Rbb_32_16 bitb_32_16 bitb_32_17 R_bl
Cb_32_16 bit_32_16 gnd C_bl
Cbb_32_16 bitb_32_16 gnd C_bl
Rb_32_17 bit_32_17 bit_32_18 R_bl
Rbb_32_17 bitb_32_17 bitb_32_18 R_bl
Cb_32_17 bit_32_17 gnd C_bl
Cbb_32_17 bitb_32_17 gnd C_bl
Rb_32_18 bit_32_18 bit_32_19 R_bl
Rbb_32_18 bitb_32_18 bitb_32_19 R_bl
Cb_32_18 bit_32_18 gnd C_bl
Cbb_32_18 bitb_32_18 gnd C_bl
Rb_32_19 bit_32_19 bit_32_20 R_bl
Rbb_32_19 bitb_32_19 bitb_32_20 R_bl
Cb_32_19 bit_32_19 gnd C_bl
Cbb_32_19 bitb_32_19 gnd C_bl
Rb_32_20 bit_32_20 bit_32_21 R_bl
Rbb_32_20 bitb_32_20 bitb_32_21 R_bl
Cb_32_20 bit_32_20 gnd C_bl
Cbb_32_20 bitb_32_20 gnd C_bl
Rb_32_21 bit_32_21 bit_32_22 R_bl
Rbb_32_21 bitb_32_21 bitb_32_22 R_bl
Cb_32_21 bit_32_21 gnd C_bl
Cbb_32_21 bitb_32_21 gnd C_bl
Rb_32_22 bit_32_22 bit_32_23 R_bl
Rbb_32_22 bitb_32_22 bitb_32_23 R_bl
Cb_32_22 bit_32_22 gnd C_bl
Cbb_32_22 bitb_32_22 gnd C_bl
Rb_32_23 bit_32_23 bit_32_24 R_bl
Rbb_32_23 bitb_32_23 bitb_32_24 R_bl
Cb_32_23 bit_32_23 gnd C_bl
Cbb_32_23 bitb_32_23 gnd C_bl
Rb_32_24 bit_32_24 bit_32_25 R_bl
Rbb_32_24 bitb_32_24 bitb_32_25 R_bl
Cb_32_24 bit_32_24 gnd C_bl
Cbb_32_24 bitb_32_24 gnd C_bl
Rb_32_25 bit_32_25 bit_32_26 R_bl
Rbb_32_25 bitb_32_25 bitb_32_26 R_bl
Cb_32_25 bit_32_25 gnd C_bl
Cbb_32_25 bitb_32_25 gnd C_bl
Rb_32_26 bit_32_26 bit_32_27 R_bl
Rbb_32_26 bitb_32_26 bitb_32_27 R_bl
Cb_32_26 bit_32_26 gnd C_bl
Cbb_32_26 bitb_32_26 gnd C_bl
Rb_32_27 bit_32_27 bit_32_28 R_bl
Rbb_32_27 bitb_32_27 bitb_32_28 R_bl
Cb_32_27 bit_32_27 gnd C_bl
Cbb_32_27 bitb_32_27 gnd C_bl
Rb_32_28 bit_32_28 bit_32_29 R_bl
Rbb_32_28 bitb_32_28 bitb_32_29 R_bl
Cb_32_28 bit_32_28 gnd C_bl
Cbb_32_28 bitb_32_28 gnd C_bl
Rb_32_29 bit_32_29 bit_32_30 R_bl
Rbb_32_29 bitb_32_29 bitb_32_30 R_bl
Cb_32_29 bit_32_29 gnd C_bl
Cbb_32_29 bitb_32_29 gnd C_bl
Rb_32_30 bit_32_30 bit_32_31 R_bl
Rbb_32_30 bitb_32_30 bitb_32_31 R_bl
Cb_32_30 bit_32_30 gnd C_bl
Cbb_32_30 bitb_32_30 gnd C_bl
Rb_32_31 bit_32_31 bit_32_32 R_bl
Rbb_32_31 bitb_32_31 bitb_32_32 R_bl
Cb_32_31 bit_32_31 gnd C_bl
Cbb_32_31 bitb_32_31 gnd C_bl
Rb_32_32 bit_32_32 bit_32_33 R_bl
Rbb_32_32 bitb_32_32 bitb_32_33 R_bl
Cb_32_32 bit_32_32 gnd C_bl
Cbb_32_32 bitb_32_32 gnd C_bl
Rb_32_33 bit_32_33 bit_32_34 R_bl
Rbb_32_33 bitb_32_33 bitb_32_34 R_bl
Cb_32_33 bit_32_33 gnd C_bl
Cbb_32_33 bitb_32_33 gnd C_bl
Rb_32_34 bit_32_34 bit_32_35 R_bl
Rbb_32_34 bitb_32_34 bitb_32_35 R_bl
Cb_32_34 bit_32_34 gnd C_bl
Cbb_32_34 bitb_32_34 gnd C_bl
Rb_32_35 bit_32_35 bit_32_36 R_bl
Rbb_32_35 bitb_32_35 bitb_32_36 R_bl
Cb_32_35 bit_32_35 gnd C_bl
Cbb_32_35 bitb_32_35 gnd C_bl
Rb_32_36 bit_32_36 bit_32_37 R_bl
Rbb_32_36 bitb_32_36 bitb_32_37 R_bl
Cb_32_36 bit_32_36 gnd C_bl
Cbb_32_36 bitb_32_36 gnd C_bl
Rb_32_37 bit_32_37 bit_32_38 R_bl
Rbb_32_37 bitb_32_37 bitb_32_38 R_bl
Cb_32_37 bit_32_37 gnd C_bl
Cbb_32_37 bitb_32_37 gnd C_bl
Rb_32_38 bit_32_38 bit_32_39 R_bl
Rbb_32_38 bitb_32_38 bitb_32_39 R_bl
Cb_32_38 bit_32_38 gnd C_bl
Cbb_32_38 bitb_32_38 gnd C_bl
Rb_32_39 bit_32_39 bit_32_40 R_bl
Rbb_32_39 bitb_32_39 bitb_32_40 R_bl
Cb_32_39 bit_32_39 gnd C_bl
Cbb_32_39 bitb_32_39 gnd C_bl
Rb_32_40 bit_32_40 bit_32_41 R_bl
Rbb_32_40 bitb_32_40 bitb_32_41 R_bl
Cb_32_40 bit_32_40 gnd C_bl
Cbb_32_40 bitb_32_40 gnd C_bl
Rb_32_41 bit_32_41 bit_32_42 R_bl
Rbb_32_41 bitb_32_41 bitb_32_42 R_bl
Cb_32_41 bit_32_41 gnd C_bl
Cbb_32_41 bitb_32_41 gnd C_bl
Rb_32_42 bit_32_42 bit_32_43 R_bl
Rbb_32_42 bitb_32_42 bitb_32_43 R_bl
Cb_32_42 bit_32_42 gnd C_bl
Cbb_32_42 bitb_32_42 gnd C_bl
Rb_32_43 bit_32_43 bit_32_44 R_bl
Rbb_32_43 bitb_32_43 bitb_32_44 R_bl
Cb_32_43 bit_32_43 gnd C_bl
Cbb_32_43 bitb_32_43 gnd C_bl
Rb_32_44 bit_32_44 bit_32_45 R_bl
Rbb_32_44 bitb_32_44 bitb_32_45 R_bl
Cb_32_44 bit_32_44 gnd C_bl
Cbb_32_44 bitb_32_44 gnd C_bl
Rb_32_45 bit_32_45 bit_32_46 R_bl
Rbb_32_45 bitb_32_45 bitb_32_46 R_bl
Cb_32_45 bit_32_45 gnd C_bl
Cbb_32_45 bitb_32_45 gnd C_bl
Rb_32_46 bit_32_46 bit_32_47 R_bl
Rbb_32_46 bitb_32_46 bitb_32_47 R_bl
Cb_32_46 bit_32_46 gnd C_bl
Cbb_32_46 bitb_32_46 gnd C_bl
Rb_32_47 bit_32_47 bit_32_48 R_bl
Rbb_32_47 bitb_32_47 bitb_32_48 R_bl
Cb_32_47 bit_32_47 gnd C_bl
Cbb_32_47 bitb_32_47 gnd C_bl
Rb_32_48 bit_32_48 bit_32_49 R_bl
Rbb_32_48 bitb_32_48 bitb_32_49 R_bl
Cb_32_48 bit_32_48 gnd C_bl
Cbb_32_48 bitb_32_48 gnd C_bl
Rb_32_49 bit_32_49 bit_32_50 R_bl
Rbb_32_49 bitb_32_49 bitb_32_50 R_bl
Cb_32_49 bit_32_49 gnd C_bl
Cbb_32_49 bitb_32_49 gnd C_bl
Rb_32_50 bit_32_50 bit_32_51 R_bl
Rbb_32_50 bitb_32_50 bitb_32_51 R_bl
Cb_32_50 bit_32_50 gnd C_bl
Cbb_32_50 bitb_32_50 gnd C_bl
Rb_32_51 bit_32_51 bit_32_52 R_bl
Rbb_32_51 bitb_32_51 bitb_32_52 R_bl
Cb_32_51 bit_32_51 gnd C_bl
Cbb_32_51 bitb_32_51 gnd C_bl
Rb_32_52 bit_32_52 bit_32_53 R_bl
Rbb_32_52 bitb_32_52 bitb_32_53 R_bl
Cb_32_52 bit_32_52 gnd C_bl
Cbb_32_52 bitb_32_52 gnd C_bl
Rb_32_53 bit_32_53 bit_32_54 R_bl
Rbb_32_53 bitb_32_53 bitb_32_54 R_bl
Cb_32_53 bit_32_53 gnd C_bl
Cbb_32_53 bitb_32_53 gnd C_bl
Rb_32_54 bit_32_54 bit_32_55 R_bl
Rbb_32_54 bitb_32_54 bitb_32_55 R_bl
Cb_32_54 bit_32_54 gnd C_bl
Cbb_32_54 bitb_32_54 gnd C_bl
Rb_32_55 bit_32_55 bit_32_56 R_bl
Rbb_32_55 bitb_32_55 bitb_32_56 R_bl
Cb_32_55 bit_32_55 gnd C_bl
Cbb_32_55 bitb_32_55 gnd C_bl
Rb_32_56 bit_32_56 bit_32_57 R_bl
Rbb_32_56 bitb_32_56 bitb_32_57 R_bl
Cb_32_56 bit_32_56 gnd C_bl
Cbb_32_56 bitb_32_56 gnd C_bl
Rb_32_57 bit_32_57 bit_32_58 R_bl
Rbb_32_57 bitb_32_57 bitb_32_58 R_bl
Cb_32_57 bit_32_57 gnd C_bl
Cbb_32_57 bitb_32_57 gnd C_bl
Rb_32_58 bit_32_58 bit_32_59 R_bl
Rbb_32_58 bitb_32_58 bitb_32_59 R_bl
Cb_32_58 bit_32_58 gnd C_bl
Cbb_32_58 bitb_32_58 gnd C_bl
Rb_32_59 bit_32_59 bit_32_60 R_bl
Rbb_32_59 bitb_32_59 bitb_32_60 R_bl
Cb_32_59 bit_32_59 gnd C_bl
Cbb_32_59 bitb_32_59 gnd C_bl
Rb_32_60 bit_32_60 bit_32_61 R_bl
Rbb_32_60 bitb_32_60 bitb_32_61 R_bl
Cb_32_60 bit_32_60 gnd C_bl
Cbb_32_60 bitb_32_60 gnd C_bl
Rb_32_61 bit_32_61 bit_32_62 R_bl
Rbb_32_61 bitb_32_61 bitb_32_62 R_bl
Cb_32_61 bit_32_61 gnd C_bl
Cbb_32_61 bitb_32_61 gnd C_bl
Rb_32_62 bit_32_62 bit_32_63 R_bl
Rbb_32_62 bitb_32_62 bitb_32_63 R_bl
Cb_32_62 bit_32_62 gnd C_bl
Cbb_32_62 bitb_32_62 gnd C_bl
Rb_32_63 bit_32_63 bit_32_64 R_bl
Rbb_32_63 bitb_32_63 bitb_32_64 R_bl
Cb_32_63 bit_32_63 gnd C_bl
Cbb_32_63 bitb_32_63 gnd C_bl
Rb_32_64 bit_32_64 bit_32_65 R_bl
Rbb_32_64 bitb_32_64 bitb_32_65 R_bl
Cb_32_64 bit_32_64 gnd C_bl
Cbb_32_64 bitb_32_64 gnd C_bl
Rb_32_65 bit_32_65 bit_32_66 R_bl
Rbb_32_65 bitb_32_65 bitb_32_66 R_bl
Cb_32_65 bit_32_65 gnd C_bl
Cbb_32_65 bitb_32_65 gnd C_bl
Rb_32_66 bit_32_66 bit_32_67 R_bl
Rbb_32_66 bitb_32_66 bitb_32_67 R_bl
Cb_32_66 bit_32_66 gnd C_bl
Cbb_32_66 bitb_32_66 gnd C_bl
Rb_32_67 bit_32_67 bit_32_68 R_bl
Rbb_32_67 bitb_32_67 bitb_32_68 R_bl
Cb_32_67 bit_32_67 gnd C_bl
Cbb_32_67 bitb_32_67 gnd C_bl
Rb_32_68 bit_32_68 bit_32_69 R_bl
Rbb_32_68 bitb_32_68 bitb_32_69 R_bl
Cb_32_68 bit_32_68 gnd C_bl
Cbb_32_68 bitb_32_68 gnd C_bl
Rb_32_69 bit_32_69 bit_32_70 R_bl
Rbb_32_69 bitb_32_69 bitb_32_70 R_bl
Cb_32_69 bit_32_69 gnd C_bl
Cbb_32_69 bitb_32_69 gnd C_bl
Rb_32_70 bit_32_70 bit_32_71 R_bl
Rbb_32_70 bitb_32_70 bitb_32_71 R_bl
Cb_32_70 bit_32_70 gnd C_bl
Cbb_32_70 bitb_32_70 gnd C_bl
Rb_32_71 bit_32_71 bit_32_72 R_bl
Rbb_32_71 bitb_32_71 bitb_32_72 R_bl
Cb_32_71 bit_32_71 gnd C_bl
Cbb_32_71 bitb_32_71 gnd C_bl
Rb_32_72 bit_32_72 bit_32_73 R_bl
Rbb_32_72 bitb_32_72 bitb_32_73 R_bl
Cb_32_72 bit_32_72 gnd C_bl
Cbb_32_72 bitb_32_72 gnd C_bl
Rb_32_73 bit_32_73 bit_32_74 R_bl
Rbb_32_73 bitb_32_73 bitb_32_74 R_bl
Cb_32_73 bit_32_73 gnd C_bl
Cbb_32_73 bitb_32_73 gnd C_bl
Rb_32_74 bit_32_74 bit_32_75 R_bl
Rbb_32_74 bitb_32_74 bitb_32_75 R_bl
Cb_32_74 bit_32_74 gnd C_bl
Cbb_32_74 bitb_32_74 gnd C_bl
Rb_32_75 bit_32_75 bit_32_76 R_bl
Rbb_32_75 bitb_32_75 bitb_32_76 R_bl
Cb_32_75 bit_32_75 gnd C_bl
Cbb_32_75 bitb_32_75 gnd C_bl
Rb_32_76 bit_32_76 bit_32_77 R_bl
Rbb_32_76 bitb_32_76 bitb_32_77 R_bl
Cb_32_76 bit_32_76 gnd C_bl
Cbb_32_76 bitb_32_76 gnd C_bl
Rb_32_77 bit_32_77 bit_32_78 R_bl
Rbb_32_77 bitb_32_77 bitb_32_78 R_bl
Cb_32_77 bit_32_77 gnd C_bl
Cbb_32_77 bitb_32_77 gnd C_bl
Rb_32_78 bit_32_78 bit_32_79 R_bl
Rbb_32_78 bitb_32_78 bitb_32_79 R_bl
Cb_32_78 bit_32_78 gnd C_bl
Cbb_32_78 bitb_32_78 gnd C_bl
Rb_32_79 bit_32_79 bit_32_80 R_bl
Rbb_32_79 bitb_32_79 bitb_32_80 R_bl
Cb_32_79 bit_32_79 gnd C_bl
Cbb_32_79 bitb_32_79 gnd C_bl
Rb_32_80 bit_32_80 bit_32_81 R_bl
Rbb_32_80 bitb_32_80 bitb_32_81 R_bl
Cb_32_80 bit_32_80 gnd C_bl
Cbb_32_80 bitb_32_80 gnd C_bl
Rb_32_81 bit_32_81 bit_32_82 R_bl
Rbb_32_81 bitb_32_81 bitb_32_82 R_bl
Cb_32_81 bit_32_81 gnd C_bl
Cbb_32_81 bitb_32_81 gnd C_bl
Rb_32_82 bit_32_82 bit_32_83 R_bl
Rbb_32_82 bitb_32_82 bitb_32_83 R_bl
Cb_32_82 bit_32_82 gnd C_bl
Cbb_32_82 bitb_32_82 gnd C_bl
Rb_32_83 bit_32_83 bit_32_84 R_bl
Rbb_32_83 bitb_32_83 bitb_32_84 R_bl
Cb_32_83 bit_32_83 gnd C_bl
Cbb_32_83 bitb_32_83 gnd C_bl
Rb_32_84 bit_32_84 bit_32_85 R_bl
Rbb_32_84 bitb_32_84 bitb_32_85 R_bl
Cb_32_84 bit_32_84 gnd C_bl
Cbb_32_84 bitb_32_84 gnd C_bl
Rb_32_85 bit_32_85 bit_32_86 R_bl
Rbb_32_85 bitb_32_85 bitb_32_86 R_bl
Cb_32_85 bit_32_85 gnd C_bl
Cbb_32_85 bitb_32_85 gnd C_bl
Rb_32_86 bit_32_86 bit_32_87 R_bl
Rbb_32_86 bitb_32_86 bitb_32_87 R_bl
Cb_32_86 bit_32_86 gnd C_bl
Cbb_32_86 bitb_32_86 gnd C_bl
Rb_32_87 bit_32_87 bit_32_88 R_bl
Rbb_32_87 bitb_32_87 bitb_32_88 R_bl
Cb_32_87 bit_32_87 gnd C_bl
Cbb_32_87 bitb_32_87 gnd C_bl
Rb_32_88 bit_32_88 bit_32_89 R_bl
Rbb_32_88 bitb_32_88 bitb_32_89 R_bl
Cb_32_88 bit_32_88 gnd C_bl
Cbb_32_88 bitb_32_88 gnd C_bl
Rb_32_89 bit_32_89 bit_32_90 R_bl
Rbb_32_89 bitb_32_89 bitb_32_90 R_bl
Cb_32_89 bit_32_89 gnd C_bl
Cbb_32_89 bitb_32_89 gnd C_bl
Rb_32_90 bit_32_90 bit_32_91 R_bl
Rbb_32_90 bitb_32_90 bitb_32_91 R_bl
Cb_32_90 bit_32_90 gnd C_bl
Cbb_32_90 bitb_32_90 gnd C_bl
Rb_32_91 bit_32_91 bit_32_92 R_bl
Rbb_32_91 bitb_32_91 bitb_32_92 R_bl
Cb_32_91 bit_32_91 gnd C_bl
Cbb_32_91 bitb_32_91 gnd C_bl
Rb_32_92 bit_32_92 bit_32_93 R_bl
Rbb_32_92 bitb_32_92 bitb_32_93 R_bl
Cb_32_92 bit_32_92 gnd C_bl
Cbb_32_92 bitb_32_92 gnd C_bl
Rb_32_93 bit_32_93 bit_32_94 R_bl
Rbb_32_93 bitb_32_93 bitb_32_94 R_bl
Cb_32_93 bit_32_93 gnd C_bl
Cbb_32_93 bitb_32_93 gnd C_bl
Rb_32_94 bit_32_94 bit_32_95 R_bl
Rbb_32_94 bitb_32_94 bitb_32_95 R_bl
Cb_32_94 bit_32_94 gnd C_bl
Cbb_32_94 bitb_32_94 gnd C_bl
Rb_32_95 bit_32_95 bit_32_96 R_bl
Rbb_32_95 bitb_32_95 bitb_32_96 R_bl
Cb_32_95 bit_32_95 gnd C_bl
Cbb_32_95 bitb_32_95 gnd C_bl
Rb_32_96 bit_32_96 bit_32_97 R_bl
Rbb_32_96 bitb_32_96 bitb_32_97 R_bl
Cb_32_96 bit_32_96 gnd C_bl
Cbb_32_96 bitb_32_96 gnd C_bl
Rb_32_97 bit_32_97 bit_32_98 R_bl
Rbb_32_97 bitb_32_97 bitb_32_98 R_bl
Cb_32_97 bit_32_97 gnd C_bl
Cbb_32_97 bitb_32_97 gnd C_bl
Rb_32_98 bit_32_98 bit_32_99 R_bl
Rbb_32_98 bitb_32_98 bitb_32_99 R_bl
Cb_32_98 bit_32_98 gnd C_bl
Cbb_32_98 bitb_32_98 gnd C_bl
Rb_32_99 bit_32_99 bit_32_100 R_bl
Rbb_32_99 bitb_32_99 bitb_32_100 R_bl
Cb_32_99 bit_32_99 gnd C_bl
Cbb_32_99 bitb_32_99 gnd C_bl
Rb_33_0 bit_33_0 bit_33_1 R_bl
Rbb_33_0 bitb_33_0 bitb_33_1 R_bl
Cb_33_0 bit_33_0 gnd C_bl
Cbb_33_0 bitb_33_0 gnd C_bl
Rb_33_1 bit_33_1 bit_33_2 R_bl
Rbb_33_1 bitb_33_1 bitb_33_2 R_bl
Cb_33_1 bit_33_1 gnd C_bl
Cbb_33_1 bitb_33_1 gnd C_bl
Rb_33_2 bit_33_2 bit_33_3 R_bl
Rbb_33_2 bitb_33_2 bitb_33_3 R_bl
Cb_33_2 bit_33_2 gnd C_bl
Cbb_33_2 bitb_33_2 gnd C_bl
Rb_33_3 bit_33_3 bit_33_4 R_bl
Rbb_33_3 bitb_33_3 bitb_33_4 R_bl
Cb_33_3 bit_33_3 gnd C_bl
Cbb_33_3 bitb_33_3 gnd C_bl
Rb_33_4 bit_33_4 bit_33_5 R_bl
Rbb_33_4 bitb_33_4 bitb_33_5 R_bl
Cb_33_4 bit_33_4 gnd C_bl
Cbb_33_4 bitb_33_4 gnd C_bl
Rb_33_5 bit_33_5 bit_33_6 R_bl
Rbb_33_5 bitb_33_5 bitb_33_6 R_bl
Cb_33_5 bit_33_5 gnd C_bl
Cbb_33_5 bitb_33_5 gnd C_bl
Rb_33_6 bit_33_6 bit_33_7 R_bl
Rbb_33_6 bitb_33_6 bitb_33_7 R_bl
Cb_33_6 bit_33_6 gnd C_bl
Cbb_33_6 bitb_33_6 gnd C_bl
Rb_33_7 bit_33_7 bit_33_8 R_bl
Rbb_33_7 bitb_33_7 bitb_33_8 R_bl
Cb_33_7 bit_33_7 gnd C_bl
Cbb_33_7 bitb_33_7 gnd C_bl
Rb_33_8 bit_33_8 bit_33_9 R_bl
Rbb_33_8 bitb_33_8 bitb_33_9 R_bl
Cb_33_8 bit_33_8 gnd C_bl
Cbb_33_8 bitb_33_8 gnd C_bl
Rb_33_9 bit_33_9 bit_33_10 R_bl
Rbb_33_9 bitb_33_9 bitb_33_10 R_bl
Cb_33_9 bit_33_9 gnd C_bl
Cbb_33_9 bitb_33_9 gnd C_bl
Rb_33_10 bit_33_10 bit_33_11 R_bl
Rbb_33_10 bitb_33_10 bitb_33_11 R_bl
Cb_33_10 bit_33_10 gnd C_bl
Cbb_33_10 bitb_33_10 gnd C_bl
Rb_33_11 bit_33_11 bit_33_12 R_bl
Rbb_33_11 bitb_33_11 bitb_33_12 R_bl
Cb_33_11 bit_33_11 gnd C_bl
Cbb_33_11 bitb_33_11 gnd C_bl
Rb_33_12 bit_33_12 bit_33_13 R_bl
Rbb_33_12 bitb_33_12 bitb_33_13 R_bl
Cb_33_12 bit_33_12 gnd C_bl
Cbb_33_12 bitb_33_12 gnd C_bl
Rb_33_13 bit_33_13 bit_33_14 R_bl
Rbb_33_13 bitb_33_13 bitb_33_14 R_bl
Cb_33_13 bit_33_13 gnd C_bl
Cbb_33_13 bitb_33_13 gnd C_bl
Rb_33_14 bit_33_14 bit_33_15 R_bl
Rbb_33_14 bitb_33_14 bitb_33_15 R_bl
Cb_33_14 bit_33_14 gnd C_bl
Cbb_33_14 bitb_33_14 gnd C_bl
Rb_33_15 bit_33_15 bit_33_16 R_bl
Rbb_33_15 bitb_33_15 bitb_33_16 R_bl
Cb_33_15 bit_33_15 gnd C_bl
Cbb_33_15 bitb_33_15 gnd C_bl
Rb_33_16 bit_33_16 bit_33_17 R_bl
Rbb_33_16 bitb_33_16 bitb_33_17 R_bl
Cb_33_16 bit_33_16 gnd C_bl
Cbb_33_16 bitb_33_16 gnd C_bl
Rb_33_17 bit_33_17 bit_33_18 R_bl
Rbb_33_17 bitb_33_17 bitb_33_18 R_bl
Cb_33_17 bit_33_17 gnd C_bl
Cbb_33_17 bitb_33_17 gnd C_bl
Rb_33_18 bit_33_18 bit_33_19 R_bl
Rbb_33_18 bitb_33_18 bitb_33_19 R_bl
Cb_33_18 bit_33_18 gnd C_bl
Cbb_33_18 bitb_33_18 gnd C_bl
Rb_33_19 bit_33_19 bit_33_20 R_bl
Rbb_33_19 bitb_33_19 bitb_33_20 R_bl
Cb_33_19 bit_33_19 gnd C_bl
Cbb_33_19 bitb_33_19 gnd C_bl
Rb_33_20 bit_33_20 bit_33_21 R_bl
Rbb_33_20 bitb_33_20 bitb_33_21 R_bl
Cb_33_20 bit_33_20 gnd C_bl
Cbb_33_20 bitb_33_20 gnd C_bl
Rb_33_21 bit_33_21 bit_33_22 R_bl
Rbb_33_21 bitb_33_21 bitb_33_22 R_bl
Cb_33_21 bit_33_21 gnd C_bl
Cbb_33_21 bitb_33_21 gnd C_bl
Rb_33_22 bit_33_22 bit_33_23 R_bl
Rbb_33_22 bitb_33_22 bitb_33_23 R_bl
Cb_33_22 bit_33_22 gnd C_bl
Cbb_33_22 bitb_33_22 gnd C_bl
Rb_33_23 bit_33_23 bit_33_24 R_bl
Rbb_33_23 bitb_33_23 bitb_33_24 R_bl
Cb_33_23 bit_33_23 gnd C_bl
Cbb_33_23 bitb_33_23 gnd C_bl
Rb_33_24 bit_33_24 bit_33_25 R_bl
Rbb_33_24 bitb_33_24 bitb_33_25 R_bl
Cb_33_24 bit_33_24 gnd C_bl
Cbb_33_24 bitb_33_24 gnd C_bl
Rb_33_25 bit_33_25 bit_33_26 R_bl
Rbb_33_25 bitb_33_25 bitb_33_26 R_bl
Cb_33_25 bit_33_25 gnd C_bl
Cbb_33_25 bitb_33_25 gnd C_bl
Rb_33_26 bit_33_26 bit_33_27 R_bl
Rbb_33_26 bitb_33_26 bitb_33_27 R_bl
Cb_33_26 bit_33_26 gnd C_bl
Cbb_33_26 bitb_33_26 gnd C_bl
Rb_33_27 bit_33_27 bit_33_28 R_bl
Rbb_33_27 bitb_33_27 bitb_33_28 R_bl
Cb_33_27 bit_33_27 gnd C_bl
Cbb_33_27 bitb_33_27 gnd C_bl
Rb_33_28 bit_33_28 bit_33_29 R_bl
Rbb_33_28 bitb_33_28 bitb_33_29 R_bl
Cb_33_28 bit_33_28 gnd C_bl
Cbb_33_28 bitb_33_28 gnd C_bl
Rb_33_29 bit_33_29 bit_33_30 R_bl
Rbb_33_29 bitb_33_29 bitb_33_30 R_bl
Cb_33_29 bit_33_29 gnd C_bl
Cbb_33_29 bitb_33_29 gnd C_bl
Rb_33_30 bit_33_30 bit_33_31 R_bl
Rbb_33_30 bitb_33_30 bitb_33_31 R_bl
Cb_33_30 bit_33_30 gnd C_bl
Cbb_33_30 bitb_33_30 gnd C_bl
Rb_33_31 bit_33_31 bit_33_32 R_bl
Rbb_33_31 bitb_33_31 bitb_33_32 R_bl
Cb_33_31 bit_33_31 gnd C_bl
Cbb_33_31 bitb_33_31 gnd C_bl
Rb_33_32 bit_33_32 bit_33_33 R_bl
Rbb_33_32 bitb_33_32 bitb_33_33 R_bl
Cb_33_32 bit_33_32 gnd C_bl
Cbb_33_32 bitb_33_32 gnd C_bl
Rb_33_33 bit_33_33 bit_33_34 R_bl
Rbb_33_33 bitb_33_33 bitb_33_34 R_bl
Cb_33_33 bit_33_33 gnd C_bl
Cbb_33_33 bitb_33_33 gnd C_bl
Rb_33_34 bit_33_34 bit_33_35 R_bl
Rbb_33_34 bitb_33_34 bitb_33_35 R_bl
Cb_33_34 bit_33_34 gnd C_bl
Cbb_33_34 bitb_33_34 gnd C_bl
Rb_33_35 bit_33_35 bit_33_36 R_bl
Rbb_33_35 bitb_33_35 bitb_33_36 R_bl
Cb_33_35 bit_33_35 gnd C_bl
Cbb_33_35 bitb_33_35 gnd C_bl
Rb_33_36 bit_33_36 bit_33_37 R_bl
Rbb_33_36 bitb_33_36 bitb_33_37 R_bl
Cb_33_36 bit_33_36 gnd C_bl
Cbb_33_36 bitb_33_36 gnd C_bl
Rb_33_37 bit_33_37 bit_33_38 R_bl
Rbb_33_37 bitb_33_37 bitb_33_38 R_bl
Cb_33_37 bit_33_37 gnd C_bl
Cbb_33_37 bitb_33_37 gnd C_bl
Rb_33_38 bit_33_38 bit_33_39 R_bl
Rbb_33_38 bitb_33_38 bitb_33_39 R_bl
Cb_33_38 bit_33_38 gnd C_bl
Cbb_33_38 bitb_33_38 gnd C_bl
Rb_33_39 bit_33_39 bit_33_40 R_bl
Rbb_33_39 bitb_33_39 bitb_33_40 R_bl
Cb_33_39 bit_33_39 gnd C_bl
Cbb_33_39 bitb_33_39 gnd C_bl
Rb_33_40 bit_33_40 bit_33_41 R_bl
Rbb_33_40 bitb_33_40 bitb_33_41 R_bl
Cb_33_40 bit_33_40 gnd C_bl
Cbb_33_40 bitb_33_40 gnd C_bl
Rb_33_41 bit_33_41 bit_33_42 R_bl
Rbb_33_41 bitb_33_41 bitb_33_42 R_bl
Cb_33_41 bit_33_41 gnd C_bl
Cbb_33_41 bitb_33_41 gnd C_bl
Rb_33_42 bit_33_42 bit_33_43 R_bl
Rbb_33_42 bitb_33_42 bitb_33_43 R_bl
Cb_33_42 bit_33_42 gnd C_bl
Cbb_33_42 bitb_33_42 gnd C_bl
Rb_33_43 bit_33_43 bit_33_44 R_bl
Rbb_33_43 bitb_33_43 bitb_33_44 R_bl
Cb_33_43 bit_33_43 gnd C_bl
Cbb_33_43 bitb_33_43 gnd C_bl
Rb_33_44 bit_33_44 bit_33_45 R_bl
Rbb_33_44 bitb_33_44 bitb_33_45 R_bl
Cb_33_44 bit_33_44 gnd C_bl
Cbb_33_44 bitb_33_44 gnd C_bl
Rb_33_45 bit_33_45 bit_33_46 R_bl
Rbb_33_45 bitb_33_45 bitb_33_46 R_bl
Cb_33_45 bit_33_45 gnd C_bl
Cbb_33_45 bitb_33_45 gnd C_bl
Rb_33_46 bit_33_46 bit_33_47 R_bl
Rbb_33_46 bitb_33_46 bitb_33_47 R_bl
Cb_33_46 bit_33_46 gnd C_bl
Cbb_33_46 bitb_33_46 gnd C_bl
Rb_33_47 bit_33_47 bit_33_48 R_bl
Rbb_33_47 bitb_33_47 bitb_33_48 R_bl
Cb_33_47 bit_33_47 gnd C_bl
Cbb_33_47 bitb_33_47 gnd C_bl
Rb_33_48 bit_33_48 bit_33_49 R_bl
Rbb_33_48 bitb_33_48 bitb_33_49 R_bl
Cb_33_48 bit_33_48 gnd C_bl
Cbb_33_48 bitb_33_48 gnd C_bl
Rb_33_49 bit_33_49 bit_33_50 R_bl
Rbb_33_49 bitb_33_49 bitb_33_50 R_bl
Cb_33_49 bit_33_49 gnd C_bl
Cbb_33_49 bitb_33_49 gnd C_bl
Rb_33_50 bit_33_50 bit_33_51 R_bl
Rbb_33_50 bitb_33_50 bitb_33_51 R_bl
Cb_33_50 bit_33_50 gnd C_bl
Cbb_33_50 bitb_33_50 gnd C_bl
Rb_33_51 bit_33_51 bit_33_52 R_bl
Rbb_33_51 bitb_33_51 bitb_33_52 R_bl
Cb_33_51 bit_33_51 gnd C_bl
Cbb_33_51 bitb_33_51 gnd C_bl
Rb_33_52 bit_33_52 bit_33_53 R_bl
Rbb_33_52 bitb_33_52 bitb_33_53 R_bl
Cb_33_52 bit_33_52 gnd C_bl
Cbb_33_52 bitb_33_52 gnd C_bl
Rb_33_53 bit_33_53 bit_33_54 R_bl
Rbb_33_53 bitb_33_53 bitb_33_54 R_bl
Cb_33_53 bit_33_53 gnd C_bl
Cbb_33_53 bitb_33_53 gnd C_bl
Rb_33_54 bit_33_54 bit_33_55 R_bl
Rbb_33_54 bitb_33_54 bitb_33_55 R_bl
Cb_33_54 bit_33_54 gnd C_bl
Cbb_33_54 bitb_33_54 gnd C_bl
Rb_33_55 bit_33_55 bit_33_56 R_bl
Rbb_33_55 bitb_33_55 bitb_33_56 R_bl
Cb_33_55 bit_33_55 gnd C_bl
Cbb_33_55 bitb_33_55 gnd C_bl
Rb_33_56 bit_33_56 bit_33_57 R_bl
Rbb_33_56 bitb_33_56 bitb_33_57 R_bl
Cb_33_56 bit_33_56 gnd C_bl
Cbb_33_56 bitb_33_56 gnd C_bl
Rb_33_57 bit_33_57 bit_33_58 R_bl
Rbb_33_57 bitb_33_57 bitb_33_58 R_bl
Cb_33_57 bit_33_57 gnd C_bl
Cbb_33_57 bitb_33_57 gnd C_bl
Rb_33_58 bit_33_58 bit_33_59 R_bl
Rbb_33_58 bitb_33_58 bitb_33_59 R_bl
Cb_33_58 bit_33_58 gnd C_bl
Cbb_33_58 bitb_33_58 gnd C_bl
Rb_33_59 bit_33_59 bit_33_60 R_bl
Rbb_33_59 bitb_33_59 bitb_33_60 R_bl
Cb_33_59 bit_33_59 gnd C_bl
Cbb_33_59 bitb_33_59 gnd C_bl
Rb_33_60 bit_33_60 bit_33_61 R_bl
Rbb_33_60 bitb_33_60 bitb_33_61 R_bl
Cb_33_60 bit_33_60 gnd C_bl
Cbb_33_60 bitb_33_60 gnd C_bl
Rb_33_61 bit_33_61 bit_33_62 R_bl
Rbb_33_61 bitb_33_61 bitb_33_62 R_bl
Cb_33_61 bit_33_61 gnd C_bl
Cbb_33_61 bitb_33_61 gnd C_bl
Rb_33_62 bit_33_62 bit_33_63 R_bl
Rbb_33_62 bitb_33_62 bitb_33_63 R_bl
Cb_33_62 bit_33_62 gnd C_bl
Cbb_33_62 bitb_33_62 gnd C_bl
Rb_33_63 bit_33_63 bit_33_64 R_bl
Rbb_33_63 bitb_33_63 bitb_33_64 R_bl
Cb_33_63 bit_33_63 gnd C_bl
Cbb_33_63 bitb_33_63 gnd C_bl
Rb_33_64 bit_33_64 bit_33_65 R_bl
Rbb_33_64 bitb_33_64 bitb_33_65 R_bl
Cb_33_64 bit_33_64 gnd C_bl
Cbb_33_64 bitb_33_64 gnd C_bl
Rb_33_65 bit_33_65 bit_33_66 R_bl
Rbb_33_65 bitb_33_65 bitb_33_66 R_bl
Cb_33_65 bit_33_65 gnd C_bl
Cbb_33_65 bitb_33_65 gnd C_bl
Rb_33_66 bit_33_66 bit_33_67 R_bl
Rbb_33_66 bitb_33_66 bitb_33_67 R_bl
Cb_33_66 bit_33_66 gnd C_bl
Cbb_33_66 bitb_33_66 gnd C_bl
Rb_33_67 bit_33_67 bit_33_68 R_bl
Rbb_33_67 bitb_33_67 bitb_33_68 R_bl
Cb_33_67 bit_33_67 gnd C_bl
Cbb_33_67 bitb_33_67 gnd C_bl
Rb_33_68 bit_33_68 bit_33_69 R_bl
Rbb_33_68 bitb_33_68 bitb_33_69 R_bl
Cb_33_68 bit_33_68 gnd C_bl
Cbb_33_68 bitb_33_68 gnd C_bl
Rb_33_69 bit_33_69 bit_33_70 R_bl
Rbb_33_69 bitb_33_69 bitb_33_70 R_bl
Cb_33_69 bit_33_69 gnd C_bl
Cbb_33_69 bitb_33_69 gnd C_bl
Rb_33_70 bit_33_70 bit_33_71 R_bl
Rbb_33_70 bitb_33_70 bitb_33_71 R_bl
Cb_33_70 bit_33_70 gnd C_bl
Cbb_33_70 bitb_33_70 gnd C_bl
Rb_33_71 bit_33_71 bit_33_72 R_bl
Rbb_33_71 bitb_33_71 bitb_33_72 R_bl
Cb_33_71 bit_33_71 gnd C_bl
Cbb_33_71 bitb_33_71 gnd C_bl
Rb_33_72 bit_33_72 bit_33_73 R_bl
Rbb_33_72 bitb_33_72 bitb_33_73 R_bl
Cb_33_72 bit_33_72 gnd C_bl
Cbb_33_72 bitb_33_72 gnd C_bl
Rb_33_73 bit_33_73 bit_33_74 R_bl
Rbb_33_73 bitb_33_73 bitb_33_74 R_bl
Cb_33_73 bit_33_73 gnd C_bl
Cbb_33_73 bitb_33_73 gnd C_bl
Rb_33_74 bit_33_74 bit_33_75 R_bl
Rbb_33_74 bitb_33_74 bitb_33_75 R_bl
Cb_33_74 bit_33_74 gnd C_bl
Cbb_33_74 bitb_33_74 gnd C_bl
Rb_33_75 bit_33_75 bit_33_76 R_bl
Rbb_33_75 bitb_33_75 bitb_33_76 R_bl
Cb_33_75 bit_33_75 gnd C_bl
Cbb_33_75 bitb_33_75 gnd C_bl
Rb_33_76 bit_33_76 bit_33_77 R_bl
Rbb_33_76 bitb_33_76 bitb_33_77 R_bl
Cb_33_76 bit_33_76 gnd C_bl
Cbb_33_76 bitb_33_76 gnd C_bl
Rb_33_77 bit_33_77 bit_33_78 R_bl
Rbb_33_77 bitb_33_77 bitb_33_78 R_bl
Cb_33_77 bit_33_77 gnd C_bl
Cbb_33_77 bitb_33_77 gnd C_bl
Rb_33_78 bit_33_78 bit_33_79 R_bl
Rbb_33_78 bitb_33_78 bitb_33_79 R_bl
Cb_33_78 bit_33_78 gnd C_bl
Cbb_33_78 bitb_33_78 gnd C_bl
Rb_33_79 bit_33_79 bit_33_80 R_bl
Rbb_33_79 bitb_33_79 bitb_33_80 R_bl
Cb_33_79 bit_33_79 gnd C_bl
Cbb_33_79 bitb_33_79 gnd C_bl
Rb_33_80 bit_33_80 bit_33_81 R_bl
Rbb_33_80 bitb_33_80 bitb_33_81 R_bl
Cb_33_80 bit_33_80 gnd C_bl
Cbb_33_80 bitb_33_80 gnd C_bl
Rb_33_81 bit_33_81 bit_33_82 R_bl
Rbb_33_81 bitb_33_81 bitb_33_82 R_bl
Cb_33_81 bit_33_81 gnd C_bl
Cbb_33_81 bitb_33_81 gnd C_bl
Rb_33_82 bit_33_82 bit_33_83 R_bl
Rbb_33_82 bitb_33_82 bitb_33_83 R_bl
Cb_33_82 bit_33_82 gnd C_bl
Cbb_33_82 bitb_33_82 gnd C_bl
Rb_33_83 bit_33_83 bit_33_84 R_bl
Rbb_33_83 bitb_33_83 bitb_33_84 R_bl
Cb_33_83 bit_33_83 gnd C_bl
Cbb_33_83 bitb_33_83 gnd C_bl
Rb_33_84 bit_33_84 bit_33_85 R_bl
Rbb_33_84 bitb_33_84 bitb_33_85 R_bl
Cb_33_84 bit_33_84 gnd C_bl
Cbb_33_84 bitb_33_84 gnd C_bl
Rb_33_85 bit_33_85 bit_33_86 R_bl
Rbb_33_85 bitb_33_85 bitb_33_86 R_bl
Cb_33_85 bit_33_85 gnd C_bl
Cbb_33_85 bitb_33_85 gnd C_bl
Rb_33_86 bit_33_86 bit_33_87 R_bl
Rbb_33_86 bitb_33_86 bitb_33_87 R_bl
Cb_33_86 bit_33_86 gnd C_bl
Cbb_33_86 bitb_33_86 gnd C_bl
Rb_33_87 bit_33_87 bit_33_88 R_bl
Rbb_33_87 bitb_33_87 bitb_33_88 R_bl
Cb_33_87 bit_33_87 gnd C_bl
Cbb_33_87 bitb_33_87 gnd C_bl
Rb_33_88 bit_33_88 bit_33_89 R_bl
Rbb_33_88 bitb_33_88 bitb_33_89 R_bl
Cb_33_88 bit_33_88 gnd C_bl
Cbb_33_88 bitb_33_88 gnd C_bl
Rb_33_89 bit_33_89 bit_33_90 R_bl
Rbb_33_89 bitb_33_89 bitb_33_90 R_bl
Cb_33_89 bit_33_89 gnd C_bl
Cbb_33_89 bitb_33_89 gnd C_bl
Rb_33_90 bit_33_90 bit_33_91 R_bl
Rbb_33_90 bitb_33_90 bitb_33_91 R_bl
Cb_33_90 bit_33_90 gnd C_bl
Cbb_33_90 bitb_33_90 gnd C_bl
Rb_33_91 bit_33_91 bit_33_92 R_bl
Rbb_33_91 bitb_33_91 bitb_33_92 R_bl
Cb_33_91 bit_33_91 gnd C_bl
Cbb_33_91 bitb_33_91 gnd C_bl
Rb_33_92 bit_33_92 bit_33_93 R_bl
Rbb_33_92 bitb_33_92 bitb_33_93 R_bl
Cb_33_92 bit_33_92 gnd C_bl
Cbb_33_92 bitb_33_92 gnd C_bl
Rb_33_93 bit_33_93 bit_33_94 R_bl
Rbb_33_93 bitb_33_93 bitb_33_94 R_bl
Cb_33_93 bit_33_93 gnd C_bl
Cbb_33_93 bitb_33_93 gnd C_bl
Rb_33_94 bit_33_94 bit_33_95 R_bl
Rbb_33_94 bitb_33_94 bitb_33_95 R_bl
Cb_33_94 bit_33_94 gnd C_bl
Cbb_33_94 bitb_33_94 gnd C_bl
Rb_33_95 bit_33_95 bit_33_96 R_bl
Rbb_33_95 bitb_33_95 bitb_33_96 R_bl
Cb_33_95 bit_33_95 gnd C_bl
Cbb_33_95 bitb_33_95 gnd C_bl
Rb_33_96 bit_33_96 bit_33_97 R_bl
Rbb_33_96 bitb_33_96 bitb_33_97 R_bl
Cb_33_96 bit_33_96 gnd C_bl
Cbb_33_96 bitb_33_96 gnd C_bl
Rb_33_97 bit_33_97 bit_33_98 R_bl
Rbb_33_97 bitb_33_97 bitb_33_98 R_bl
Cb_33_97 bit_33_97 gnd C_bl
Cbb_33_97 bitb_33_97 gnd C_bl
Rb_33_98 bit_33_98 bit_33_99 R_bl
Rbb_33_98 bitb_33_98 bitb_33_99 R_bl
Cb_33_98 bit_33_98 gnd C_bl
Cbb_33_98 bitb_33_98 gnd C_bl
Rb_33_99 bit_33_99 bit_33_100 R_bl
Rbb_33_99 bitb_33_99 bitb_33_100 R_bl
Cb_33_99 bit_33_99 gnd C_bl
Cbb_33_99 bitb_33_99 gnd C_bl
Rb_34_0 bit_34_0 bit_34_1 R_bl
Rbb_34_0 bitb_34_0 bitb_34_1 R_bl
Cb_34_0 bit_34_0 gnd C_bl
Cbb_34_0 bitb_34_0 gnd C_bl
Rb_34_1 bit_34_1 bit_34_2 R_bl
Rbb_34_1 bitb_34_1 bitb_34_2 R_bl
Cb_34_1 bit_34_1 gnd C_bl
Cbb_34_1 bitb_34_1 gnd C_bl
Rb_34_2 bit_34_2 bit_34_3 R_bl
Rbb_34_2 bitb_34_2 bitb_34_3 R_bl
Cb_34_2 bit_34_2 gnd C_bl
Cbb_34_2 bitb_34_2 gnd C_bl
Rb_34_3 bit_34_3 bit_34_4 R_bl
Rbb_34_3 bitb_34_3 bitb_34_4 R_bl
Cb_34_3 bit_34_3 gnd C_bl
Cbb_34_3 bitb_34_3 gnd C_bl
Rb_34_4 bit_34_4 bit_34_5 R_bl
Rbb_34_4 bitb_34_4 bitb_34_5 R_bl
Cb_34_4 bit_34_4 gnd C_bl
Cbb_34_4 bitb_34_4 gnd C_bl
Rb_34_5 bit_34_5 bit_34_6 R_bl
Rbb_34_5 bitb_34_5 bitb_34_6 R_bl
Cb_34_5 bit_34_5 gnd C_bl
Cbb_34_5 bitb_34_5 gnd C_bl
Rb_34_6 bit_34_6 bit_34_7 R_bl
Rbb_34_6 bitb_34_6 bitb_34_7 R_bl
Cb_34_6 bit_34_6 gnd C_bl
Cbb_34_6 bitb_34_6 gnd C_bl
Rb_34_7 bit_34_7 bit_34_8 R_bl
Rbb_34_7 bitb_34_7 bitb_34_8 R_bl
Cb_34_7 bit_34_7 gnd C_bl
Cbb_34_7 bitb_34_7 gnd C_bl
Rb_34_8 bit_34_8 bit_34_9 R_bl
Rbb_34_8 bitb_34_8 bitb_34_9 R_bl
Cb_34_8 bit_34_8 gnd C_bl
Cbb_34_8 bitb_34_8 gnd C_bl
Rb_34_9 bit_34_9 bit_34_10 R_bl
Rbb_34_9 bitb_34_9 bitb_34_10 R_bl
Cb_34_9 bit_34_9 gnd C_bl
Cbb_34_9 bitb_34_9 gnd C_bl
Rb_34_10 bit_34_10 bit_34_11 R_bl
Rbb_34_10 bitb_34_10 bitb_34_11 R_bl
Cb_34_10 bit_34_10 gnd C_bl
Cbb_34_10 bitb_34_10 gnd C_bl
Rb_34_11 bit_34_11 bit_34_12 R_bl
Rbb_34_11 bitb_34_11 bitb_34_12 R_bl
Cb_34_11 bit_34_11 gnd C_bl
Cbb_34_11 bitb_34_11 gnd C_bl
Rb_34_12 bit_34_12 bit_34_13 R_bl
Rbb_34_12 bitb_34_12 bitb_34_13 R_bl
Cb_34_12 bit_34_12 gnd C_bl
Cbb_34_12 bitb_34_12 gnd C_bl
Rb_34_13 bit_34_13 bit_34_14 R_bl
Rbb_34_13 bitb_34_13 bitb_34_14 R_bl
Cb_34_13 bit_34_13 gnd C_bl
Cbb_34_13 bitb_34_13 gnd C_bl
Rb_34_14 bit_34_14 bit_34_15 R_bl
Rbb_34_14 bitb_34_14 bitb_34_15 R_bl
Cb_34_14 bit_34_14 gnd C_bl
Cbb_34_14 bitb_34_14 gnd C_bl
Rb_34_15 bit_34_15 bit_34_16 R_bl
Rbb_34_15 bitb_34_15 bitb_34_16 R_bl
Cb_34_15 bit_34_15 gnd C_bl
Cbb_34_15 bitb_34_15 gnd C_bl
Rb_34_16 bit_34_16 bit_34_17 R_bl
Rbb_34_16 bitb_34_16 bitb_34_17 R_bl
Cb_34_16 bit_34_16 gnd C_bl
Cbb_34_16 bitb_34_16 gnd C_bl
Rb_34_17 bit_34_17 bit_34_18 R_bl
Rbb_34_17 bitb_34_17 bitb_34_18 R_bl
Cb_34_17 bit_34_17 gnd C_bl
Cbb_34_17 bitb_34_17 gnd C_bl
Rb_34_18 bit_34_18 bit_34_19 R_bl
Rbb_34_18 bitb_34_18 bitb_34_19 R_bl
Cb_34_18 bit_34_18 gnd C_bl
Cbb_34_18 bitb_34_18 gnd C_bl
Rb_34_19 bit_34_19 bit_34_20 R_bl
Rbb_34_19 bitb_34_19 bitb_34_20 R_bl
Cb_34_19 bit_34_19 gnd C_bl
Cbb_34_19 bitb_34_19 gnd C_bl
Rb_34_20 bit_34_20 bit_34_21 R_bl
Rbb_34_20 bitb_34_20 bitb_34_21 R_bl
Cb_34_20 bit_34_20 gnd C_bl
Cbb_34_20 bitb_34_20 gnd C_bl
Rb_34_21 bit_34_21 bit_34_22 R_bl
Rbb_34_21 bitb_34_21 bitb_34_22 R_bl
Cb_34_21 bit_34_21 gnd C_bl
Cbb_34_21 bitb_34_21 gnd C_bl
Rb_34_22 bit_34_22 bit_34_23 R_bl
Rbb_34_22 bitb_34_22 bitb_34_23 R_bl
Cb_34_22 bit_34_22 gnd C_bl
Cbb_34_22 bitb_34_22 gnd C_bl
Rb_34_23 bit_34_23 bit_34_24 R_bl
Rbb_34_23 bitb_34_23 bitb_34_24 R_bl
Cb_34_23 bit_34_23 gnd C_bl
Cbb_34_23 bitb_34_23 gnd C_bl
Rb_34_24 bit_34_24 bit_34_25 R_bl
Rbb_34_24 bitb_34_24 bitb_34_25 R_bl
Cb_34_24 bit_34_24 gnd C_bl
Cbb_34_24 bitb_34_24 gnd C_bl
Rb_34_25 bit_34_25 bit_34_26 R_bl
Rbb_34_25 bitb_34_25 bitb_34_26 R_bl
Cb_34_25 bit_34_25 gnd C_bl
Cbb_34_25 bitb_34_25 gnd C_bl
Rb_34_26 bit_34_26 bit_34_27 R_bl
Rbb_34_26 bitb_34_26 bitb_34_27 R_bl
Cb_34_26 bit_34_26 gnd C_bl
Cbb_34_26 bitb_34_26 gnd C_bl
Rb_34_27 bit_34_27 bit_34_28 R_bl
Rbb_34_27 bitb_34_27 bitb_34_28 R_bl
Cb_34_27 bit_34_27 gnd C_bl
Cbb_34_27 bitb_34_27 gnd C_bl
Rb_34_28 bit_34_28 bit_34_29 R_bl
Rbb_34_28 bitb_34_28 bitb_34_29 R_bl
Cb_34_28 bit_34_28 gnd C_bl
Cbb_34_28 bitb_34_28 gnd C_bl
Rb_34_29 bit_34_29 bit_34_30 R_bl
Rbb_34_29 bitb_34_29 bitb_34_30 R_bl
Cb_34_29 bit_34_29 gnd C_bl
Cbb_34_29 bitb_34_29 gnd C_bl
Rb_34_30 bit_34_30 bit_34_31 R_bl
Rbb_34_30 bitb_34_30 bitb_34_31 R_bl
Cb_34_30 bit_34_30 gnd C_bl
Cbb_34_30 bitb_34_30 gnd C_bl
Rb_34_31 bit_34_31 bit_34_32 R_bl
Rbb_34_31 bitb_34_31 bitb_34_32 R_bl
Cb_34_31 bit_34_31 gnd C_bl
Cbb_34_31 bitb_34_31 gnd C_bl
Rb_34_32 bit_34_32 bit_34_33 R_bl
Rbb_34_32 bitb_34_32 bitb_34_33 R_bl
Cb_34_32 bit_34_32 gnd C_bl
Cbb_34_32 bitb_34_32 gnd C_bl
Rb_34_33 bit_34_33 bit_34_34 R_bl
Rbb_34_33 bitb_34_33 bitb_34_34 R_bl
Cb_34_33 bit_34_33 gnd C_bl
Cbb_34_33 bitb_34_33 gnd C_bl
Rb_34_34 bit_34_34 bit_34_35 R_bl
Rbb_34_34 bitb_34_34 bitb_34_35 R_bl
Cb_34_34 bit_34_34 gnd C_bl
Cbb_34_34 bitb_34_34 gnd C_bl
Rb_34_35 bit_34_35 bit_34_36 R_bl
Rbb_34_35 bitb_34_35 bitb_34_36 R_bl
Cb_34_35 bit_34_35 gnd C_bl
Cbb_34_35 bitb_34_35 gnd C_bl
Rb_34_36 bit_34_36 bit_34_37 R_bl
Rbb_34_36 bitb_34_36 bitb_34_37 R_bl
Cb_34_36 bit_34_36 gnd C_bl
Cbb_34_36 bitb_34_36 gnd C_bl
Rb_34_37 bit_34_37 bit_34_38 R_bl
Rbb_34_37 bitb_34_37 bitb_34_38 R_bl
Cb_34_37 bit_34_37 gnd C_bl
Cbb_34_37 bitb_34_37 gnd C_bl
Rb_34_38 bit_34_38 bit_34_39 R_bl
Rbb_34_38 bitb_34_38 bitb_34_39 R_bl
Cb_34_38 bit_34_38 gnd C_bl
Cbb_34_38 bitb_34_38 gnd C_bl
Rb_34_39 bit_34_39 bit_34_40 R_bl
Rbb_34_39 bitb_34_39 bitb_34_40 R_bl
Cb_34_39 bit_34_39 gnd C_bl
Cbb_34_39 bitb_34_39 gnd C_bl
Rb_34_40 bit_34_40 bit_34_41 R_bl
Rbb_34_40 bitb_34_40 bitb_34_41 R_bl
Cb_34_40 bit_34_40 gnd C_bl
Cbb_34_40 bitb_34_40 gnd C_bl
Rb_34_41 bit_34_41 bit_34_42 R_bl
Rbb_34_41 bitb_34_41 bitb_34_42 R_bl
Cb_34_41 bit_34_41 gnd C_bl
Cbb_34_41 bitb_34_41 gnd C_bl
Rb_34_42 bit_34_42 bit_34_43 R_bl
Rbb_34_42 bitb_34_42 bitb_34_43 R_bl
Cb_34_42 bit_34_42 gnd C_bl
Cbb_34_42 bitb_34_42 gnd C_bl
Rb_34_43 bit_34_43 bit_34_44 R_bl
Rbb_34_43 bitb_34_43 bitb_34_44 R_bl
Cb_34_43 bit_34_43 gnd C_bl
Cbb_34_43 bitb_34_43 gnd C_bl
Rb_34_44 bit_34_44 bit_34_45 R_bl
Rbb_34_44 bitb_34_44 bitb_34_45 R_bl
Cb_34_44 bit_34_44 gnd C_bl
Cbb_34_44 bitb_34_44 gnd C_bl
Rb_34_45 bit_34_45 bit_34_46 R_bl
Rbb_34_45 bitb_34_45 bitb_34_46 R_bl
Cb_34_45 bit_34_45 gnd C_bl
Cbb_34_45 bitb_34_45 gnd C_bl
Rb_34_46 bit_34_46 bit_34_47 R_bl
Rbb_34_46 bitb_34_46 bitb_34_47 R_bl
Cb_34_46 bit_34_46 gnd C_bl
Cbb_34_46 bitb_34_46 gnd C_bl
Rb_34_47 bit_34_47 bit_34_48 R_bl
Rbb_34_47 bitb_34_47 bitb_34_48 R_bl
Cb_34_47 bit_34_47 gnd C_bl
Cbb_34_47 bitb_34_47 gnd C_bl
Rb_34_48 bit_34_48 bit_34_49 R_bl
Rbb_34_48 bitb_34_48 bitb_34_49 R_bl
Cb_34_48 bit_34_48 gnd C_bl
Cbb_34_48 bitb_34_48 gnd C_bl
Rb_34_49 bit_34_49 bit_34_50 R_bl
Rbb_34_49 bitb_34_49 bitb_34_50 R_bl
Cb_34_49 bit_34_49 gnd C_bl
Cbb_34_49 bitb_34_49 gnd C_bl
Rb_34_50 bit_34_50 bit_34_51 R_bl
Rbb_34_50 bitb_34_50 bitb_34_51 R_bl
Cb_34_50 bit_34_50 gnd C_bl
Cbb_34_50 bitb_34_50 gnd C_bl
Rb_34_51 bit_34_51 bit_34_52 R_bl
Rbb_34_51 bitb_34_51 bitb_34_52 R_bl
Cb_34_51 bit_34_51 gnd C_bl
Cbb_34_51 bitb_34_51 gnd C_bl
Rb_34_52 bit_34_52 bit_34_53 R_bl
Rbb_34_52 bitb_34_52 bitb_34_53 R_bl
Cb_34_52 bit_34_52 gnd C_bl
Cbb_34_52 bitb_34_52 gnd C_bl
Rb_34_53 bit_34_53 bit_34_54 R_bl
Rbb_34_53 bitb_34_53 bitb_34_54 R_bl
Cb_34_53 bit_34_53 gnd C_bl
Cbb_34_53 bitb_34_53 gnd C_bl
Rb_34_54 bit_34_54 bit_34_55 R_bl
Rbb_34_54 bitb_34_54 bitb_34_55 R_bl
Cb_34_54 bit_34_54 gnd C_bl
Cbb_34_54 bitb_34_54 gnd C_bl
Rb_34_55 bit_34_55 bit_34_56 R_bl
Rbb_34_55 bitb_34_55 bitb_34_56 R_bl
Cb_34_55 bit_34_55 gnd C_bl
Cbb_34_55 bitb_34_55 gnd C_bl
Rb_34_56 bit_34_56 bit_34_57 R_bl
Rbb_34_56 bitb_34_56 bitb_34_57 R_bl
Cb_34_56 bit_34_56 gnd C_bl
Cbb_34_56 bitb_34_56 gnd C_bl
Rb_34_57 bit_34_57 bit_34_58 R_bl
Rbb_34_57 bitb_34_57 bitb_34_58 R_bl
Cb_34_57 bit_34_57 gnd C_bl
Cbb_34_57 bitb_34_57 gnd C_bl
Rb_34_58 bit_34_58 bit_34_59 R_bl
Rbb_34_58 bitb_34_58 bitb_34_59 R_bl
Cb_34_58 bit_34_58 gnd C_bl
Cbb_34_58 bitb_34_58 gnd C_bl
Rb_34_59 bit_34_59 bit_34_60 R_bl
Rbb_34_59 bitb_34_59 bitb_34_60 R_bl
Cb_34_59 bit_34_59 gnd C_bl
Cbb_34_59 bitb_34_59 gnd C_bl
Rb_34_60 bit_34_60 bit_34_61 R_bl
Rbb_34_60 bitb_34_60 bitb_34_61 R_bl
Cb_34_60 bit_34_60 gnd C_bl
Cbb_34_60 bitb_34_60 gnd C_bl
Rb_34_61 bit_34_61 bit_34_62 R_bl
Rbb_34_61 bitb_34_61 bitb_34_62 R_bl
Cb_34_61 bit_34_61 gnd C_bl
Cbb_34_61 bitb_34_61 gnd C_bl
Rb_34_62 bit_34_62 bit_34_63 R_bl
Rbb_34_62 bitb_34_62 bitb_34_63 R_bl
Cb_34_62 bit_34_62 gnd C_bl
Cbb_34_62 bitb_34_62 gnd C_bl
Rb_34_63 bit_34_63 bit_34_64 R_bl
Rbb_34_63 bitb_34_63 bitb_34_64 R_bl
Cb_34_63 bit_34_63 gnd C_bl
Cbb_34_63 bitb_34_63 gnd C_bl
Rb_34_64 bit_34_64 bit_34_65 R_bl
Rbb_34_64 bitb_34_64 bitb_34_65 R_bl
Cb_34_64 bit_34_64 gnd C_bl
Cbb_34_64 bitb_34_64 gnd C_bl
Rb_34_65 bit_34_65 bit_34_66 R_bl
Rbb_34_65 bitb_34_65 bitb_34_66 R_bl
Cb_34_65 bit_34_65 gnd C_bl
Cbb_34_65 bitb_34_65 gnd C_bl
Rb_34_66 bit_34_66 bit_34_67 R_bl
Rbb_34_66 bitb_34_66 bitb_34_67 R_bl
Cb_34_66 bit_34_66 gnd C_bl
Cbb_34_66 bitb_34_66 gnd C_bl
Rb_34_67 bit_34_67 bit_34_68 R_bl
Rbb_34_67 bitb_34_67 bitb_34_68 R_bl
Cb_34_67 bit_34_67 gnd C_bl
Cbb_34_67 bitb_34_67 gnd C_bl
Rb_34_68 bit_34_68 bit_34_69 R_bl
Rbb_34_68 bitb_34_68 bitb_34_69 R_bl
Cb_34_68 bit_34_68 gnd C_bl
Cbb_34_68 bitb_34_68 gnd C_bl
Rb_34_69 bit_34_69 bit_34_70 R_bl
Rbb_34_69 bitb_34_69 bitb_34_70 R_bl
Cb_34_69 bit_34_69 gnd C_bl
Cbb_34_69 bitb_34_69 gnd C_bl
Rb_34_70 bit_34_70 bit_34_71 R_bl
Rbb_34_70 bitb_34_70 bitb_34_71 R_bl
Cb_34_70 bit_34_70 gnd C_bl
Cbb_34_70 bitb_34_70 gnd C_bl
Rb_34_71 bit_34_71 bit_34_72 R_bl
Rbb_34_71 bitb_34_71 bitb_34_72 R_bl
Cb_34_71 bit_34_71 gnd C_bl
Cbb_34_71 bitb_34_71 gnd C_bl
Rb_34_72 bit_34_72 bit_34_73 R_bl
Rbb_34_72 bitb_34_72 bitb_34_73 R_bl
Cb_34_72 bit_34_72 gnd C_bl
Cbb_34_72 bitb_34_72 gnd C_bl
Rb_34_73 bit_34_73 bit_34_74 R_bl
Rbb_34_73 bitb_34_73 bitb_34_74 R_bl
Cb_34_73 bit_34_73 gnd C_bl
Cbb_34_73 bitb_34_73 gnd C_bl
Rb_34_74 bit_34_74 bit_34_75 R_bl
Rbb_34_74 bitb_34_74 bitb_34_75 R_bl
Cb_34_74 bit_34_74 gnd C_bl
Cbb_34_74 bitb_34_74 gnd C_bl
Rb_34_75 bit_34_75 bit_34_76 R_bl
Rbb_34_75 bitb_34_75 bitb_34_76 R_bl
Cb_34_75 bit_34_75 gnd C_bl
Cbb_34_75 bitb_34_75 gnd C_bl
Rb_34_76 bit_34_76 bit_34_77 R_bl
Rbb_34_76 bitb_34_76 bitb_34_77 R_bl
Cb_34_76 bit_34_76 gnd C_bl
Cbb_34_76 bitb_34_76 gnd C_bl
Rb_34_77 bit_34_77 bit_34_78 R_bl
Rbb_34_77 bitb_34_77 bitb_34_78 R_bl
Cb_34_77 bit_34_77 gnd C_bl
Cbb_34_77 bitb_34_77 gnd C_bl
Rb_34_78 bit_34_78 bit_34_79 R_bl
Rbb_34_78 bitb_34_78 bitb_34_79 R_bl
Cb_34_78 bit_34_78 gnd C_bl
Cbb_34_78 bitb_34_78 gnd C_bl
Rb_34_79 bit_34_79 bit_34_80 R_bl
Rbb_34_79 bitb_34_79 bitb_34_80 R_bl
Cb_34_79 bit_34_79 gnd C_bl
Cbb_34_79 bitb_34_79 gnd C_bl
Rb_34_80 bit_34_80 bit_34_81 R_bl
Rbb_34_80 bitb_34_80 bitb_34_81 R_bl
Cb_34_80 bit_34_80 gnd C_bl
Cbb_34_80 bitb_34_80 gnd C_bl
Rb_34_81 bit_34_81 bit_34_82 R_bl
Rbb_34_81 bitb_34_81 bitb_34_82 R_bl
Cb_34_81 bit_34_81 gnd C_bl
Cbb_34_81 bitb_34_81 gnd C_bl
Rb_34_82 bit_34_82 bit_34_83 R_bl
Rbb_34_82 bitb_34_82 bitb_34_83 R_bl
Cb_34_82 bit_34_82 gnd C_bl
Cbb_34_82 bitb_34_82 gnd C_bl
Rb_34_83 bit_34_83 bit_34_84 R_bl
Rbb_34_83 bitb_34_83 bitb_34_84 R_bl
Cb_34_83 bit_34_83 gnd C_bl
Cbb_34_83 bitb_34_83 gnd C_bl
Rb_34_84 bit_34_84 bit_34_85 R_bl
Rbb_34_84 bitb_34_84 bitb_34_85 R_bl
Cb_34_84 bit_34_84 gnd C_bl
Cbb_34_84 bitb_34_84 gnd C_bl
Rb_34_85 bit_34_85 bit_34_86 R_bl
Rbb_34_85 bitb_34_85 bitb_34_86 R_bl
Cb_34_85 bit_34_85 gnd C_bl
Cbb_34_85 bitb_34_85 gnd C_bl
Rb_34_86 bit_34_86 bit_34_87 R_bl
Rbb_34_86 bitb_34_86 bitb_34_87 R_bl
Cb_34_86 bit_34_86 gnd C_bl
Cbb_34_86 bitb_34_86 gnd C_bl
Rb_34_87 bit_34_87 bit_34_88 R_bl
Rbb_34_87 bitb_34_87 bitb_34_88 R_bl
Cb_34_87 bit_34_87 gnd C_bl
Cbb_34_87 bitb_34_87 gnd C_bl
Rb_34_88 bit_34_88 bit_34_89 R_bl
Rbb_34_88 bitb_34_88 bitb_34_89 R_bl
Cb_34_88 bit_34_88 gnd C_bl
Cbb_34_88 bitb_34_88 gnd C_bl
Rb_34_89 bit_34_89 bit_34_90 R_bl
Rbb_34_89 bitb_34_89 bitb_34_90 R_bl
Cb_34_89 bit_34_89 gnd C_bl
Cbb_34_89 bitb_34_89 gnd C_bl
Rb_34_90 bit_34_90 bit_34_91 R_bl
Rbb_34_90 bitb_34_90 bitb_34_91 R_bl
Cb_34_90 bit_34_90 gnd C_bl
Cbb_34_90 bitb_34_90 gnd C_bl
Rb_34_91 bit_34_91 bit_34_92 R_bl
Rbb_34_91 bitb_34_91 bitb_34_92 R_bl
Cb_34_91 bit_34_91 gnd C_bl
Cbb_34_91 bitb_34_91 gnd C_bl
Rb_34_92 bit_34_92 bit_34_93 R_bl
Rbb_34_92 bitb_34_92 bitb_34_93 R_bl
Cb_34_92 bit_34_92 gnd C_bl
Cbb_34_92 bitb_34_92 gnd C_bl
Rb_34_93 bit_34_93 bit_34_94 R_bl
Rbb_34_93 bitb_34_93 bitb_34_94 R_bl
Cb_34_93 bit_34_93 gnd C_bl
Cbb_34_93 bitb_34_93 gnd C_bl
Rb_34_94 bit_34_94 bit_34_95 R_bl
Rbb_34_94 bitb_34_94 bitb_34_95 R_bl
Cb_34_94 bit_34_94 gnd C_bl
Cbb_34_94 bitb_34_94 gnd C_bl
Rb_34_95 bit_34_95 bit_34_96 R_bl
Rbb_34_95 bitb_34_95 bitb_34_96 R_bl
Cb_34_95 bit_34_95 gnd C_bl
Cbb_34_95 bitb_34_95 gnd C_bl
Rb_34_96 bit_34_96 bit_34_97 R_bl
Rbb_34_96 bitb_34_96 bitb_34_97 R_bl
Cb_34_96 bit_34_96 gnd C_bl
Cbb_34_96 bitb_34_96 gnd C_bl
Rb_34_97 bit_34_97 bit_34_98 R_bl
Rbb_34_97 bitb_34_97 bitb_34_98 R_bl
Cb_34_97 bit_34_97 gnd C_bl
Cbb_34_97 bitb_34_97 gnd C_bl
Rb_34_98 bit_34_98 bit_34_99 R_bl
Rbb_34_98 bitb_34_98 bitb_34_99 R_bl
Cb_34_98 bit_34_98 gnd C_bl
Cbb_34_98 bitb_34_98 gnd C_bl
Rb_34_99 bit_34_99 bit_34_100 R_bl
Rbb_34_99 bitb_34_99 bitb_34_100 R_bl
Cb_34_99 bit_34_99 gnd C_bl
Cbb_34_99 bitb_34_99 gnd C_bl
Rb_35_0 bit_35_0 bit_35_1 R_bl
Rbb_35_0 bitb_35_0 bitb_35_1 R_bl
Cb_35_0 bit_35_0 gnd C_bl
Cbb_35_0 bitb_35_0 gnd C_bl
Rb_35_1 bit_35_1 bit_35_2 R_bl
Rbb_35_1 bitb_35_1 bitb_35_2 R_bl
Cb_35_1 bit_35_1 gnd C_bl
Cbb_35_1 bitb_35_1 gnd C_bl
Rb_35_2 bit_35_2 bit_35_3 R_bl
Rbb_35_2 bitb_35_2 bitb_35_3 R_bl
Cb_35_2 bit_35_2 gnd C_bl
Cbb_35_2 bitb_35_2 gnd C_bl
Rb_35_3 bit_35_3 bit_35_4 R_bl
Rbb_35_3 bitb_35_3 bitb_35_4 R_bl
Cb_35_3 bit_35_3 gnd C_bl
Cbb_35_3 bitb_35_3 gnd C_bl
Rb_35_4 bit_35_4 bit_35_5 R_bl
Rbb_35_4 bitb_35_4 bitb_35_5 R_bl
Cb_35_4 bit_35_4 gnd C_bl
Cbb_35_4 bitb_35_4 gnd C_bl
Rb_35_5 bit_35_5 bit_35_6 R_bl
Rbb_35_5 bitb_35_5 bitb_35_6 R_bl
Cb_35_5 bit_35_5 gnd C_bl
Cbb_35_5 bitb_35_5 gnd C_bl
Rb_35_6 bit_35_6 bit_35_7 R_bl
Rbb_35_6 bitb_35_6 bitb_35_7 R_bl
Cb_35_6 bit_35_6 gnd C_bl
Cbb_35_6 bitb_35_6 gnd C_bl
Rb_35_7 bit_35_7 bit_35_8 R_bl
Rbb_35_7 bitb_35_7 bitb_35_8 R_bl
Cb_35_7 bit_35_7 gnd C_bl
Cbb_35_7 bitb_35_7 gnd C_bl
Rb_35_8 bit_35_8 bit_35_9 R_bl
Rbb_35_8 bitb_35_8 bitb_35_9 R_bl
Cb_35_8 bit_35_8 gnd C_bl
Cbb_35_8 bitb_35_8 gnd C_bl
Rb_35_9 bit_35_9 bit_35_10 R_bl
Rbb_35_9 bitb_35_9 bitb_35_10 R_bl
Cb_35_9 bit_35_9 gnd C_bl
Cbb_35_9 bitb_35_9 gnd C_bl
Rb_35_10 bit_35_10 bit_35_11 R_bl
Rbb_35_10 bitb_35_10 bitb_35_11 R_bl
Cb_35_10 bit_35_10 gnd C_bl
Cbb_35_10 bitb_35_10 gnd C_bl
Rb_35_11 bit_35_11 bit_35_12 R_bl
Rbb_35_11 bitb_35_11 bitb_35_12 R_bl
Cb_35_11 bit_35_11 gnd C_bl
Cbb_35_11 bitb_35_11 gnd C_bl
Rb_35_12 bit_35_12 bit_35_13 R_bl
Rbb_35_12 bitb_35_12 bitb_35_13 R_bl
Cb_35_12 bit_35_12 gnd C_bl
Cbb_35_12 bitb_35_12 gnd C_bl
Rb_35_13 bit_35_13 bit_35_14 R_bl
Rbb_35_13 bitb_35_13 bitb_35_14 R_bl
Cb_35_13 bit_35_13 gnd C_bl
Cbb_35_13 bitb_35_13 gnd C_bl
Rb_35_14 bit_35_14 bit_35_15 R_bl
Rbb_35_14 bitb_35_14 bitb_35_15 R_bl
Cb_35_14 bit_35_14 gnd C_bl
Cbb_35_14 bitb_35_14 gnd C_bl
Rb_35_15 bit_35_15 bit_35_16 R_bl
Rbb_35_15 bitb_35_15 bitb_35_16 R_bl
Cb_35_15 bit_35_15 gnd C_bl
Cbb_35_15 bitb_35_15 gnd C_bl
Rb_35_16 bit_35_16 bit_35_17 R_bl
Rbb_35_16 bitb_35_16 bitb_35_17 R_bl
Cb_35_16 bit_35_16 gnd C_bl
Cbb_35_16 bitb_35_16 gnd C_bl
Rb_35_17 bit_35_17 bit_35_18 R_bl
Rbb_35_17 bitb_35_17 bitb_35_18 R_bl
Cb_35_17 bit_35_17 gnd C_bl
Cbb_35_17 bitb_35_17 gnd C_bl
Rb_35_18 bit_35_18 bit_35_19 R_bl
Rbb_35_18 bitb_35_18 bitb_35_19 R_bl
Cb_35_18 bit_35_18 gnd C_bl
Cbb_35_18 bitb_35_18 gnd C_bl
Rb_35_19 bit_35_19 bit_35_20 R_bl
Rbb_35_19 bitb_35_19 bitb_35_20 R_bl
Cb_35_19 bit_35_19 gnd C_bl
Cbb_35_19 bitb_35_19 gnd C_bl
Rb_35_20 bit_35_20 bit_35_21 R_bl
Rbb_35_20 bitb_35_20 bitb_35_21 R_bl
Cb_35_20 bit_35_20 gnd C_bl
Cbb_35_20 bitb_35_20 gnd C_bl
Rb_35_21 bit_35_21 bit_35_22 R_bl
Rbb_35_21 bitb_35_21 bitb_35_22 R_bl
Cb_35_21 bit_35_21 gnd C_bl
Cbb_35_21 bitb_35_21 gnd C_bl
Rb_35_22 bit_35_22 bit_35_23 R_bl
Rbb_35_22 bitb_35_22 bitb_35_23 R_bl
Cb_35_22 bit_35_22 gnd C_bl
Cbb_35_22 bitb_35_22 gnd C_bl
Rb_35_23 bit_35_23 bit_35_24 R_bl
Rbb_35_23 bitb_35_23 bitb_35_24 R_bl
Cb_35_23 bit_35_23 gnd C_bl
Cbb_35_23 bitb_35_23 gnd C_bl
Rb_35_24 bit_35_24 bit_35_25 R_bl
Rbb_35_24 bitb_35_24 bitb_35_25 R_bl
Cb_35_24 bit_35_24 gnd C_bl
Cbb_35_24 bitb_35_24 gnd C_bl
Rb_35_25 bit_35_25 bit_35_26 R_bl
Rbb_35_25 bitb_35_25 bitb_35_26 R_bl
Cb_35_25 bit_35_25 gnd C_bl
Cbb_35_25 bitb_35_25 gnd C_bl
Rb_35_26 bit_35_26 bit_35_27 R_bl
Rbb_35_26 bitb_35_26 bitb_35_27 R_bl
Cb_35_26 bit_35_26 gnd C_bl
Cbb_35_26 bitb_35_26 gnd C_bl
Rb_35_27 bit_35_27 bit_35_28 R_bl
Rbb_35_27 bitb_35_27 bitb_35_28 R_bl
Cb_35_27 bit_35_27 gnd C_bl
Cbb_35_27 bitb_35_27 gnd C_bl
Rb_35_28 bit_35_28 bit_35_29 R_bl
Rbb_35_28 bitb_35_28 bitb_35_29 R_bl
Cb_35_28 bit_35_28 gnd C_bl
Cbb_35_28 bitb_35_28 gnd C_bl
Rb_35_29 bit_35_29 bit_35_30 R_bl
Rbb_35_29 bitb_35_29 bitb_35_30 R_bl
Cb_35_29 bit_35_29 gnd C_bl
Cbb_35_29 bitb_35_29 gnd C_bl
Rb_35_30 bit_35_30 bit_35_31 R_bl
Rbb_35_30 bitb_35_30 bitb_35_31 R_bl
Cb_35_30 bit_35_30 gnd C_bl
Cbb_35_30 bitb_35_30 gnd C_bl
Rb_35_31 bit_35_31 bit_35_32 R_bl
Rbb_35_31 bitb_35_31 bitb_35_32 R_bl
Cb_35_31 bit_35_31 gnd C_bl
Cbb_35_31 bitb_35_31 gnd C_bl
Rb_35_32 bit_35_32 bit_35_33 R_bl
Rbb_35_32 bitb_35_32 bitb_35_33 R_bl
Cb_35_32 bit_35_32 gnd C_bl
Cbb_35_32 bitb_35_32 gnd C_bl
Rb_35_33 bit_35_33 bit_35_34 R_bl
Rbb_35_33 bitb_35_33 bitb_35_34 R_bl
Cb_35_33 bit_35_33 gnd C_bl
Cbb_35_33 bitb_35_33 gnd C_bl
Rb_35_34 bit_35_34 bit_35_35 R_bl
Rbb_35_34 bitb_35_34 bitb_35_35 R_bl
Cb_35_34 bit_35_34 gnd C_bl
Cbb_35_34 bitb_35_34 gnd C_bl
Rb_35_35 bit_35_35 bit_35_36 R_bl
Rbb_35_35 bitb_35_35 bitb_35_36 R_bl
Cb_35_35 bit_35_35 gnd C_bl
Cbb_35_35 bitb_35_35 gnd C_bl
Rb_35_36 bit_35_36 bit_35_37 R_bl
Rbb_35_36 bitb_35_36 bitb_35_37 R_bl
Cb_35_36 bit_35_36 gnd C_bl
Cbb_35_36 bitb_35_36 gnd C_bl
Rb_35_37 bit_35_37 bit_35_38 R_bl
Rbb_35_37 bitb_35_37 bitb_35_38 R_bl
Cb_35_37 bit_35_37 gnd C_bl
Cbb_35_37 bitb_35_37 gnd C_bl
Rb_35_38 bit_35_38 bit_35_39 R_bl
Rbb_35_38 bitb_35_38 bitb_35_39 R_bl
Cb_35_38 bit_35_38 gnd C_bl
Cbb_35_38 bitb_35_38 gnd C_bl
Rb_35_39 bit_35_39 bit_35_40 R_bl
Rbb_35_39 bitb_35_39 bitb_35_40 R_bl
Cb_35_39 bit_35_39 gnd C_bl
Cbb_35_39 bitb_35_39 gnd C_bl
Rb_35_40 bit_35_40 bit_35_41 R_bl
Rbb_35_40 bitb_35_40 bitb_35_41 R_bl
Cb_35_40 bit_35_40 gnd C_bl
Cbb_35_40 bitb_35_40 gnd C_bl
Rb_35_41 bit_35_41 bit_35_42 R_bl
Rbb_35_41 bitb_35_41 bitb_35_42 R_bl
Cb_35_41 bit_35_41 gnd C_bl
Cbb_35_41 bitb_35_41 gnd C_bl
Rb_35_42 bit_35_42 bit_35_43 R_bl
Rbb_35_42 bitb_35_42 bitb_35_43 R_bl
Cb_35_42 bit_35_42 gnd C_bl
Cbb_35_42 bitb_35_42 gnd C_bl
Rb_35_43 bit_35_43 bit_35_44 R_bl
Rbb_35_43 bitb_35_43 bitb_35_44 R_bl
Cb_35_43 bit_35_43 gnd C_bl
Cbb_35_43 bitb_35_43 gnd C_bl
Rb_35_44 bit_35_44 bit_35_45 R_bl
Rbb_35_44 bitb_35_44 bitb_35_45 R_bl
Cb_35_44 bit_35_44 gnd C_bl
Cbb_35_44 bitb_35_44 gnd C_bl
Rb_35_45 bit_35_45 bit_35_46 R_bl
Rbb_35_45 bitb_35_45 bitb_35_46 R_bl
Cb_35_45 bit_35_45 gnd C_bl
Cbb_35_45 bitb_35_45 gnd C_bl
Rb_35_46 bit_35_46 bit_35_47 R_bl
Rbb_35_46 bitb_35_46 bitb_35_47 R_bl
Cb_35_46 bit_35_46 gnd C_bl
Cbb_35_46 bitb_35_46 gnd C_bl
Rb_35_47 bit_35_47 bit_35_48 R_bl
Rbb_35_47 bitb_35_47 bitb_35_48 R_bl
Cb_35_47 bit_35_47 gnd C_bl
Cbb_35_47 bitb_35_47 gnd C_bl
Rb_35_48 bit_35_48 bit_35_49 R_bl
Rbb_35_48 bitb_35_48 bitb_35_49 R_bl
Cb_35_48 bit_35_48 gnd C_bl
Cbb_35_48 bitb_35_48 gnd C_bl
Rb_35_49 bit_35_49 bit_35_50 R_bl
Rbb_35_49 bitb_35_49 bitb_35_50 R_bl
Cb_35_49 bit_35_49 gnd C_bl
Cbb_35_49 bitb_35_49 gnd C_bl
Rb_35_50 bit_35_50 bit_35_51 R_bl
Rbb_35_50 bitb_35_50 bitb_35_51 R_bl
Cb_35_50 bit_35_50 gnd C_bl
Cbb_35_50 bitb_35_50 gnd C_bl
Rb_35_51 bit_35_51 bit_35_52 R_bl
Rbb_35_51 bitb_35_51 bitb_35_52 R_bl
Cb_35_51 bit_35_51 gnd C_bl
Cbb_35_51 bitb_35_51 gnd C_bl
Rb_35_52 bit_35_52 bit_35_53 R_bl
Rbb_35_52 bitb_35_52 bitb_35_53 R_bl
Cb_35_52 bit_35_52 gnd C_bl
Cbb_35_52 bitb_35_52 gnd C_bl
Rb_35_53 bit_35_53 bit_35_54 R_bl
Rbb_35_53 bitb_35_53 bitb_35_54 R_bl
Cb_35_53 bit_35_53 gnd C_bl
Cbb_35_53 bitb_35_53 gnd C_bl
Rb_35_54 bit_35_54 bit_35_55 R_bl
Rbb_35_54 bitb_35_54 bitb_35_55 R_bl
Cb_35_54 bit_35_54 gnd C_bl
Cbb_35_54 bitb_35_54 gnd C_bl
Rb_35_55 bit_35_55 bit_35_56 R_bl
Rbb_35_55 bitb_35_55 bitb_35_56 R_bl
Cb_35_55 bit_35_55 gnd C_bl
Cbb_35_55 bitb_35_55 gnd C_bl
Rb_35_56 bit_35_56 bit_35_57 R_bl
Rbb_35_56 bitb_35_56 bitb_35_57 R_bl
Cb_35_56 bit_35_56 gnd C_bl
Cbb_35_56 bitb_35_56 gnd C_bl
Rb_35_57 bit_35_57 bit_35_58 R_bl
Rbb_35_57 bitb_35_57 bitb_35_58 R_bl
Cb_35_57 bit_35_57 gnd C_bl
Cbb_35_57 bitb_35_57 gnd C_bl
Rb_35_58 bit_35_58 bit_35_59 R_bl
Rbb_35_58 bitb_35_58 bitb_35_59 R_bl
Cb_35_58 bit_35_58 gnd C_bl
Cbb_35_58 bitb_35_58 gnd C_bl
Rb_35_59 bit_35_59 bit_35_60 R_bl
Rbb_35_59 bitb_35_59 bitb_35_60 R_bl
Cb_35_59 bit_35_59 gnd C_bl
Cbb_35_59 bitb_35_59 gnd C_bl
Rb_35_60 bit_35_60 bit_35_61 R_bl
Rbb_35_60 bitb_35_60 bitb_35_61 R_bl
Cb_35_60 bit_35_60 gnd C_bl
Cbb_35_60 bitb_35_60 gnd C_bl
Rb_35_61 bit_35_61 bit_35_62 R_bl
Rbb_35_61 bitb_35_61 bitb_35_62 R_bl
Cb_35_61 bit_35_61 gnd C_bl
Cbb_35_61 bitb_35_61 gnd C_bl
Rb_35_62 bit_35_62 bit_35_63 R_bl
Rbb_35_62 bitb_35_62 bitb_35_63 R_bl
Cb_35_62 bit_35_62 gnd C_bl
Cbb_35_62 bitb_35_62 gnd C_bl
Rb_35_63 bit_35_63 bit_35_64 R_bl
Rbb_35_63 bitb_35_63 bitb_35_64 R_bl
Cb_35_63 bit_35_63 gnd C_bl
Cbb_35_63 bitb_35_63 gnd C_bl
Rb_35_64 bit_35_64 bit_35_65 R_bl
Rbb_35_64 bitb_35_64 bitb_35_65 R_bl
Cb_35_64 bit_35_64 gnd C_bl
Cbb_35_64 bitb_35_64 gnd C_bl
Rb_35_65 bit_35_65 bit_35_66 R_bl
Rbb_35_65 bitb_35_65 bitb_35_66 R_bl
Cb_35_65 bit_35_65 gnd C_bl
Cbb_35_65 bitb_35_65 gnd C_bl
Rb_35_66 bit_35_66 bit_35_67 R_bl
Rbb_35_66 bitb_35_66 bitb_35_67 R_bl
Cb_35_66 bit_35_66 gnd C_bl
Cbb_35_66 bitb_35_66 gnd C_bl
Rb_35_67 bit_35_67 bit_35_68 R_bl
Rbb_35_67 bitb_35_67 bitb_35_68 R_bl
Cb_35_67 bit_35_67 gnd C_bl
Cbb_35_67 bitb_35_67 gnd C_bl
Rb_35_68 bit_35_68 bit_35_69 R_bl
Rbb_35_68 bitb_35_68 bitb_35_69 R_bl
Cb_35_68 bit_35_68 gnd C_bl
Cbb_35_68 bitb_35_68 gnd C_bl
Rb_35_69 bit_35_69 bit_35_70 R_bl
Rbb_35_69 bitb_35_69 bitb_35_70 R_bl
Cb_35_69 bit_35_69 gnd C_bl
Cbb_35_69 bitb_35_69 gnd C_bl
Rb_35_70 bit_35_70 bit_35_71 R_bl
Rbb_35_70 bitb_35_70 bitb_35_71 R_bl
Cb_35_70 bit_35_70 gnd C_bl
Cbb_35_70 bitb_35_70 gnd C_bl
Rb_35_71 bit_35_71 bit_35_72 R_bl
Rbb_35_71 bitb_35_71 bitb_35_72 R_bl
Cb_35_71 bit_35_71 gnd C_bl
Cbb_35_71 bitb_35_71 gnd C_bl
Rb_35_72 bit_35_72 bit_35_73 R_bl
Rbb_35_72 bitb_35_72 bitb_35_73 R_bl
Cb_35_72 bit_35_72 gnd C_bl
Cbb_35_72 bitb_35_72 gnd C_bl
Rb_35_73 bit_35_73 bit_35_74 R_bl
Rbb_35_73 bitb_35_73 bitb_35_74 R_bl
Cb_35_73 bit_35_73 gnd C_bl
Cbb_35_73 bitb_35_73 gnd C_bl
Rb_35_74 bit_35_74 bit_35_75 R_bl
Rbb_35_74 bitb_35_74 bitb_35_75 R_bl
Cb_35_74 bit_35_74 gnd C_bl
Cbb_35_74 bitb_35_74 gnd C_bl
Rb_35_75 bit_35_75 bit_35_76 R_bl
Rbb_35_75 bitb_35_75 bitb_35_76 R_bl
Cb_35_75 bit_35_75 gnd C_bl
Cbb_35_75 bitb_35_75 gnd C_bl
Rb_35_76 bit_35_76 bit_35_77 R_bl
Rbb_35_76 bitb_35_76 bitb_35_77 R_bl
Cb_35_76 bit_35_76 gnd C_bl
Cbb_35_76 bitb_35_76 gnd C_bl
Rb_35_77 bit_35_77 bit_35_78 R_bl
Rbb_35_77 bitb_35_77 bitb_35_78 R_bl
Cb_35_77 bit_35_77 gnd C_bl
Cbb_35_77 bitb_35_77 gnd C_bl
Rb_35_78 bit_35_78 bit_35_79 R_bl
Rbb_35_78 bitb_35_78 bitb_35_79 R_bl
Cb_35_78 bit_35_78 gnd C_bl
Cbb_35_78 bitb_35_78 gnd C_bl
Rb_35_79 bit_35_79 bit_35_80 R_bl
Rbb_35_79 bitb_35_79 bitb_35_80 R_bl
Cb_35_79 bit_35_79 gnd C_bl
Cbb_35_79 bitb_35_79 gnd C_bl
Rb_35_80 bit_35_80 bit_35_81 R_bl
Rbb_35_80 bitb_35_80 bitb_35_81 R_bl
Cb_35_80 bit_35_80 gnd C_bl
Cbb_35_80 bitb_35_80 gnd C_bl
Rb_35_81 bit_35_81 bit_35_82 R_bl
Rbb_35_81 bitb_35_81 bitb_35_82 R_bl
Cb_35_81 bit_35_81 gnd C_bl
Cbb_35_81 bitb_35_81 gnd C_bl
Rb_35_82 bit_35_82 bit_35_83 R_bl
Rbb_35_82 bitb_35_82 bitb_35_83 R_bl
Cb_35_82 bit_35_82 gnd C_bl
Cbb_35_82 bitb_35_82 gnd C_bl
Rb_35_83 bit_35_83 bit_35_84 R_bl
Rbb_35_83 bitb_35_83 bitb_35_84 R_bl
Cb_35_83 bit_35_83 gnd C_bl
Cbb_35_83 bitb_35_83 gnd C_bl
Rb_35_84 bit_35_84 bit_35_85 R_bl
Rbb_35_84 bitb_35_84 bitb_35_85 R_bl
Cb_35_84 bit_35_84 gnd C_bl
Cbb_35_84 bitb_35_84 gnd C_bl
Rb_35_85 bit_35_85 bit_35_86 R_bl
Rbb_35_85 bitb_35_85 bitb_35_86 R_bl
Cb_35_85 bit_35_85 gnd C_bl
Cbb_35_85 bitb_35_85 gnd C_bl
Rb_35_86 bit_35_86 bit_35_87 R_bl
Rbb_35_86 bitb_35_86 bitb_35_87 R_bl
Cb_35_86 bit_35_86 gnd C_bl
Cbb_35_86 bitb_35_86 gnd C_bl
Rb_35_87 bit_35_87 bit_35_88 R_bl
Rbb_35_87 bitb_35_87 bitb_35_88 R_bl
Cb_35_87 bit_35_87 gnd C_bl
Cbb_35_87 bitb_35_87 gnd C_bl
Rb_35_88 bit_35_88 bit_35_89 R_bl
Rbb_35_88 bitb_35_88 bitb_35_89 R_bl
Cb_35_88 bit_35_88 gnd C_bl
Cbb_35_88 bitb_35_88 gnd C_bl
Rb_35_89 bit_35_89 bit_35_90 R_bl
Rbb_35_89 bitb_35_89 bitb_35_90 R_bl
Cb_35_89 bit_35_89 gnd C_bl
Cbb_35_89 bitb_35_89 gnd C_bl
Rb_35_90 bit_35_90 bit_35_91 R_bl
Rbb_35_90 bitb_35_90 bitb_35_91 R_bl
Cb_35_90 bit_35_90 gnd C_bl
Cbb_35_90 bitb_35_90 gnd C_bl
Rb_35_91 bit_35_91 bit_35_92 R_bl
Rbb_35_91 bitb_35_91 bitb_35_92 R_bl
Cb_35_91 bit_35_91 gnd C_bl
Cbb_35_91 bitb_35_91 gnd C_bl
Rb_35_92 bit_35_92 bit_35_93 R_bl
Rbb_35_92 bitb_35_92 bitb_35_93 R_bl
Cb_35_92 bit_35_92 gnd C_bl
Cbb_35_92 bitb_35_92 gnd C_bl
Rb_35_93 bit_35_93 bit_35_94 R_bl
Rbb_35_93 bitb_35_93 bitb_35_94 R_bl
Cb_35_93 bit_35_93 gnd C_bl
Cbb_35_93 bitb_35_93 gnd C_bl
Rb_35_94 bit_35_94 bit_35_95 R_bl
Rbb_35_94 bitb_35_94 bitb_35_95 R_bl
Cb_35_94 bit_35_94 gnd C_bl
Cbb_35_94 bitb_35_94 gnd C_bl
Rb_35_95 bit_35_95 bit_35_96 R_bl
Rbb_35_95 bitb_35_95 bitb_35_96 R_bl
Cb_35_95 bit_35_95 gnd C_bl
Cbb_35_95 bitb_35_95 gnd C_bl
Rb_35_96 bit_35_96 bit_35_97 R_bl
Rbb_35_96 bitb_35_96 bitb_35_97 R_bl
Cb_35_96 bit_35_96 gnd C_bl
Cbb_35_96 bitb_35_96 gnd C_bl
Rb_35_97 bit_35_97 bit_35_98 R_bl
Rbb_35_97 bitb_35_97 bitb_35_98 R_bl
Cb_35_97 bit_35_97 gnd C_bl
Cbb_35_97 bitb_35_97 gnd C_bl
Rb_35_98 bit_35_98 bit_35_99 R_bl
Rbb_35_98 bitb_35_98 bitb_35_99 R_bl
Cb_35_98 bit_35_98 gnd C_bl
Cbb_35_98 bitb_35_98 gnd C_bl
Rb_35_99 bit_35_99 bit_35_100 R_bl
Rbb_35_99 bitb_35_99 bitb_35_100 R_bl
Cb_35_99 bit_35_99 gnd C_bl
Cbb_35_99 bitb_35_99 gnd C_bl
Rb_36_0 bit_36_0 bit_36_1 R_bl
Rbb_36_0 bitb_36_0 bitb_36_1 R_bl
Cb_36_0 bit_36_0 gnd C_bl
Cbb_36_0 bitb_36_0 gnd C_bl
Rb_36_1 bit_36_1 bit_36_2 R_bl
Rbb_36_1 bitb_36_1 bitb_36_2 R_bl
Cb_36_1 bit_36_1 gnd C_bl
Cbb_36_1 bitb_36_1 gnd C_bl
Rb_36_2 bit_36_2 bit_36_3 R_bl
Rbb_36_2 bitb_36_2 bitb_36_3 R_bl
Cb_36_2 bit_36_2 gnd C_bl
Cbb_36_2 bitb_36_2 gnd C_bl
Rb_36_3 bit_36_3 bit_36_4 R_bl
Rbb_36_3 bitb_36_3 bitb_36_4 R_bl
Cb_36_3 bit_36_3 gnd C_bl
Cbb_36_3 bitb_36_3 gnd C_bl
Rb_36_4 bit_36_4 bit_36_5 R_bl
Rbb_36_4 bitb_36_4 bitb_36_5 R_bl
Cb_36_4 bit_36_4 gnd C_bl
Cbb_36_4 bitb_36_4 gnd C_bl
Rb_36_5 bit_36_5 bit_36_6 R_bl
Rbb_36_5 bitb_36_5 bitb_36_6 R_bl
Cb_36_5 bit_36_5 gnd C_bl
Cbb_36_5 bitb_36_5 gnd C_bl
Rb_36_6 bit_36_6 bit_36_7 R_bl
Rbb_36_6 bitb_36_6 bitb_36_7 R_bl
Cb_36_6 bit_36_6 gnd C_bl
Cbb_36_6 bitb_36_6 gnd C_bl
Rb_36_7 bit_36_7 bit_36_8 R_bl
Rbb_36_7 bitb_36_7 bitb_36_8 R_bl
Cb_36_7 bit_36_7 gnd C_bl
Cbb_36_7 bitb_36_7 gnd C_bl
Rb_36_8 bit_36_8 bit_36_9 R_bl
Rbb_36_8 bitb_36_8 bitb_36_9 R_bl
Cb_36_8 bit_36_8 gnd C_bl
Cbb_36_8 bitb_36_8 gnd C_bl
Rb_36_9 bit_36_9 bit_36_10 R_bl
Rbb_36_9 bitb_36_9 bitb_36_10 R_bl
Cb_36_9 bit_36_9 gnd C_bl
Cbb_36_9 bitb_36_9 gnd C_bl
Rb_36_10 bit_36_10 bit_36_11 R_bl
Rbb_36_10 bitb_36_10 bitb_36_11 R_bl
Cb_36_10 bit_36_10 gnd C_bl
Cbb_36_10 bitb_36_10 gnd C_bl
Rb_36_11 bit_36_11 bit_36_12 R_bl
Rbb_36_11 bitb_36_11 bitb_36_12 R_bl
Cb_36_11 bit_36_11 gnd C_bl
Cbb_36_11 bitb_36_11 gnd C_bl
Rb_36_12 bit_36_12 bit_36_13 R_bl
Rbb_36_12 bitb_36_12 bitb_36_13 R_bl
Cb_36_12 bit_36_12 gnd C_bl
Cbb_36_12 bitb_36_12 gnd C_bl
Rb_36_13 bit_36_13 bit_36_14 R_bl
Rbb_36_13 bitb_36_13 bitb_36_14 R_bl
Cb_36_13 bit_36_13 gnd C_bl
Cbb_36_13 bitb_36_13 gnd C_bl
Rb_36_14 bit_36_14 bit_36_15 R_bl
Rbb_36_14 bitb_36_14 bitb_36_15 R_bl
Cb_36_14 bit_36_14 gnd C_bl
Cbb_36_14 bitb_36_14 gnd C_bl
Rb_36_15 bit_36_15 bit_36_16 R_bl
Rbb_36_15 bitb_36_15 bitb_36_16 R_bl
Cb_36_15 bit_36_15 gnd C_bl
Cbb_36_15 bitb_36_15 gnd C_bl
Rb_36_16 bit_36_16 bit_36_17 R_bl
Rbb_36_16 bitb_36_16 bitb_36_17 R_bl
Cb_36_16 bit_36_16 gnd C_bl
Cbb_36_16 bitb_36_16 gnd C_bl
Rb_36_17 bit_36_17 bit_36_18 R_bl
Rbb_36_17 bitb_36_17 bitb_36_18 R_bl
Cb_36_17 bit_36_17 gnd C_bl
Cbb_36_17 bitb_36_17 gnd C_bl
Rb_36_18 bit_36_18 bit_36_19 R_bl
Rbb_36_18 bitb_36_18 bitb_36_19 R_bl
Cb_36_18 bit_36_18 gnd C_bl
Cbb_36_18 bitb_36_18 gnd C_bl
Rb_36_19 bit_36_19 bit_36_20 R_bl
Rbb_36_19 bitb_36_19 bitb_36_20 R_bl
Cb_36_19 bit_36_19 gnd C_bl
Cbb_36_19 bitb_36_19 gnd C_bl
Rb_36_20 bit_36_20 bit_36_21 R_bl
Rbb_36_20 bitb_36_20 bitb_36_21 R_bl
Cb_36_20 bit_36_20 gnd C_bl
Cbb_36_20 bitb_36_20 gnd C_bl
Rb_36_21 bit_36_21 bit_36_22 R_bl
Rbb_36_21 bitb_36_21 bitb_36_22 R_bl
Cb_36_21 bit_36_21 gnd C_bl
Cbb_36_21 bitb_36_21 gnd C_bl
Rb_36_22 bit_36_22 bit_36_23 R_bl
Rbb_36_22 bitb_36_22 bitb_36_23 R_bl
Cb_36_22 bit_36_22 gnd C_bl
Cbb_36_22 bitb_36_22 gnd C_bl
Rb_36_23 bit_36_23 bit_36_24 R_bl
Rbb_36_23 bitb_36_23 bitb_36_24 R_bl
Cb_36_23 bit_36_23 gnd C_bl
Cbb_36_23 bitb_36_23 gnd C_bl
Rb_36_24 bit_36_24 bit_36_25 R_bl
Rbb_36_24 bitb_36_24 bitb_36_25 R_bl
Cb_36_24 bit_36_24 gnd C_bl
Cbb_36_24 bitb_36_24 gnd C_bl
Rb_36_25 bit_36_25 bit_36_26 R_bl
Rbb_36_25 bitb_36_25 bitb_36_26 R_bl
Cb_36_25 bit_36_25 gnd C_bl
Cbb_36_25 bitb_36_25 gnd C_bl
Rb_36_26 bit_36_26 bit_36_27 R_bl
Rbb_36_26 bitb_36_26 bitb_36_27 R_bl
Cb_36_26 bit_36_26 gnd C_bl
Cbb_36_26 bitb_36_26 gnd C_bl
Rb_36_27 bit_36_27 bit_36_28 R_bl
Rbb_36_27 bitb_36_27 bitb_36_28 R_bl
Cb_36_27 bit_36_27 gnd C_bl
Cbb_36_27 bitb_36_27 gnd C_bl
Rb_36_28 bit_36_28 bit_36_29 R_bl
Rbb_36_28 bitb_36_28 bitb_36_29 R_bl
Cb_36_28 bit_36_28 gnd C_bl
Cbb_36_28 bitb_36_28 gnd C_bl
Rb_36_29 bit_36_29 bit_36_30 R_bl
Rbb_36_29 bitb_36_29 bitb_36_30 R_bl
Cb_36_29 bit_36_29 gnd C_bl
Cbb_36_29 bitb_36_29 gnd C_bl
Rb_36_30 bit_36_30 bit_36_31 R_bl
Rbb_36_30 bitb_36_30 bitb_36_31 R_bl
Cb_36_30 bit_36_30 gnd C_bl
Cbb_36_30 bitb_36_30 gnd C_bl
Rb_36_31 bit_36_31 bit_36_32 R_bl
Rbb_36_31 bitb_36_31 bitb_36_32 R_bl
Cb_36_31 bit_36_31 gnd C_bl
Cbb_36_31 bitb_36_31 gnd C_bl
Rb_36_32 bit_36_32 bit_36_33 R_bl
Rbb_36_32 bitb_36_32 bitb_36_33 R_bl
Cb_36_32 bit_36_32 gnd C_bl
Cbb_36_32 bitb_36_32 gnd C_bl
Rb_36_33 bit_36_33 bit_36_34 R_bl
Rbb_36_33 bitb_36_33 bitb_36_34 R_bl
Cb_36_33 bit_36_33 gnd C_bl
Cbb_36_33 bitb_36_33 gnd C_bl
Rb_36_34 bit_36_34 bit_36_35 R_bl
Rbb_36_34 bitb_36_34 bitb_36_35 R_bl
Cb_36_34 bit_36_34 gnd C_bl
Cbb_36_34 bitb_36_34 gnd C_bl
Rb_36_35 bit_36_35 bit_36_36 R_bl
Rbb_36_35 bitb_36_35 bitb_36_36 R_bl
Cb_36_35 bit_36_35 gnd C_bl
Cbb_36_35 bitb_36_35 gnd C_bl
Rb_36_36 bit_36_36 bit_36_37 R_bl
Rbb_36_36 bitb_36_36 bitb_36_37 R_bl
Cb_36_36 bit_36_36 gnd C_bl
Cbb_36_36 bitb_36_36 gnd C_bl
Rb_36_37 bit_36_37 bit_36_38 R_bl
Rbb_36_37 bitb_36_37 bitb_36_38 R_bl
Cb_36_37 bit_36_37 gnd C_bl
Cbb_36_37 bitb_36_37 gnd C_bl
Rb_36_38 bit_36_38 bit_36_39 R_bl
Rbb_36_38 bitb_36_38 bitb_36_39 R_bl
Cb_36_38 bit_36_38 gnd C_bl
Cbb_36_38 bitb_36_38 gnd C_bl
Rb_36_39 bit_36_39 bit_36_40 R_bl
Rbb_36_39 bitb_36_39 bitb_36_40 R_bl
Cb_36_39 bit_36_39 gnd C_bl
Cbb_36_39 bitb_36_39 gnd C_bl
Rb_36_40 bit_36_40 bit_36_41 R_bl
Rbb_36_40 bitb_36_40 bitb_36_41 R_bl
Cb_36_40 bit_36_40 gnd C_bl
Cbb_36_40 bitb_36_40 gnd C_bl
Rb_36_41 bit_36_41 bit_36_42 R_bl
Rbb_36_41 bitb_36_41 bitb_36_42 R_bl
Cb_36_41 bit_36_41 gnd C_bl
Cbb_36_41 bitb_36_41 gnd C_bl
Rb_36_42 bit_36_42 bit_36_43 R_bl
Rbb_36_42 bitb_36_42 bitb_36_43 R_bl
Cb_36_42 bit_36_42 gnd C_bl
Cbb_36_42 bitb_36_42 gnd C_bl
Rb_36_43 bit_36_43 bit_36_44 R_bl
Rbb_36_43 bitb_36_43 bitb_36_44 R_bl
Cb_36_43 bit_36_43 gnd C_bl
Cbb_36_43 bitb_36_43 gnd C_bl
Rb_36_44 bit_36_44 bit_36_45 R_bl
Rbb_36_44 bitb_36_44 bitb_36_45 R_bl
Cb_36_44 bit_36_44 gnd C_bl
Cbb_36_44 bitb_36_44 gnd C_bl
Rb_36_45 bit_36_45 bit_36_46 R_bl
Rbb_36_45 bitb_36_45 bitb_36_46 R_bl
Cb_36_45 bit_36_45 gnd C_bl
Cbb_36_45 bitb_36_45 gnd C_bl
Rb_36_46 bit_36_46 bit_36_47 R_bl
Rbb_36_46 bitb_36_46 bitb_36_47 R_bl
Cb_36_46 bit_36_46 gnd C_bl
Cbb_36_46 bitb_36_46 gnd C_bl
Rb_36_47 bit_36_47 bit_36_48 R_bl
Rbb_36_47 bitb_36_47 bitb_36_48 R_bl
Cb_36_47 bit_36_47 gnd C_bl
Cbb_36_47 bitb_36_47 gnd C_bl
Rb_36_48 bit_36_48 bit_36_49 R_bl
Rbb_36_48 bitb_36_48 bitb_36_49 R_bl
Cb_36_48 bit_36_48 gnd C_bl
Cbb_36_48 bitb_36_48 gnd C_bl
Rb_36_49 bit_36_49 bit_36_50 R_bl
Rbb_36_49 bitb_36_49 bitb_36_50 R_bl
Cb_36_49 bit_36_49 gnd C_bl
Cbb_36_49 bitb_36_49 gnd C_bl
Rb_36_50 bit_36_50 bit_36_51 R_bl
Rbb_36_50 bitb_36_50 bitb_36_51 R_bl
Cb_36_50 bit_36_50 gnd C_bl
Cbb_36_50 bitb_36_50 gnd C_bl
Rb_36_51 bit_36_51 bit_36_52 R_bl
Rbb_36_51 bitb_36_51 bitb_36_52 R_bl
Cb_36_51 bit_36_51 gnd C_bl
Cbb_36_51 bitb_36_51 gnd C_bl
Rb_36_52 bit_36_52 bit_36_53 R_bl
Rbb_36_52 bitb_36_52 bitb_36_53 R_bl
Cb_36_52 bit_36_52 gnd C_bl
Cbb_36_52 bitb_36_52 gnd C_bl
Rb_36_53 bit_36_53 bit_36_54 R_bl
Rbb_36_53 bitb_36_53 bitb_36_54 R_bl
Cb_36_53 bit_36_53 gnd C_bl
Cbb_36_53 bitb_36_53 gnd C_bl
Rb_36_54 bit_36_54 bit_36_55 R_bl
Rbb_36_54 bitb_36_54 bitb_36_55 R_bl
Cb_36_54 bit_36_54 gnd C_bl
Cbb_36_54 bitb_36_54 gnd C_bl
Rb_36_55 bit_36_55 bit_36_56 R_bl
Rbb_36_55 bitb_36_55 bitb_36_56 R_bl
Cb_36_55 bit_36_55 gnd C_bl
Cbb_36_55 bitb_36_55 gnd C_bl
Rb_36_56 bit_36_56 bit_36_57 R_bl
Rbb_36_56 bitb_36_56 bitb_36_57 R_bl
Cb_36_56 bit_36_56 gnd C_bl
Cbb_36_56 bitb_36_56 gnd C_bl
Rb_36_57 bit_36_57 bit_36_58 R_bl
Rbb_36_57 bitb_36_57 bitb_36_58 R_bl
Cb_36_57 bit_36_57 gnd C_bl
Cbb_36_57 bitb_36_57 gnd C_bl
Rb_36_58 bit_36_58 bit_36_59 R_bl
Rbb_36_58 bitb_36_58 bitb_36_59 R_bl
Cb_36_58 bit_36_58 gnd C_bl
Cbb_36_58 bitb_36_58 gnd C_bl
Rb_36_59 bit_36_59 bit_36_60 R_bl
Rbb_36_59 bitb_36_59 bitb_36_60 R_bl
Cb_36_59 bit_36_59 gnd C_bl
Cbb_36_59 bitb_36_59 gnd C_bl
Rb_36_60 bit_36_60 bit_36_61 R_bl
Rbb_36_60 bitb_36_60 bitb_36_61 R_bl
Cb_36_60 bit_36_60 gnd C_bl
Cbb_36_60 bitb_36_60 gnd C_bl
Rb_36_61 bit_36_61 bit_36_62 R_bl
Rbb_36_61 bitb_36_61 bitb_36_62 R_bl
Cb_36_61 bit_36_61 gnd C_bl
Cbb_36_61 bitb_36_61 gnd C_bl
Rb_36_62 bit_36_62 bit_36_63 R_bl
Rbb_36_62 bitb_36_62 bitb_36_63 R_bl
Cb_36_62 bit_36_62 gnd C_bl
Cbb_36_62 bitb_36_62 gnd C_bl
Rb_36_63 bit_36_63 bit_36_64 R_bl
Rbb_36_63 bitb_36_63 bitb_36_64 R_bl
Cb_36_63 bit_36_63 gnd C_bl
Cbb_36_63 bitb_36_63 gnd C_bl
Rb_36_64 bit_36_64 bit_36_65 R_bl
Rbb_36_64 bitb_36_64 bitb_36_65 R_bl
Cb_36_64 bit_36_64 gnd C_bl
Cbb_36_64 bitb_36_64 gnd C_bl
Rb_36_65 bit_36_65 bit_36_66 R_bl
Rbb_36_65 bitb_36_65 bitb_36_66 R_bl
Cb_36_65 bit_36_65 gnd C_bl
Cbb_36_65 bitb_36_65 gnd C_bl
Rb_36_66 bit_36_66 bit_36_67 R_bl
Rbb_36_66 bitb_36_66 bitb_36_67 R_bl
Cb_36_66 bit_36_66 gnd C_bl
Cbb_36_66 bitb_36_66 gnd C_bl
Rb_36_67 bit_36_67 bit_36_68 R_bl
Rbb_36_67 bitb_36_67 bitb_36_68 R_bl
Cb_36_67 bit_36_67 gnd C_bl
Cbb_36_67 bitb_36_67 gnd C_bl
Rb_36_68 bit_36_68 bit_36_69 R_bl
Rbb_36_68 bitb_36_68 bitb_36_69 R_bl
Cb_36_68 bit_36_68 gnd C_bl
Cbb_36_68 bitb_36_68 gnd C_bl
Rb_36_69 bit_36_69 bit_36_70 R_bl
Rbb_36_69 bitb_36_69 bitb_36_70 R_bl
Cb_36_69 bit_36_69 gnd C_bl
Cbb_36_69 bitb_36_69 gnd C_bl
Rb_36_70 bit_36_70 bit_36_71 R_bl
Rbb_36_70 bitb_36_70 bitb_36_71 R_bl
Cb_36_70 bit_36_70 gnd C_bl
Cbb_36_70 bitb_36_70 gnd C_bl
Rb_36_71 bit_36_71 bit_36_72 R_bl
Rbb_36_71 bitb_36_71 bitb_36_72 R_bl
Cb_36_71 bit_36_71 gnd C_bl
Cbb_36_71 bitb_36_71 gnd C_bl
Rb_36_72 bit_36_72 bit_36_73 R_bl
Rbb_36_72 bitb_36_72 bitb_36_73 R_bl
Cb_36_72 bit_36_72 gnd C_bl
Cbb_36_72 bitb_36_72 gnd C_bl
Rb_36_73 bit_36_73 bit_36_74 R_bl
Rbb_36_73 bitb_36_73 bitb_36_74 R_bl
Cb_36_73 bit_36_73 gnd C_bl
Cbb_36_73 bitb_36_73 gnd C_bl
Rb_36_74 bit_36_74 bit_36_75 R_bl
Rbb_36_74 bitb_36_74 bitb_36_75 R_bl
Cb_36_74 bit_36_74 gnd C_bl
Cbb_36_74 bitb_36_74 gnd C_bl
Rb_36_75 bit_36_75 bit_36_76 R_bl
Rbb_36_75 bitb_36_75 bitb_36_76 R_bl
Cb_36_75 bit_36_75 gnd C_bl
Cbb_36_75 bitb_36_75 gnd C_bl
Rb_36_76 bit_36_76 bit_36_77 R_bl
Rbb_36_76 bitb_36_76 bitb_36_77 R_bl
Cb_36_76 bit_36_76 gnd C_bl
Cbb_36_76 bitb_36_76 gnd C_bl
Rb_36_77 bit_36_77 bit_36_78 R_bl
Rbb_36_77 bitb_36_77 bitb_36_78 R_bl
Cb_36_77 bit_36_77 gnd C_bl
Cbb_36_77 bitb_36_77 gnd C_bl
Rb_36_78 bit_36_78 bit_36_79 R_bl
Rbb_36_78 bitb_36_78 bitb_36_79 R_bl
Cb_36_78 bit_36_78 gnd C_bl
Cbb_36_78 bitb_36_78 gnd C_bl
Rb_36_79 bit_36_79 bit_36_80 R_bl
Rbb_36_79 bitb_36_79 bitb_36_80 R_bl
Cb_36_79 bit_36_79 gnd C_bl
Cbb_36_79 bitb_36_79 gnd C_bl
Rb_36_80 bit_36_80 bit_36_81 R_bl
Rbb_36_80 bitb_36_80 bitb_36_81 R_bl
Cb_36_80 bit_36_80 gnd C_bl
Cbb_36_80 bitb_36_80 gnd C_bl
Rb_36_81 bit_36_81 bit_36_82 R_bl
Rbb_36_81 bitb_36_81 bitb_36_82 R_bl
Cb_36_81 bit_36_81 gnd C_bl
Cbb_36_81 bitb_36_81 gnd C_bl
Rb_36_82 bit_36_82 bit_36_83 R_bl
Rbb_36_82 bitb_36_82 bitb_36_83 R_bl
Cb_36_82 bit_36_82 gnd C_bl
Cbb_36_82 bitb_36_82 gnd C_bl
Rb_36_83 bit_36_83 bit_36_84 R_bl
Rbb_36_83 bitb_36_83 bitb_36_84 R_bl
Cb_36_83 bit_36_83 gnd C_bl
Cbb_36_83 bitb_36_83 gnd C_bl
Rb_36_84 bit_36_84 bit_36_85 R_bl
Rbb_36_84 bitb_36_84 bitb_36_85 R_bl
Cb_36_84 bit_36_84 gnd C_bl
Cbb_36_84 bitb_36_84 gnd C_bl
Rb_36_85 bit_36_85 bit_36_86 R_bl
Rbb_36_85 bitb_36_85 bitb_36_86 R_bl
Cb_36_85 bit_36_85 gnd C_bl
Cbb_36_85 bitb_36_85 gnd C_bl
Rb_36_86 bit_36_86 bit_36_87 R_bl
Rbb_36_86 bitb_36_86 bitb_36_87 R_bl
Cb_36_86 bit_36_86 gnd C_bl
Cbb_36_86 bitb_36_86 gnd C_bl
Rb_36_87 bit_36_87 bit_36_88 R_bl
Rbb_36_87 bitb_36_87 bitb_36_88 R_bl
Cb_36_87 bit_36_87 gnd C_bl
Cbb_36_87 bitb_36_87 gnd C_bl
Rb_36_88 bit_36_88 bit_36_89 R_bl
Rbb_36_88 bitb_36_88 bitb_36_89 R_bl
Cb_36_88 bit_36_88 gnd C_bl
Cbb_36_88 bitb_36_88 gnd C_bl
Rb_36_89 bit_36_89 bit_36_90 R_bl
Rbb_36_89 bitb_36_89 bitb_36_90 R_bl
Cb_36_89 bit_36_89 gnd C_bl
Cbb_36_89 bitb_36_89 gnd C_bl
Rb_36_90 bit_36_90 bit_36_91 R_bl
Rbb_36_90 bitb_36_90 bitb_36_91 R_bl
Cb_36_90 bit_36_90 gnd C_bl
Cbb_36_90 bitb_36_90 gnd C_bl
Rb_36_91 bit_36_91 bit_36_92 R_bl
Rbb_36_91 bitb_36_91 bitb_36_92 R_bl
Cb_36_91 bit_36_91 gnd C_bl
Cbb_36_91 bitb_36_91 gnd C_bl
Rb_36_92 bit_36_92 bit_36_93 R_bl
Rbb_36_92 bitb_36_92 bitb_36_93 R_bl
Cb_36_92 bit_36_92 gnd C_bl
Cbb_36_92 bitb_36_92 gnd C_bl
Rb_36_93 bit_36_93 bit_36_94 R_bl
Rbb_36_93 bitb_36_93 bitb_36_94 R_bl
Cb_36_93 bit_36_93 gnd C_bl
Cbb_36_93 bitb_36_93 gnd C_bl
Rb_36_94 bit_36_94 bit_36_95 R_bl
Rbb_36_94 bitb_36_94 bitb_36_95 R_bl
Cb_36_94 bit_36_94 gnd C_bl
Cbb_36_94 bitb_36_94 gnd C_bl
Rb_36_95 bit_36_95 bit_36_96 R_bl
Rbb_36_95 bitb_36_95 bitb_36_96 R_bl
Cb_36_95 bit_36_95 gnd C_bl
Cbb_36_95 bitb_36_95 gnd C_bl
Rb_36_96 bit_36_96 bit_36_97 R_bl
Rbb_36_96 bitb_36_96 bitb_36_97 R_bl
Cb_36_96 bit_36_96 gnd C_bl
Cbb_36_96 bitb_36_96 gnd C_bl
Rb_36_97 bit_36_97 bit_36_98 R_bl
Rbb_36_97 bitb_36_97 bitb_36_98 R_bl
Cb_36_97 bit_36_97 gnd C_bl
Cbb_36_97 bitb_36_97 gnd C_bl
Rb_36_98 bit_36_98 bit_36_99 R_bl
Rbb_36_98 bitb_36_98 bitb_36_99 R_bl
Cb_36_98 bit_36_98 gnd C_bl
Cbb_36_98 bitb_36_98 gnd C_bl
Rb_36_99 bit_36_99 bit_36_100 R_bl
Rbb_36_99 bitb_36_99 bitb_36_100 R_bl
Cb_36_99 bit_36_99 gnd C_bl
Cbb_36_99 bitb_36_99 gnd C_bl
Rb_37_0 bit_37_0 bit_37_1 R_bl
Rbb_37_0 bitb_37_0 bitb_37_1 R_bl
Cb_37_0 bit_37_0 gnd C_bl
Cbb_37_0 bitb_37_0 gnd C_bl
Rb_37_1 bit_37_1 bit_37_2 R_bl
Rbb_37_1 bitb_37_1 bitb_37_2 R_bl
Cb_37_1 bit_37_1 gnd C_bl
Cbb_37_1 bitb_37_1 gnd C_bl
Rb_37_2 bit_37_2 bit_37_3 R_bl
Rbb_37_2 bitb_37_2 bitb_37_3 R_bl
Cb_37_2 bit_37_2 gnd C_bl
Cbb_37_2 bitb_37_2 gnd C_bl
Rb_37_3 bit_37_3 bit_37_4 R_bl
Rbb_37_3 bitb_37_3 bitb_37_4 R_bl
Cb_37_3 bit_37_3 gnd C_bl
Cbb_37_3 bitb_37_3 gnd C_bl
Rb_37_4 bit_37_4 bit_37_5 R_bl
Rbb_37_4 bitb_37_4 bitb_37_5 R_bl
Cb_37_4 bit_37_4 gnd C_bl
Cbb_37_4 bitb_37_4 gnd C_bl
Rb_37_5 bit_37_5 bit_37_6 R_bl
Rbb_37_5 bitb_37_5 bitb_37_6 R_bl
Cb_37_5 bit_37_5 gnd C_bl
Cbb_37_5 bitb_37_5 gnd C_bl
Rb_37_6 bit_37_6 bit_37_7 R_bl
Rbb_37_6 bitb_37_6 bitb_37_7 R_bl
Cb_37_6 bit_37_6 gnd C_bl
Cbb_37_6 bitb_37_6 gnd C_bl
Rb_37_7 bit_37_7 bit_37_8 R_bl
Rbb_37_7 bitb_37_7 bitb_37_8 R_bl
Cb_37_7 bit_37_7 gnd C_bl
Cbb_37_7 bitb_37_7 gnd C_bl
Rb_37_8 bit_37_8 bit_37_9 R_bl
Rbb_37_8 bitb_37_8 bitb_37_9 R_bl
Cb_37_8 bit_37_8 gnd C_bl
Cbb_37_8 bitb_37_8 gnd C_bl
Rb_37_9 bit_37_9 bit_37_10 R_bl
Rbb_37_9 bitb_37_9 bitb_37_10 R_bl
Cb_37_9 bit_37_9 gnd C_bl
Cbb_37_9 bitb_37_9 gnd C_bl
Rb_37_10 bit_37_10 bit_37_11 R_bl
Rbb_37_10 bitb_37_10 bitb_37_11 R_bl
Cb_37_10 bit_37_10 gnd C_bl
Cbb_37_10 bitb_37_10 gnd C_bl
Rb_37_11 bit_37_11 bit_37_12 R_bl
Rbb_37_11 bitb_37_11 bitb_37_12 R_bl
Cb_37_11 bit_37_11 gnd C_bl
Cbb_37_11 bitb_37_11 gnd C_bl
Rb_37_12 bit_37_12 bit_37_13 R_bl
Rbb_37_12 bitb_37_12 bitb_37_13 R_bl
Cb_37_12 bit_37_12 gnd C_bl
Cbb_37_12 bitb_37_12 gnd C_bl
Rb_37_13 bit_37_13 bit_37_14 R_bl
Rbb_37_13 bitb_37_13 bitb_37_14 R_bl
Cb_37_13 bit_37_13 gnd C_bl
Cbb_37_13 bitb_37_13 gnd C_bl
Rb_37_14 bit_37_14 bit_37_15 R_bl
Rbb_37_14 bitb_37_14 bitb_37_15 R_bl
Cb_37_14 bit_37_14 gnd C_bl
Cbb_37_14 bitb_37_14 gnd C_bl
Rb_37_15 bit_37_15 bit_37_16 R_bl
Rbb_37_15 bitb_37_15 bitb_37_16 R_bl
Cb_37_15 bit_37_15 gnd C_bl
Cbb_37_15 bitb_37_15 gnd C_bl
Rb_37_16 bit_37_16 bit_37_17 R_bl
Rbb_37_16 bitb_37_16 bitb_37_17 R_bl
Cb_37_16 bit_37_16 gnd C_bl
Cbb_37_16 bitb_37_16 gnd C_bl
Rb_37_17 bit_37_17 bit_37_18 R_bl
Rbb_37_17 bitb_37_17 bitb_37_18 R_bl
Cb_37_17 bit_37_17 gnd C_bl
Cbb_37_17 bitb_37_17 gnd C_bl
Rb_37_18 bit_37_18 bit_37_19 R_bl
Rbb_37_18 bitb_37_18 bitb_37_19 R_bl
Cb_37_18 bit_37_18 gnd C_bl
Cbb_37_18 bitb_37_18 gnd C_bl
Rb_37_19 bit_37_19 bit_37_20 R_bl
Rbb_37_19 bitb_37_19 bitb_37_20 R_bl
Cb_37_19 bit_37_19 gnd C_bl
Cbb_37_19 bitb_37_19 gnd C_bl
Rb_37_20 bit_37_20 bit_37_21 R_bl
Rbb_37_20 bitb_37_20 bitb_37_21 R_bl
Cb_37_20 bit_37_20 gnd C_bl
Cbb_37_20 bitb_37_20 gnd C_bl
Rb_37_21 bit_37_21 bit_37_22 R_bl
Rbb_37_21 bitb_37_21 bitb_37_22 R_bl
Cb_37_21 bit_37_21 gnd C_bl
Cbb_37_21 bitb_37_21 gnd C_bl
Rb_37_22 bit_37_22 bit_37_23 R_bl
Rbb_37_22 bitb_37_22 bitb_37_23 R_bl
Cb_37_22 bit_37_22 gnd C_bl
Cbb_37_22 bitb_37_22 gnd C_bl
Rb_37_23 bit_37_23 bit_37_24 R_bl
Rbb_37_23 bitb_37_23 bitb_37_24 R_bl
Cb_37_23 bit_37_23 gnd C_bl
Cbb_37_23 bitb_37_23 gnd C_bl
Rb_37_24 bit_37_24 bit_37_25 R_bl
Rbb_37_24 bitb_37_24 bitb_37_25 R_bl
Cb_37_24 bit_37_24 gnd C_bl
Cbb_37_24 bitb_37_24 gnd C_bl
Rb_37_25 bit_37_25 bit_37_26 R_bl
Rbb_37_25 bitb_37_25 bitb_37_26 R_bl
Cb_37_25 bit_37_25 gnd C_bl
Cbb_37_25 bitb_37_25 gnd C_bl
Rb_37_26 bit_37_26 bit_37_27 R_bl
Rbb_37_26 bitb_37_26 bitb_37_27 R_bl
Cb_37_26 bit_37_26 gnd C_bl
Cbb_37_26 bitb_37_26 gnd C_bl
Rb_37_27 bit_37_27 bit_37_28 R_bl
Rbb_37_27 bitb_37_27 bitb_37_28 R_bl
Cb_37_27 bit_37_27 gnd C_bl
Cbb_37_27 bitb_37_27 gnd C_bl
Rb_37_28 bit_37_28 bit_37_29 R_bl
Rbb_37_28 bitb_37_28 bitb_37_29 R_bl
Cb_37_28 bit_37_28 gnd C_bl
Cbb_37_28 bitb_37_28 gnd C_bl
Rb_37_29 bit_37_29 bit_37_30 R_bl
Rbb_37_29 bitb_37_29 bitb_37_30 R_bl
Cb_37_29 bit_37_29 gnd C_bl
Cbb_37_29 bitb_37_29 gnd C_bl
Rb_37_30 bit_37_30 bit_37_31 R_bl
Rbb_37_30 bitb_37_30 bitb_37_31 R_bl
Cb_37_30 bit_37_30 gnd C_bl
Cbb_37_30 bitb_37_30 gnd C_bl
Rb_37_31 bit_37_31 bit_37_32 R_bl
Rbb_37_31 bitb_37_31 bitb_37_32 R_bl
Cb_37_31 bit_37_31 gnd C_bl
Cbb_37_31 bitb_37_31 gnd C_bl
Rb_37_32 bit_37_32 bit_37_33 R_bl
Rbb_37_32 bitb_37_32 bitb_37_33 R_bl
Cb_37_32 bit_37_32 gnd C_bl
Cbb_37_32 bitb_37_32 gnd C_bl
Rb_37_33 bit_37_33 bit_37_34 R_bl
Rbb_37_33 bitb_37_33 bitb_37_34 R_bl
Cb_37_33 bit_37_33 gnd C_bl
Cbb_37_33 bitb_37_33 gnd C_bl
Rb_37_34 bit_37_34 bit_37_35 R_bl
Rbb_37_34 bitb_37_34 bitb_37_35 R_bl
Cb_37_34 bit_37_34 gnd C_bl
Cbb_37_34 bitb_37_34 gnd C_bl
Rb_37_35 bit_37_35 bit_37_36 R_bl
Rbb_37_35 bitb_37_35 bitb_37_36 R_bl
Cb_37_35 bit_37_35 gnd C_bl
Cbb_37_35 bitb_37_35 gnd C_bl
Rb_37_36 bit_37_36 bit_37_37 R_bl
Rbb_37_36 bitb_37_36 bitb_37_37 R_bl
Cb_37_36 bit_37_36 gnd C_bl
Cbb_37_36 bitb_37_36 gnd C_bl
Rb_37_37 bit_37_37 bit_37_38 R_bl
Rbb_37_37 bitb_37_37 bitb_37_38 R_bl
Cb_37_37 bit_37_37 gnd C_bl
Cbb_37_37 bitb_37_37 gnd C_bl
Rb_37_38 bit_37_38 bit_37_39 R_bl
Rbb_37_38 bitb_37_38 bitb_37_39 R_bl
Cb_37_38 bit_37_38 gnd C_bl
Cbb_37_38 bitb_37_38 gnd C_bl
Rb_37_39 bit_37_39 bit_37_40 R_bl
Rbb_37_39 bitb_37_39 bitb_37_40 R_bl
Cb_37_39 bit_37_39 gnd C_bl
Cbb_37_39 bitb_37_39 gnd C_bl
Rb_37_40 bit_37_40 bit_37_41 R_bl
Rbb_37_40 bitb_37_40 bitb_37_41 R_bl
Cb_37_40 bit_37_40 gnd C_bl
Cbb_37_40 bitb_37_40 gnd C_bl
Rb_37_41 bit_37_41 bit_37_42 R_bl
Rbb_37_41 bitb_37_41 bitb_37_42 R_bl
Cb_37_41 bit_37_41 gnd C_bl
Cbb_37_41 bitb_37_41 gnd C_bl
Rb_37_42 bit_37_42 bit_37_43 R_bl
Rbb_37_42 bitb_37_42 bitb_37_43 R_bl
Cb_37_42 bit_37_42 gnd C_bl
Cbb_37_42 bitb_37_42 gnd C_bl
Rb_37_43 bit_37_43 bit_37_44 R_bl
Rbb_37_43 bitb_37_43 bitb_37_44 R_bl
Cb_37_43 bit_37_43 gnd C_bl
Cbb_37_43 bitb_37_43 gnd C_bl
Rb_37_44 bit_37_44 bit_37_45 R_bl
Rbb_37_44 bitb_37_44 bitb_37_45 R_bl
Cb_37_44 bit_37_44 gnd C_bl
Cbb_37_44 bitb_37_44 gnd C_bl
Rb_37_45 bit_37_45 bit_37_46 R_bl
Rbb_37_45 bitb_37_45 bitb_37_46 R_bl
Cb_37_45 bit_37_45 gnd C_bl
Cbb_37_45 bitb_37_45 gnd C_bl
Rb_37_46 bit_37_46 bit_37_47 R_bl
Rbb_37_46 bitb_37_46 bitb_37_47 R_bl
Cb_37_46 bit_37_46 gnd C_bl
Cbb_37_46 bitb_37_46 gnd C_bl
Rb_37_47 bit_37_47 bit_37_48 R_bl
Rbb_37_47 bitb_37_47 bitb_37_48 R_bl
Cb_37_47 bit_37_47 gnd C_bl
Cbb_37_47 bitb_37_47 gnd C_bl
Rb_37_48 bit_37_48 bit_37_49 R_bl
Rbb_37_48 bitb_37_48 bitb_37_49 R_bl
Cb_37_48 bit_37_48 gnd C_bl
Cbb_37_48 bitb_37_48 gnd C_bl
Rb_37_49 bit_37_49 bit_37_50 R_bl
Rbb_37_49 bitb_37_49 bitb_37_50 R_bl
Cb_37_49 bit_37_49 gnd C_bl
Cbb_37_49 bitb_37_49 gnd C_bl
Rb_37_50 bit_37_50 bit_37_51 R_bl
Rbb_37_50 bitb_37_50 bitb_37_51 R_bl
Cb_37_50 bit_37_50 gnd C_bl
Cbb_37_50 bitb_37_50 gnd C_bl
Rb_37_51 bit_37_51 bit_37_52 R_bl
Rbb_37_51 bitb_37_51 bitb_37_52 R_bl
Cb_37_51 bit_37_51 gnd C_bl
Cbb_37_51 bitb_37_51 gnd C_bl
Rb_37_52 bit_37_52 bit_37_53 R_bl
Rbb_37_52 bitb_37_52 bitb_37_53 R_bl
Cb_37_52 bit_37_52 gnd C_bl
Cbb_37_52 bitb_37_52 gnd C_bl
Rb_37_53 bit_37_53 bit_37_54 R_bl
Rbb_37_53 bitb_37_53 bitb_37_54 R_bl
Cb_37_53 bit_37_53 gnd C_bl
Cbb_37_53 bitb_37_53 gnd C_bl
Rb_37_54 bit_37_54 bit_37_55 R_bl
Rbb_37_54 bitb_37_54 bitb_37_55 R_bl
Cb_37_54 bit_37_54 gnd C_bl
Cbb_37_54 bitb_37_54 gnd C_bl
Rb_37_55 bit_37_55 bit_37_56 R_bl
Rbb_37_55 bitb_37_55 bitb_37_56 R_bl
Cb_37_55 bit_37_55 gnd C_bl
Cbb_37_55 bitb_37_55 gnd C_bl
Rb_37_56 bit_37_56 bit_37_57 R_bl
Rbb_37_56 bitb_37_56 bitb_37_57 R_bl
Cb_37_56 bit_37_56 gnd C_bl
Cbb_37_56 bitb_37_56 gnd C_bl
Rb_37_57 bit_37_57 bit_37_58 R_bl
Rbb_37_57 bitb_37_57 bitb_37_58 R_bl
Cb_37_57 bit_37_57 gnd C_bl
Cbb_37_57 bitb_37_57 gnd C_bl
Rb_37_58 bit_37_58 bit_37_59 R_bl
Rbb_37_58 bitb_37_58 bitb_37_59 R_bl
Cb_37_58 bit_37_58 gnd C_bl
Cbb_37_58 bitb_37_58 gnd C_bl
Rb_37_59 bit_37_59 bit_37_60 R_bl
Rbb_37_59 bitb_37_59 bitb_37_60 R_bl
Cb_37_59 bit_37_59 gnd C_bl
Cbb_37_59 bitb_37_59 gnd C_bl
Rb_37_60 bit_37_60 bit_37_61 R_bl
Rbb_37_60 bitb_37_60 bitb_37_61 R_bl
Cb_37_60 bit_37_60 gnd C_bl
Cbb_37_60 bitb_37_60 gnd C_bl
Rb_37_61 bit_37_61 bit_37_62 R_bl
Rbb_37_61 bitb_37_61 bitb_37_62 R_bl
Cb_37_61 bit_37_61 gnd C_bl
Cbb_37_61 bitb_37_61 gnd C_bl
Rb_37_62 bit_37_62 bit_37_63 R_bl
Rbb_37_62 bitb_37_62 bitb_37_63 R_bl
Cb_37_62 bit_37_62 gnd C_bl
Cbb_37_62 bitb_37_62 gnd C_bl
Rb_37_63 bit_37_63 bit_37_64 R_bl
Rbb_37_63 bitb_37_63 bitb_37_64 R_bl
Cb_37_63 bit_37_63 gnd C_bl
Cbb_37_63 bitb_37_63 gnd C_bl
Rb_37_64 bit_37_64 bit_37_65 R_bl
Rbb_37_64 bitb_37_64 bitb_37_65 R_bl
Cb_37_64 bit_37_64 gnd C_bl
Cbb_37_64 bitb_37_64 gnd C_bl
Rb_37_65 bit_37_65 bit_37_66 R_bl
Rbb_37_65 bitb_37_65 bitb_37_66 R_bl
Cb_37_65 bit_37_65 gnd C_bl
Cbb_37_65 bitb_37_65 gnd C_bl
Rb_37_66 bit_37_66 bit_37_67 R_bl
Rbb_37_66 bitb_37_66 bitb_37_67 R_bl
Cb_37_66 bit_37_66 gnd C_bl
Cbb_37_66 bitb_37_66 gnd C_bl
Rb_37_67 bit_37_67 bit_37_68 R_bl
Rbb_37_67 bitb_37_67 bitb_37_68 R_bl
Cb_37_67 bit_37_67 gnd C_bl
Cbb_37_67 bitb_37_67 gnd C_bl
Rb_37_68 bit_37_68 bit_37_69 R_bl
Rbb_37_68 bitb_37_68 bitb_37_69 R_bl
Cb_37_68 bit_37_68 gnd C_bl
Cbb_37_68 bitb_37_68 gnd C_bl
Rb_37_69 bit_37_69 bit_37_70 R_bl
Rbb_37_69 bitb_37_69 bitb_37_70 R_bl
Cb_37_69 bit_37_69 gnd C_bl
Cbb_37_69 bitb_37_69 gnd C_bl
Rb_37_70 bit_37_70 bit_37_71 R_bl
Rbb_37_70 bitb_37_70 bitb_37_71 R_bl
Cb_37_70 bit_37_70 gnd C_bl
Cbb_37_70 bitb_37_70 gnd C_bl
Rb_37_71 bit_37_71 bit_37_72 R_bl
Rbb_37_71 bitb_37_71 bitb_37_72 R_bl
Cb_37_71 bit_37_71 gnd C_bl
Cbb_37_71 bitb_37_71 gnd C_bl
Rb_37_72 bit_37_72 bit_37_73 R_bl
Rbb_37_72 bitb_37_72 bitb_37_73 R_bl
Cb_37_72 bit_37_72 gnd C_bl
Cbb_37_72 bitb_37_72 gnd C_bl
Rb_37_73 bit_37_73 bit_37_74 R_bl
Rbb_37_73 bitb_37_73 bitb_37_74 R_bl
Cb_37_73 bit_37_73 gnd C_bl
Cbb_37_73 bitb_37_73 gnd C_bl
Rb_37_74 bit_37_74 bit_37_75 R_bl
Rbb_37_74 bitb_37_74 bitb_37_75 R_bl
Cb_37_74 bit_37_74 gnd C_bl
Cbb_37_74 bitb_37_74 gnd C_bl
Rb_37_75 bit_37_75 bit_37_76 R_bl
Rbb_37_75 bitb_37_75 bitb_37_76 R_bl
Cb_37_75 bit_37_75 gnd C_bl
Cbb_37_75 bitb_37_75 gnd C_bl
Rb_37_76 bit_37_76 bit_37_77 R_bl
Rbb_37_76 bitb_37_76 bitb_37_77 R_bl
Cb_37_76 bit_37_76 gnd C_bl
Cbb_37_76 bitb_37_76 gnd C_bl
Rb_37_77 bit_37_77 bit_37_78 R_bl
Rbb_37_77 bitb_37_77 bitb_37_78 R_bl
Cb_37_77 bit_37_77 gnd C_bl
Cbb_37_77 bitb_37_77 gnd C_bl
Rb_37_78 bit_37_78 bit_37_79 R_bl
Rbb_37_78 bitb_37_78 bitb_37_79 R_bl
Cb_37_78 bit_37_78 gnd C_bl
Cbb_37_78 bitb_37_78 gnd C_bl
Rb_37_79 bit_37_79 bit_37_80 R_bl
Rbb_37_79 bitb_37_79 bitb_37_80 R_bl
Cb_37_79 bit_37_79 gnd C_bl
Cbb_37_79 bitb_37_79 gnd C_bl
Rb_37_80 bit_37_80 bit_37_81 R_bl
Rbb_37_80 bitb_37_80 bitb_37_81 R_bl
Cb_37_80 bit_37_80 gnd C_bl
Cbb_37_80 bitb_37_80 gnd C_bl
Rb_37_81 bit_37_81 bit_37_82 R_bl
Rbb_37_81 bitb_37_81 bitb_37_82 R_bl
Cb_37_81 bit_37_81 gnd C_bl
Cbb_37_81 bitb_37_81 gnd C_bl
Rb_37_82 bit_37_82 bit_37_83 R_bl
Rbb_37_82 bitb_37_82 bitb_37_83 R_bl
Cb_37_82 bit_37_82 gnd C_bl
Cbb_37_82 bitb_37_82 gnd C_bl
Rb_37_83 bit_37_83 bit_37_84 R_bl
Rbb_37_83 bitb_37_83 bitb_37_84 R_bl
Cb_37_83 bit_37_83 gnd C_bl
Cbb_37_83 bitb_37_83 gnd C_bl
Rb_37_84 bit_37_84 bit_37_85 R_bl
Rbb_37_84 bitb_37_84 bitb_37_85 R_bl
Cb_37_84 bit_37_84 gnd C_bl
Cbb_37_84 bitb_37_84 gnd C_bl
Rb_37_85 bit_37_85 bit_37_86 R_bl
Rbb_37_85 bitb_37_85 bitb_37_86 R_bl
Cb_37_85 bit_37_85 gnd C_bl
Cbb_37_85 bitb_37_85 gnd C_bl
Rb_37_86 bit_37_86 bit_37_87 R_bl
Rbb_37_86 bitb_37_86 bitb_37_87 R_bl
Cb_37_86 bit_37_86 gnd C_bl
Cbb_37_86 bitb_37_86 gnd C_bl
Rb_37_87 bit_37_87 bit_37_88 R_bl
Rbb_37_87 bitb_37_87 bitb_37_88 R_bl
Cb_37_87 bit_37_87 gnd C_bl
Cbb_37_87 bitb_37_87 gnd C_bl
Rb_37_88 bit_37_88 bit_37_89 R_bl
Rbb_37_88 bitb_37_88 bitb_37_89 R_bl
Cb_37_88 bit_37_88 gnd C_bl
Cbb_37_88 bitb_37_88 gnd C_bl
Rb_37_89 bit_37_89 bit_37_90 R_bl
Rbb_37_89 bitb_37_89 bitb_37_90 R_bl
Cb_37_89 bit_37_89 gnd C_bl
Cbb_37_89 bitb_37_89 gnd C_bl
Rb_37_90 bit_37_90 bit_37_91 R_bl
Rbb_37_90 bitb_37_90 bitb_37_91 R_bl
Cb_37_90 bit_37_90 gnd C_bl
Cbb_37_90 bitb_37_90 gnd C_bl
Rb_37_91 bit_37_91 bit_37_92 R_bl
Rbb_37_91 bitb_37_91 bitb_37_92 R_bl
Cb_37_91 bit_37_91 gnd C_bl
Cbb_37_91 bitb_37_91 gnd C_bl
Rb_37_92 bit_37_92 bit_37_93 R_bl
Rbb_37_92 bitb_37_92 bitb_37_93 R_bl
Cb_37_92 bit_37_92 gnd C_bl
Cbb_37_92 bitb_37_92 gnd C_bl
Rb_37_93 bit_37_93 bit_37_94 R_bl
Rbb_37_93 bitb_37_93 bitb_37_94 R_bl
Cb_37_93 bit_37_93 gnd C_bl
Cbb_37_93 bitb_37_93 gnd C_bl
Rb_37_94 bit_37_94 bit_37_95 R_bl
Rbb_37_94 bitb_37_94 bitb_37_95 R_bl
Cb_37_94 bit_37_94 gnd C_bl
Cbb_37_94 bitb_37_94 gnd C_bl
Rb_37_95 bit_37_95 bit_37_96 R_bl
Rbb_37_95 bitb_37_95 bitb_37_96 R_bl
Cb_37_95 bit_37_95 gnd C_bl
Cbb_37_95 bitb_37_95 gnd C_bl
Rb_37_96 bit_37_96 bit_37_97 R_bl
Rbb_37_96 bitb_37_96 bitb_37_97 R_bl
Cb_37_96 bit_37_96 gnd C_bl
Cbb_37_96 bitb_37_96 gnd C_bl
Rb_37_97 bit_37_97 bit_37_98 R_bl
Rbb_37_97 bitb_37_97 bitb_37_98 R_bl
Cb_37_97 bit_37_97 gnd C_bl
Cbb_37_97 bitb_37_97 gnd C_bl
Rb_37_98 bit_37_98 bit_37_99 R_bl
Rbb_37_98 bitb_37_98 bitb_37_99 R_bl
Cb_37_98 bit_37_98 gnd C_bl
Cbb_37_98 bitb_37_98 gnd C_bl
Rb_37_99 bit_37_99 bit_37_100 R_bl
Rbb_37_99 bitb_37_99 bitb_37_100 R_bl
Cb_37_99 bit_37_99 gnd C_bl
Cbb_37_99 bitb_37_99 gnd C_bl
Rb_38_0 bit_38_0 bit_38_1 R_bl
Rbb_38_0 bitb_38_0 bitb_38_1 R_bl
Cb_38_0 bit_38_0 gnd C_bl
Cbb_38_0 bitb_38_0 gnd C_bl
Rb_38_1 bit_38_1 bit_38_2 R_bl
Rbb_38_1 bitb_38_1 bitb_38_2 R_bl
Cb_38_1 bit_38_1 gnd C_bl
Cbb_38_1 bitb_38_1 gnd C_bl
Rb_38_2 bit_38_2 bit_38_3 R_bl
Rbb_38_2 bitb_38_2 bitb_38_3 R_bl
Cb_38_2 bit_38_2 gnd C_bl
Cbb_38_2 bitb_38_2 gnd C_bl
Rb_38_3 bit_38_3 bit_38_4 R_bl
Rbb_38_3 bitb_38_3 bitb_38_4 R_bl
Cb_38_3 bit_38_3 gnd C_bl
Cbb_38_3 bitb_38_3 gnd C_bl
Rb_38_4 bit_38_4 bit_38_5 R_bl
Rbb_38_4 bitb_38_4 bitb_38_5 R_bl
Cb_38_4 bit_38_4 gnd C_bl
Cbb_38_4 bitb_38_4 gnd C_bl
Rb_38_5 bit_38_5 bit_38_6 R_bl
Rbb_38_5 bitb_38_5 bitb_38_6 R_bl
Cb_38_5 bit_38_5 gnd C_bl
Cbb_38_5 bitb_38_5 gnd C_bl
Rb_38_6 bit_38_6 bit_38_7 R_bl
Rbb_38_6 bitb_38_6 bitb_38_7 R_bl
Cb_38_6 bit_38_6 gnd C_bl
Cbb_38_6 bitb_38_6 gnd C_bl
Rb_38_7 bit_38_7 bit_38_8 R_bl
Rbb_38_7 bitb_38_7 bitb_38_8 R_bl
Cb_38_7 bit_38_7 gnd C_bl
Cbb_38_7 bitb_38_7 gnd C_bl
Rb_38_8 bit_38_8 bit_38_9 R_bl
Rbb_38_8 bitb_38_8 bitb_38_9 R_bl
Cb_38_8 bit_38_8 gnd C_bl
Cbb_38_8 bitb_38_8 gnd C_bl
Rb_38_9 bit_38_9 bit_38_10 R_bl
Rbb_38_9 bitb_38_9 bitb_38_10 R_bl
Cb_38_9 bit_38_9 gnd C_bl
Cbb_38_9 bitb_38_9 gnd C_bl
Rb_38_10 bit_38_10 bit_38_11 R_bl
Rbb_38_10 bitb_38_10 bitb_38_11 R_bl
Cb_38_10 bit_38_10 gnd C_bl
Cbb_38_10 bitb_38_10 gnd C_bl
Rb_38_11 bit_38_11 bit_38_12 R_bl
Rbb_38_11 bitb_38_11 bitb_38_12 R_bl
Cb_38_11 bit_38_11 gnd C_bl
Cbb_38_11 bitb_38_11 gnd C_bl
Rb_38_12 bit_38_12 bit_38_13 R_bl
Rbb_38_12 bitb_38_12 bitb_38_13 R_bl
Cb_38_12 bit_38_12 gnd C_bl
Cbb_38_12 bitb_38_12 gnd C_bl
Rb_38_13 bit_38_13 bit_38_14 R_bl
Rbb_38_13 bitb_38_13 bitb_38_14 R_bl
Cb_38_13 bit_38_13 gnd C_bl
Cbb_38_13 bitb_38_13 gnd C_bl
Rb_38_14 bit_38_14 bit_38_15 R_bl
Rbb_38_14 bitb_38_14 bitb_38_15 R_bl
Cb_38_14 bit_38_14 gnd C_bl
Cbb_38_14 bitb_38_14 gnd C_bl
Rb_38_15 bit_38_15 bit_38_16 R_bl
Rbb_38_15 bitb_38_15 bitb_38_16 R_bl
Cb_38_15 bit_38_15 gnd C_bl
Cbb_38_15 bitb_38_15 gnd C_bl
Rb_38_16 bit_38_16 bit_38_17 R_bl
Rbb_38_16 bitb_38_16 bitb_38_17 R_bl
Cb_38_16 bit_38_16 gnd C_bl
Cbb_38_16 bitb_38_16 gnd C_bl
Rb_38_17 bit_38_17 bit_38_18 R_bl
Rbb_38_17 bitb_38_17 bitb_38_18 R_bl
Cb_38_17 bit_38_17 gnd C_bl
Cbb_38_17 bitb_38_17 gnd C_bl
Rb_38_18 bit_38_18 bit_38_19 R_bl
Rbb_38_18 bitb_38_18 bitb_38_19 R_bl
Cb_38_18 bit_38_18 gnd C_bl
Cbb_38_18 bitb_38_18 gnd C_bl
Rb_38_19 bit_38_19 bit_38_20 R_bl
Rbb_38_19 bitb_38_19 bitb_38_20 R_bl
Cb_38_19 bit_38_19 gnd C_bl
Cbb_38_19 bitb_38_19 gnd C_bl
Rb_38_20 bit_38_20 bit_38_21 R_bl
Rbb_38_20 bitb_38_20 bitb_38_21 R_bl
Cb_38_20 bit_38_20 gnd C_bl
Cbb_38_20 bitb_38_20 gnd C_bl
Rb_38_21 bit_38_21 bit_38_22 R_bl
Rbb_38_21 bitb_38_21 bitb_38_22 R_bl
Cb_38_21 bit_38_21 gnd C_bl
Cbb_38_21 bitb_38_21 gnd C_bl
Rb_38_22 bit_38_22 bit_38_23 R_bl
Rbb_38_22 bitb_38_22 bitb_38_23 R_bl
Cb_38_22 bit_38_22 gnd C_bl
Cbb_38_22 bitb_38_22 gnd C_bl
Rb_38_23 bit_38_23 bit_38_24 R_bl
Rbb_38_23 bitb_38_23 bitb_38_24 R_bl
Cb_38_23 bit_38_23 gnd C_bl
Cbb_38_23 bitb_38_23 gnd C_bl
Rb_38_24 bit_38_24 bit_38_25 R_bl
Rbb_38_24 bitb_38_24 bitb_38_25 R_bl
Cb_38_24 bit_38_24 gnd C_bl
Cbb_38_24 bitb_38_24 gnd C_bl
Rb_38_25 bit_38_25 bit_38_26 R_bl
Rbb_38_25 bitb_38_25 bitb_38_26 R_bl
Cb_38_25 bit_38_25 gnd C_bl
Cbb_38_25 bitb_38_25 gnd C_bl
Rb_38_26 bit_38_26 bit_38_27 R_bl
Rbb_38_26 bitb_38_26 bitb_38_27 R_bl
Cb_38_26 bit_38_26 gnd C_bl
Cbb_38_26 bitb_38_26 gnd C_bl
Rb_38_27 bit_38_27 bit_38_28 R_bl
Rbb_38_27 bitb_38_27 bitb_38_28 R_bl
Cb_38_27 bit_38_27 gnd C_bl
Cbb_38_27 bitb_38_27 gnd C_bl
Rb_38_28 bit_38_28 bit_38_29 R_bl
Rbb_38_28 bitb_38_28 bitb_38_29 R_bl
Cb_38_28 bit_38_28 gnd C_bl
Cbb_38_28 bitb_38_28 gnd C_bl
Rb_38_29 bit_38_29 bit_38_30 R_bl
Rbb_38_29 bitb_38_29 bitb_38_30 R_bl
Cb_38_29 bit_38_29 gnd C_bl
Cbb_38_29 bitb_38_29 gnd C_bl
Rb_38_30 bit_38_30 bit_38_31 R_bl
Rbb_38_30 bitb_38_30 bitb_38_31 R_bl
Cb_38_30 bit_38_30 gnd C_bl
Cbb_38_30 bitb_38_30 gnd C_bl
Rb_38_31 bit_38_31 bit_38_32 R_bl
Rbb_38_31 bitb_38_31 bitb_38_32 R_bl
Cb_38_31 bit_38_31 gnd C_bl
Cbb_38_31 bitb_38_31 gnd C_bl
Rb_38_32 bit_38_32 bit_38_33 R_bl
Rbb_38_32 bitb_38_32 bitb_38_33 R_bl
Cb_38_32 bit_38_32 gnd C_bl
Cbb_38_32 bitb_38_32 gnd C_bl
Rb_38_33 bit_38_33 bit_38_34 R_bl
Rbb_38_33 bitb_38_33 bitb_38_34 R_bl
Cb_38_33 bit_38_33 gnd C_bl
Cbb_38_33 bitb_38_33 gnd C_bl
Rb_38_34 bit_38_34 bit_38_35 R_bl
Rbb_38_34 bitb_38_34 bitb_38_35 R_bl
Cb_38_34 bit_38_34 gnd C_bl
Cbb_38_34 bitb_38_34 gnd C_bl
Rb_38_35 bit_38_35 bit_38_36 R_bl
Rbb_38_35 bitb_38_35 bitb_38_36 R_bl
Cb_38_35 bit_38_35 gnd C_bl
Cbb_38_35 bitb_38_35 gnd C_bl
Rb_38_36 bit_38_36 bit_38_37 R_bl
Rbb_38_36 bitb_38_36 bitb_38_37 R_bl
Cb_38_36 bit_38_36 gnd C_bl
Cbb_38_36 bitb_38_36 gnd C_bl
Rb_38_37 bit_38_37 bit_38_38 R_bl
Rbb_38_37 bitb_38_37 bitb_38_38 R_bl
Cb_38_37 bit_38_37 gnd C_bl
Cbb_38_37 bitb_38_37 gnd C_bl
Rb_38_38 bit_38_38 bit_38_39 R_bl
Rbb_38_38 bitb_38_38 bitb_38_39 R_bl
Cb_38_38 bit_38_38 gnd C_bl
Cbb_38_38 bitb_38_38 gnd C_bl
Rb_38_39 bit_38_39 bit_38_40 R_bl
Rbb_38_39 bitb_38_39 bitb_38_40 R_bl
Cb_38_39 bit_38_39 gnd C_bl
Cbb_38_39 bitb_38_39 gnd C_bl
Rb_38_40 bit_38_40 bit_38_41 R_bl
Rbb_38_40 bitb_38_40 bitb_38_41 R_bl
Cb_38_40 bit_38_40 gnd C_bl
Cbb_38_40 bitb_38_40 gnd C_bl
Rb_38_41 bit_38_41 bit_38_42 R_bl
Rbb_38_41 bitb_38_41 bitb_38_42 R_bl
Cb_38_41 bit_38_41 gnd C_bl
Cbb_38_41 bitb_38_41 gnd C_bl
Rb_38_42 bit_38_42 bit_38_43 R_bl
Rbb_38_42 bitb_38_42 bitb_38_43 R_bl
Cb_38_42 bit_38_42 gnd C_bl
Cbb_38_42 bitb_38_42 gnd C_bl
Rb_38_43 bit_38_43 bit_38_44 R_bl
Rbb_38_43 bitb_38_43 bitb_38_44 R_bl
Cb_38_43 bit_38_43 gnd C_bl
Cbb_38_43 bitb_38_43 gnd C_bl
Rb_38_44 bit_38_44 bit_38_45 R_bl
Rbb_38_44 bitb_38_44 bitb_38_45 R_bl
Cb_38_44 bit_38_44 gnd C_bl
Cbb_38_44 bitb_38_44 gnd C_bl
Rb_38_45 bit_38_45 bit_38_46 R_bl
Rbb_38_45 bitb_38_45 bitb_38_46 R_bl
Cb_38_45 bit_38_45 gnd C_bl
Cbb_38_45 bitb_38_45 gnd C_bl
Rb_38_46 bit_38_46 bit_38_47 R_bl
Rbb_38_46 bitb_38_46 bitb_38_47 R_bl
Cb_38_46 bit_38_46 gnd C_bl
Cbb_38_46 bitb_38_46 gnd C_bl
Rb_38_47 bit_38_47 bit_38_48 R_bl
Rbb_38_47 bitb_38_47 bitb_38_48 R_bl
Cb_38_47 bit_38_47 gnd C_bl
Cbb_38_47 bitb_38_47 gnd C_bl
Rb_38_48 bit_38_48 bit_38_49 R_bl
Rbb_38_48 bitb_38_48 bitb_38_49 R_bl
Cb_38_48 bit_38_48 gnd C_bl
Cbb_38_48 bitb_38_48 gnd C_bl
Rb_38_49 bit_38_49 bit_38_50 R_bl
Rbb_38_49 bitb_38_49 bitb_38_50 R_bl
Cb_38_49 bit_38_49 gnd C_bl
Cbb_38_49 bitb_38_49 gnd C_bl
Rb_38_50 bit_38_50 bit_38_51 R_bl
Rbb_38_50 bitb_38_50 bitb_38_51 R_bl
Cb_38_50 bit_38_50 gnd C_bl
Cbb_38_50 bitb_38_50 gnd C_bl
Rb_38_51 bit_38_51 bit_38_52 R_bl
Rbb_38_51 bitb_38_51 bitb_38_52 R_bl
Cb_38_51 bit_38_51 gnd C_bl
Cbb_38_51 bitb_38_51 gnd C_bl
Rb_38_52 bit_38_52 bit_38_53 R_bl
Rbb_38_52 bitb_38_52 bitb_38_53 R_bl
Cb_38_52 bit_38_52 gnd C_bl
Cbb_38_52 bitb_38_52 gnd C_bl
Rb_38_53 bit_38_53 bit_38_54 R_bl
Rbb_38_53 bitb_38_53 bitb_38_54 R_bl
Cb_38_53 bit_38_53 gnd C_bl
Cbb_38_53 bitb_38_53 gnd C_bl
Rb_38_54 bit_38_54 bit_38_55 R_bl
Rbb_38_54 bitb_38_54 bitb_38_55 R_bl
Cb_38_54 bit_38_54 gnd C_bl
Cbb_38_54 bitb_38_54 gnd C_bl
Rb_38_55 bit_38_55 bit_38_56 R_bl
Rbb_38_55 bitb_38_55 bitb_38_56 R_bl
Cb_38_55 bit_38_55 gnd C_bl
Cbb_38_55 bitb_38_55 gnd C_bl
Rb_38_56 bit_38_56 bit_38_57 R_bl
Rbb_38_56 bitb_38_56 bitb_38_57 R_bl
Cb_38_56 bit_38_56 gnd C_bl
Cbb_38_56 bitb_38_56 gnd C_bl
Rb_38_57 bit_38_57 bit_38_58 R_bl
Rbb_38_57 bitb_38_57 bitb_38_58 R_bl
Cb_38_57 bit_38_57 gnd C_bl
Cbb_38_57 bitb_38_57 gnd C_bl
Rb_38_58 bit_38_58 bit_38_59 R_bl
Rbb_38_58 bitb_38_58 bitb_38_59 R_bl
Cb_38_58 bit_38_58 gnd C_bl
Cbb_38_58 bitb_38_58 gnd C_bl
Rb_38_59 bit_38_59 bit_38_60 R_bl
Rbb_38_59 bitb_38_59 bitb_38_60 R_bl
Cb_38_59 bit_38_59 gnd C_bl
Cbb_38_59 bitb_38_59 gnd C_bl
Rb_38_60 bit_38_60 bit_38_61 R_bl
Rbb_38_60 bitb_38_60 bitb_38_61 R_bl
Cb_38_60 bit_38_60 gnd C_bl
Cbb_38_60 bitb_38_60 gnd C_bl
Rb_38_61 bit_38_61 bit_38_62 R_bl
Rbb_38_61 bitb_38_61 bitb_38_62 R_bl
Cb_38_61 bit_38_61 gnd C_bl
Cbb_38_61 bitb_38_61 gnd C_bl
Rb_38_62 bit_38_62 bit_38_63 R_bl
Rbb_38_62 bitb_38_62 bitb_38_63 R_bl
Cb_38_62 bit_38_62 gnd C_bl
Cbb_38_62 bitb_38_62 gnd C_bl
Rb_38_63 bit_38_63 bit_38_64 R_bl
Rbb_38_63 bitb_38_63 bitb_38_64 R_bl
Cb_38_63 bit_38_63 gnd C_bl
Cbb_38_63 bitb_38_63 gnd C_bl
Rb_38_64 bit_38_64 bit_38_65 R_bl
Rbb_38_64 bitb_38_64 bitb_38_65 R_bl
Cb_38_64 bit_38_64 gnd C_bl
Cbb_38_64 bitb_38_64 gnd C_bl
Rb_38_65 bit_38_65 bit_38_66 R_bl
Rbb_38_65 bitb_38_65 bitb_38_66 R_bl
Cb_38_65 bit_38_65 gnd C_bl
Cbb_38_65 bitb_38_65 gnd C_bl
Rb_38_66 bit_38_66 bit_38_67 R_bl
Rbb_38_66 bitb_38_66 bitb_38_67 R_bl
Cb_38_66 bit_38_66 gnd C_bl
Cbb_38_66 bitb_38_66 gnd C_bl
Rb_38_67 bit_38_67 bit_38_68 R_bl
Rbb_38_67 bitb_38_67 bitb_38_68 R_bl
Cb_38_67 bit_38_67 gnd C_bl
Cbb_38_67 bitb_38_67 gnd C_bl
Rb_38_68 bit_38_68 bit_38_69 R_bl
Rbb_38_68 bitb_38_68 bitb_38_69 R_bl
Cb_38_68 bit_38_68 gnd C_bl
Cbb_38_68 bitb_38_68 gnd C_bl
Rb_38_69 bit_38_69 bit_38_70 R_bl
Rbb_38_69 bitb_38_69 bitb_38_70 R_bl
Cb_38_69 bit_38_69 gnd C_bl
Cbb_38_69 bitb_38_69 gnd C_bl
Rb_38_70 bit_38_70 bit_38_71 R_bl
Rbb_38_70 bitb_38_70 bitb_38_71 R_bl
Cb_38_70 bit_38_70 gnd C_bl
Cbb_38_70 bitb_38_70 gnd C_bl
Rb_38_71 bit_38_71 bit_38_72 R_bl
Rbb_38_71 bitb_38_71 bitb_38_72 R_bl
Cb_38_71 bit_38_71 gnd C_bl
Cbb_38_71 bitb_38_71 gnd C_bl
Rb_38_72 bit_38_72 bit_38_73 R_bl
Rbb_38_72 bitb_38_72 bitb_38_73 R_bl
Cb_38_72 bit_38_72 gnd C_bl
Cbb_38_72 bitb_38_72 gnd C_bl
Rb_38_73 bit_38_73 bit_38_74 R_bl
Rbb_38_73 bitb_38_73 bitb_38_74 R_bl
Cb_38_73 bit_38_73 gnd C_bl
Cbb_38_73 bitb_38_73 gnd C_bl
Rb_38_74 bit_38_74 bit_38_75 R_bl
Rbb_38_74 bitb_38_74 bitb_38_75 R_bl
Cb_38_74 bit_38_74 gnd C_bl
Cbb_38_74 bitb_38_74 gnd C_bl
Rb_38_75 bit_38_75 bit_38_76 R_bl
Rbb_38_75 bitb_38_75 bitb_38_76 R_bl
Cb_38_75 bit_38_75 gnd C_bl
Cbb_38_75 bitb_38_75 gnd C_bl
Rb_38_76 bit_38_76 bit_38_77 R_bl
Rbb_38_76 bitb_38_76 bitb_38_77 R_bl
Cb_38_76 bit_38_76 gnd C_bl
Cbb_38_76 bitb_38_76 gnd C_bl
Rb_38_77 bit_38_77 bit_38_78 R_bl
Rbb_38_77 bitb_38_77 bitb_38_78 R_bl
Cb_38_77 bit_38_77 gnd C_bl
Cbb_38_77 bitb_38_77 gnd C_bl
Rb_38_78 bit_38_78 bit_38_79 R_bl
Rbb_38_78 bitb_38_78 bitb_38_79 R_bl
Cb_38_78 bit_38_78 gnd C_bl
Cbb_38_78 bitb_38_78 gnd C_bl
Rb_38_79 bit_38_79 bit_38_80 R_bl
Rbb_38_79 bitb_38_79 bitb_38_80 R_bl
Cb_38_79 bit_38_79 gnd C_bl
Cbb_38_79 bitb_38_79 gnd C_bl
Rb_38_80 bit_38_80 bit_38_81 R_bl
Rbb_38_80 bitb_38_80 bitb_38_81 R_bl
Cb_38_80 bit_38_80 gnd C_bl
Cbb_38_80 bitb_38_80 gnd C_bl
Rb_38_81 bit_38_81 bit_38_82 R_bl
Rbb_38_81 bitb_38_81 bitb_38_82 R_bl
Cb_38_81 bit_38_81 gnd C_bl
Cbb_38_81 bitb_38_81 gnd C_bl
Rb_38_82 bit_38_82 bit_38_83 R_bl
Rbb_38_82 bitb_38_82 bitb_38_83 R_bl
Cb_38_82 bit_38_82 gnd C_bl
Cbb_38_82 bitb_38_82 gnd C_bl
Rb_38_83 bit_38_83 bit_38_84 R_bl
Rbb_38_83 bitb_38_83 bitb_38_84 R_bl
Cb_38_83 bit_38_83 gnd C_bl
Cbb_38_83 bitb_38_83 gnd C_bl
Rb_38_84 bit_38_84 bit_38_85 R_bl
Rbb_38_84 bitb_38_84 bitb_38_85 R_bl
Cb_38_84 bit_38_84 gnd C_bl
Cbb_38_84 bitb_38_84 gnd C_bl
Rb_38_85 bit_38_85 bit_38_86 R_bl
Rbb_38_85 bitb_38_85 bitb_38_86 R_bl
Cb_38_85 bit_38_85 gnd C_bl
Cbb_38_85 bitb_38_85 gnd C_bl
Rb_38_86 bit_38_86 bit_38_87 R_bl
Rbb_38_86 bitb_38_86 bitb_38_87 R_bl
Cb_38_86 bit_38_86 gnd C_bl
Cbb_38_86 bitb_38_86 gnd C_bl
Rb_38_87 bit_38_87 bit_38_88 R_bl
Rbb_38_87 bitb_38_87 bitb_38_88 R_bl
Cb_38_87 bit_38_87 gnd C_bl
Cbb_38_87 bitb_38_87 gnd C_bl
Rb_38_88 bit_38_88 bit_38_89 R_bl
Rbb_38_88 bitb_38_88 bitb_38_89 R_bl
Cb_38_88 bit_38_88 gnd C_bl
Cbb_38_88 bitb_38_88 gnd C_bl
Rb_38_89 bit_38_89 bit_38_90 R_bl
Rbb_38_89 bitb_38_89 bitb_38_90 R_bl
Cb_38_89 bit_38_89 gnd C_bl
Cbb_38_89 bitb_38_89 gnd C_bl
Rb_38_90 bit_38_90 bit_38_91 R_bl
Rbb_38_90 bitb_38_90 bitb_38_91 R_bl
Cb_38_90 bit_38_90 gnd C_bl
Cbb_38_90 bitb_38_90 gnd C_bl
Rb_38_91 bit_38_91 bit_38_92 R_bl
Rbb_38_91 bitb_38_91 bitb_38_92 R_bl
Cb_38_91 bit_38_91 gnd C_bl
Cbb_38_91 bitb_38_91 gnd C_bl
Rb_38_92 bit_38_92 bit_38_93 R_bl
Rbb_38_92 bitb_38_92 bitb_38_93 R_bl
Cb_38_92 bit_38_92 gnd C_bl
Cbb_38_92 bitb_38_92 gnd C_bl
Rb_38_93 bit_38_93 bit_38_94 R_bl
Rbb_38_93 bitb_38_93 bitb_38_94 R_bl
Cb_38_93 bit_38_93 gnd C_bl
Cbb_38_93 bitb_38_93 gnd C_bl
Rb_38_94 bit_38_94 bit_38_95 R_bl
Rbb_38_94 bitb_38_94 bitb_38_95 R_bl
Cb_38_94 bit_38_94 gnd C_bl
Cbb_38_94 bitb_38_94 gnd C_bl
Rb_38_95 bit_38_95 bit_38_96 R_bl
Rbb_38_95 bitb_38_95 bitb_38_96 R_bl
Cb_38_95 bit_38_95 gnd C_bl
Cbb_38_95 bitb_38_95 gnd C_bl
Rb_38_96 bit_38_96 bit_38_97 R_bl
Rbb_38_96 bitb_38_96 bitb_38_97 R_bl
Cb_38_96 bit_38_96 gnd C_bl
Cbb_38_96 bitb_38_96 gnd C_bl
Rb_38_97 bit_38_97 bit_38_98 R_bl
Rbb_38_97 bitb_38_97 bitb_38_98 R_bl
Cb_38_97 bit_38_97 gnd C_bl
Cbb_38_97 bitb_38_97 gnd C_bl
Rb_38_98 bit_38_98 bit_38_99 R_bl
Rbb_38_98 bitb_38_98 bitb_38_99 R_bl
Cb_38_98 bit_38_98 gnd C_bl
Cbb_38_98 bitb_38_98 gnd C_bl
Rb_38_99 bit_38_99 bit_38_100 R_bl
Rbb_38_99 bitb_38_99 bitb_38_100 R_bl
Cb_38_99 bit_38_99 gnd C_bl
Cbb_38_99 bitb_38_99 gnd C_bl
Rb_39_0 bit_39_0 bit_39_1 R_bl
Rbb_39_0 bitb_39_0 bitb_39_1 R_bl
Cb_39_0 bit_39_0 gnd C_bl
Cbb_39_0 bitb_39_0 gnd C_bl
Rb_39_1 bit_39_1 bit_39_2 R_bl
Rbb_39_1 bitb_39_1 bitb_39_2 R_bl
Cb_39_1 bit_39_1 gnd C_bl
Cbb_39_1 bitb_39_1 gnd C_bl
Rb_39_2 bit_39_2 bit_39_3 R_bl
Rbb_39_2 bitb_39_2 bitb_39_3 R_bl
Cb_39_2 bit_39_2 gnd C_bl
Cbb_39_2 bitb_39_2 gnd C_bl
Rb_39_3 bit_39_3 bit_39_4 R_bl
Rbb_39_3 bitb_39_3 bitb_39_4 R_bl
Cb_39_3 bit_39_3 gnd C_bl
Cbb_39_3 bitb_39_3 gnd C_bl
Rb_39_4 bit_39_4 bit_39_5 R_bl
Rbb_39_4 bitb_39_4 bitb_39_5 R_bl
Cb_39_4 bit_39_4 gnd C_bl
Cbb_39_4 bitb_39_4 gnd C_bl
Rb_39_5 bit_39_5 bit_39_6 R_bl
Rbb_39_5 bitb_39_5 bitb_39_6 R_bl
Cb_39_5 bit_39_5 gnd C_bl
Cbb_39_5 bitb_39_5 gnd C_bl
Rb_39_6 bit_39_6 bit_39_7 R_bl
Rbb_39_6 bitb_39_6 bitb_39_7 R_bl
Cb_39_6 bit_39_6 gnd C_bl
Cbb_39_6 bitb_39_6 gnd C_bl
Rb_39_7 bit_39_7 bit_39_8 R_bl
Rbb_39_7 bitb_39_7 bitb_39_8 R_bl
Cb_39_7 bit_39_7 gnd C_bl
Cbb_39_7 bitb_39_7 gnd C_bl
Rb_39_8 bit_39_8 bit_39_9 R_bl
Rbb_39_8 bitb_39_8 bitb_39_9 R_bl
Cb_39_8 bit_39_8 gnd C_bl
Cbb_39_8 bitb_39_8 gnd C_bl
Rb_39_9 bit_39_9 bit_39_10 R_bl
Rbb_39_9 bitb_39_9 bitb_39_10 R_bl
Cb_39_9 bit_39_9 gnd C_bl
Cbb_39_9 bitb_39_9 gnd C_bl
Rb_39_10 bit_39_10 bit_39_11 R_bl
Rbb_39_10 bitb_39_10 bitb_39_11 R_bl
Cb_39_10 bit_39_10 gnd C_bl
Cbb_39_10 bitb_39_10 gnd C_bl
Rb_39_11 bit_39_11 bit_39_12 R_bl
Rbb_39_11 bitb_39_11 bitb_39_12 R_bl
Cb_39_11 bit_39_11 gnd C_bl
Cbb_39_11 bitb_39_11 gnd C_bl
Rb_39_12 bit_39_12 bit_39_13 R_bl
Rbb_39_12 bitb_39_12 bitb_39_13 R_bl
Cb_39_12 bit_39_12 gnd C_bl
Cbb_39_12 bitb_39_12 gnd C_bl
Rb_39_13 bit_39_13 bit_39_14 R_bl
Rbb_39_13 bitb_39_13 bitb_39_14 R_bl
Cb_39_13 bit_39_13 gnd C_bl
Cbb_39_13 bitb_39_13 gnd C_bl
Rb_39_14 bit_39_14 bit_39_15 R_bl
Rbb_39_14 bitb_39_14 bitb_39_15 R_bl
Cb_39_14 bit_39_14 gnd C_bl
Cbb_39_14 bitb_39_14 gnd C_bl
Rb_39_15 bit_39_15 bit_39_16 R_bl
Rbb_39_15 bitb_39_15 bitb_39_16 R_bl
Cb_39_15 bit_39_15 gnd C_bl
Cbb_39_15 bitb_39_15 gnd C_bl
Rb_39_16 bit_39_16 bit_39_17 R_bl
Rbb_39_16 bitb_39_16 bitb_39_17 R_bl
Cb_39_16 bit_39_16 gnd C_bl
Cbb_39_16 bitb_39_16 gnd C_bl
Rb_39_17 bit_39_17 bit_39_18 R_bl
Rbb_39_17 bitb_39_17 bitb_39_18 R_bl
Cb_39_17 bit_39_17 gnd C_bl
Cbb_39_17 bitb_39_17 gnd C_bl
Rb_39_18 bit_39_18 bit_39_19 R_bl
Rbb_39_18 bitb_39_18 bitb_39_19 R_bl
Cb_39_18 bit_39_18 gnd C_bl
Cbb_39_18 bitb_39_18 gnd C_bl
Rb_39_19 bit_39_19 bit_39_20 R_bl
Rbb_39_19 bitb_39_19 bitb_39_20 R_bl
Cb_39_19 bit_39_19 gnd C_bl
Cbb_39_19 bitb_39_19 gnd C_bl
Rb_39_20 bit_39_20 bit_39_21 R_bl
Rbb_39_20 bitb_39_20 bitb_39_21 R_bl
Cb_39_20 bit_39_20 gnd C_bl
Cbb_39_20 bitb_39_20 gnd C_bl
Rb_39_21 bit_39_21 bit_39_22 R_bl
Rbb_39_21 bitb_39_21 bitb_39_22 R_bl
Cb_39_21 bit_39_21 gnd C_bl
Cbb_39_21 bitb_39_21 gnd C_bl
Rb_39_22 bit_39_22 bit_39_23 R_bl
Rbb_39_22 bitb_39_22 bitb_39_23 R_bl
Cb_39_22 bit_39_22 gnd C_bl
Cbb_39_22 bitb_39_22 gnd C_bl
Rb_39_23 bit_39_23 bit_39_24 R_bl
Rbb_39_23 bitb_39_23 bitb_39_24 R_bl
Cb_39_23 bit_39_23 gnd C_bl
Cbb_39_23 bitb_39_23 gnd C_bl
Rb_39_24 bit_39_24 bit_39_25 R_bl
Rbb_39_24 bitb_39_24 bitb_39_25 R_bl
Cb_39_24 bit_39_24 gnd C_bl
Cbb_39_24 bitb_39_24 gnd C_bl
Rb_39_25 bit_39_25 bit_39_26 R_bl
Rbb_39_25 bitb_39_25 bitb_39_26 R_bl
Cb_39_25 bit_39_25 gnd C_bl
Cbb_39_25 bitb_39_25 gnd C_bl
Rb_39_26 bit_39_26 bit_39_27 R_bl
Rbb_39_26 bitb_39_26 bitb_39_27 R_bl
Cb_39_26 bit_39_26 gnd C_bl
Cbb_39_26 bitb_39_26 gnd C_bl
Rb_39_27 bit_39_27 bit_39_28 R_bl
Rbb_39_27 bitb_39_27 bitb_39_28 R_bl
Cb_39_27 bit_39_27 gnd C_bl
Cbb_39_27 bitb_39_27 gnd C_bl
Rb_39_28 bit_39_28 bit_39_29 R_bl
Rbb_39_28 bitb_39_28 bitb_39_29 R_bl
Cb_39_28 bit_39_28 gnd C_bl
Cbb_39_28 bitb_39_28 gnd C_bl
Rb_39_29 bit_39_29 bit_39_30 R_bl
Rbb_39_29 bitb_39_29 bitb_39_30 R_bl
Cb_39_29 bit_39_29 gnd C_bl
Cbb_39_29 bitb_39_29 gnd C_bl
Rb_39_30 bit_39_30 bit_39_31 R_bl
Rbb_39_30 bitb_39_30 bitb_39_31 R_bl
Cb_39_30 bit_39_30 gnd C_bl
Cbb_39_30 bitb_39_30 gnd C_bl
Rb_39_31 bit_39_31 bit_39_32 R_bl
Rbb_39_31 bitb_39_31 bitb_39_32 R_bl
Cb_39_31 bit_39_31 gnd C_bl
Cbb_39_31 bitb_39_31 gnd C_bl
Rb_39_32 bit_39_32 bit_39_33 R_bl
Rbb_39_32 bitb_39_32 bitb_39_33 R_bl
Cb_39_32 bit_39_32 gnd C_bl
Cbb_39_32 bitb_39_32 gnd C_bl
Rb_39_33 bit_39_33 bit_39_34 R_bl
Rbb_39_33 bitb_39_33 bitb_39_34 R_bl
Cb_39_33 bit_39_33 gnd C_bl
Cbb_39_33 bitb_39_33 gnd C_bl
Rb_39_34 bit_39_34 bit_39_35 R_bl
Rbb_39_34 bitb_39_34 bitb_39_35 R_bl
Cb_39_34 bit_39_34 gnd C_bl
Cbb_39_34 bitb_39_34 gnd C_bl
Rb_39_35 bit_39_35 bit_39_36 R_bl
Rbb_39_35 bitb_39_35 bitb_39_36 R_bl
Cb_39_35 bit_39_35 gnd C_bl
Cbb_39_35 bitb_39_35 gnd C_bl
Rb_39_36 bit_39_36 bit_39_37 R_bl
Rbb_39_36 bitb_39_36 bitb_39_37 R_bl
Cb_39_36 bit_39_36 gnd C_bl
Cbb_39_36 bitb_39_36 gnd C_bl
Rb_39_37 bit_39_37 bit_39_38 R_bl
Rbb_39_37 bitb_39_37 bitb_39_38 R_bl
Cb_39_37 bit_39_37 gnd C_bl
Cbb_39_37 bitb_39_37 gnd C_bl
Rb_39_38 bit_39_38 bit_39_39 R_bl
Rbb_39_38 bitb_39_38 bitb_39_39 R_bl
Cb_39_38 bit_39_38 gnd C_bl
Cbb_39_38 bitb_39_38 gnd C_bl
Rb_39_39 bit_39_39 bit_39_40 R_bl
Rbb_39_39 bitb_39_39 bitb_39_40 R_bl
Cb_39_39 bit_39_39 gnd C_bl
Cbb_39_39 bitb_39_39 gnd C_bl
Rb_39_40 bit_39_40 bit_39_41 R_bl
Rbb_39_40 bitb_39_40 bitb_39_41 R_bl
Cb_39_40 bit_39_40 gnd C_bl
Cbb_39_40 bitb_39_40 gnd C_bl
Rb_39_41 bit_39_41 bit_39_42 R_bl
Rbb_39_41 bitb_39_41 bitb_39_42 R_bl
Cb_39_41 bit_39_41 gnd C_bl
Cbb_39_41 bitb_39_41 gnd C_bl
Rb_39_42 bit_39_42 bit_39_43 R_bl
Rbb_39_42 bitb_39_42 bitb_39_43 R_bl
Cb_39_42 bit_39_42 gnd C_bl
Cbb_39_42 bitb_39_42 gnd C_bl
Rb_39_43 bit_39_43 bit_39_44 R_bl
Rbb_39_43 bitb_39_43 bitb_39_44 R_bl
Cb_39_43 bit_39_43 gnd C_bl
Cbb_39_43 bitb_39_43 gnd C_bl
Rb_39_44 bit_39_44 bit_39_45 R_bl
Rbb_39_44 bitb_39_44 bitb_39_45 R_bl
Cb_39_44 bit_39_44 gnd C_bl
Cbb_39_44 bitb_39_44 gnd C_bl
Rb_39_45 bit_39_45 bit_39_46 R_bl
Rbb_39_45 bitb_39_45 bitb_39_46 R_bl
Cb_39_45 bit_39_45 gnd C_bl
Cbb_39_45 bitb_39_45 gnd C_bl
Rb_39_46 bit_39_46 bit_39_47 R_bl
Rbb_39_46 bitb_39_46 bitb_39_47 R_bl
Cb_39_46 bit_39_46 gnd C_bl
Cbb_39_46 bitb_39_46 gnd C_bl
Rb_39_47 bit_39_47 bit_39_48 R_bl
Rbb_39_47 bitb_39_47 bitb_39_48 R_bl
Cb_39_47 bit_39_47 gnd C_bl
Cbb_39_47 bitb_39_47 gnd C_bl
Rb_39_48 bit_39_48 bit_39_49 R_bl
Rbb_39_48 bitb_39_48 bitb_39_49 R_bl
Cb_39_48 bit_39_48 gnd C_bl
Cbb_39_48 bitb_39_48 gnd C_bl
Rb_39_49 bit_39_49 bit_39_50 R_bl
Rbb_39_49 bitb_39_49 bitb_39_50 R_bl
Cb_39_49 bit_39_49 gnd C_bl
Cbb_39_49 bitb_39_49 gnd C_bl
Rb_39_50 bit_39_50 bit_39_51 R_bl
Rbb_39_50 bitb_39_50 bitb_39_51 R_bl
Cb_39_50 bit_39_50 gnd C_bl
Cbb_39_50 bitb_39_50 gnd C_bl
Rb_39_51 bit_39_51 bit_39_52 R_bl
Rbb_39_51 bitb_39_51 bitb_39_52 R_bl
Cb_39_51 bit_39_51 gnd C_bl
Cbb_39_51 bitb_39_51 gnd C_bl
Rb_39_52 bit_39_52 bit_39_53 R_bl
Rbb_39_52 bitb_39_52 bitb_39_53 R_bl
Cb_39_52 bit_39_52 gnd C_bl
Cbb_39_52 bitb_39_52 gnd C_bl
Rb_39_53 bit_39_53 bit_39_54 R_bl
Rbb_39_53 bitb_39_53 bitb_39_54 R_bl
Cb_39_53 bit_39_53 gnd C_bl
Cbb_39_53 bitb_39_53 gnd C_bl
Rb_39_54 bit_39_54 bit_39_55 R_bl
Rbb_39_54 bitb_39_54 bitb_39_55 R_bl
Cb_39_54 bit_39_54 gnd C_bl
Cbb_39_54 bitb_39_54 gnd C_bl
Rb_39_55 bit_39_55 bit_39_56 R_bl
Rbb_39_55 bitb_39_55 bitb_39_56 R_bl
Cb_39_55 bit_39_55 gnd C_bl
Cbb_39_55 bitb_39_55 gnd C_bl
Rb_39_56 bit_39_56 bit_39_57 R_bl
Rbb_39_56 bitb_39_56 bitb_39_57 R_bl
Cb_39_56 bit_39_56 gnd C_bl
Cbb_39_56 bitb_39_56 gnd C_bl
Rb_39_57 bit_39_57 bit_39_58 R_bl
Rbb_39_57 bitb_39_57 bitb_39_58 R_bl
Cb_39_57 bit_39_57 gnd C_bl
Cbb_39_57 bitb_39_57 gnd C_bl
Rb_39_58 bit_39_58 bit_39_59 R_bl
Rbb_39_58 bitb_39_58 bitb_39_59 R_bl
Cb_39_58 bit_39_58 gnd C_bl
Cbb_39_58 bitb_39_58 gnd C_bl
Rb_39_59 bit_39_59 bit_39_60 R_bl
Rbb_39_59 bitb_39_59 bitb_39_60 R_bl
Cb_39_59 bit_39_59 gnd C_bl
Cbb_39_59 bitb_39_59 gnd C_bl
Rb_39_60 bit_39_60 bit_39_61 R_bl
Rbb_39_60 bitb_39_60 bitb_39_61 R_bl
Cb_39_60 bit_39_60 gnd C_bl
Cbb_39_60 bitb_39_60 gnd C_bl
Rb_39_61 bit_39_61 bit_39_62 R_bl
Rbb_39_61 bitb_39_61 bitb_39_62 R_bl
Cb_39_61 bit_39_61 gnd C_bl
Cbb_39_61 bitb_39_61 gnd C_bl
Rb_39_62 bit_39_62 bit_39_63 R_bl
Rbb_39_62 bitb_39_62 bitb_39_63 R_bl
Cb_39_62 bit_39_62 gnd C_bl
Cbb_39_62 bitb_39_62 gnd C_bl
Rb_39_63 bit_39_63 bit_39_64 R_bl
Rbb_39_63 bitb_39_63 bitb_39_64 R_bl
Cb_39_63 bit_39_63 gnd C_bl
Cbb_39_63 bitb_39_63 gnd C_bl
Rb_39_64 bit_39_64 bit_39_65 R_bl
Rbb_39_64 bitb_39_64 bitb_39_65 R_bl
Cb_39_64 bit_39_64 gnd C_bl
Cbb_39_64 bitb_39_64 gnd C_bl
Rb_39_65 bit_39_65 bit_39_66 R_bl
Rbb_39_65 bitb_39_65 bitb_39_66 R_bl
Cb_39_65 bit_39_65 gnd C_bl
Cbb_39_65 bitb_39_65 gnd C_bl
Rb_39_66 bit_39_66 bit_39_67 R_bl
Rbb_39_66 bitb_39_66 bitb_39_67 R_bl
Cb_39_66 bit_39_66 gnd C_bl
Cbb_39_66 bitb_39_66 gnd C_bl
Rb_39_67 bit_39_67 bit_39_68 R_bl
Rbb_39_67 bitb_39_67 bitb_39_68 R_bl
Cb_39_67 bit_39_67 gnd C_bl
Cbb_39_67 bitb_39_67 gnd C_bl
Rb_39_68 bit_39_68 bit_39_69 R_bl
Rbb_39_68 bitb_39_68 bitb_39_69 R_bl
Cb_39_68 bit_39_68 gnd C_bl
Cbb_39_68 bitb_39_68 gnd C_bl
Rb_39_69 bit_39_69 bit_39_70 R_bl
Rbb_39_69 bitb_39_69 bitb_39_70 R_bl
Cb_39_69 bit_39_69 gnd C_bl
Cbb_39_69 bitb_39_69 gnd C_bl
Rb_39_70 bit_39_70 bit_39_71 R_bl
Rbb_39_70 bitb_39_70 bitb_39_71 R_bl
Cb_39_70 bit_39_70 gnd C_bl
Cbb_39_70 bitb_39_70 gnd C_bl
Rb_39_71 bit_39_71 bit_39_72 R_bl
Rbb_39_71 bitb_39_71 bitb_39_72 R_bl
Cb_39_71 bit_39_71 gnd C_bl
Cbb_39_71 bitb_39_71 gnd C_bl
Rb_39_72 bit_39_72 bit_39_73 R_bl
Rbb_39_72 bitb_39_72 bitb_39_73 R_bl
Cb_39_72 bit_39_72 gnd C_bl
Cbb_39_72 bitb_39_72 gnd C_bl
Rb_39_73 bit_39_73 bit_39_74 R_bl
Rbb_39_73 bitb_39_73 bitb_39_74 R_bl
Cb_39_73 bit_39_73 gnd C_bl
Cbb_39_73 bitb_39_73 gnd C_bl
Rb_39_74 bit_39_74 bit_39_75 R_bl
Rbb_39_74 bitb_39_74 bitb_39_75 R_bl
Cb_39_74 bit_39_74 gnd C_bl
Cbb_39_74 bitb_39_74 gnd C_bl
Rb_39_75 bit_39_75 bit_39_76 R_bl
Rbb_39_75 bitb_39_75 bitb_39_76 R_bl
Cb_39_75 bit_39_75 gnd C_bl
Cbb_39_75 bitb_39_75 gnd C_bl
Rb_39_76 bit_39_76 bit_39_77 R_bl
Rbb_39_76 bitb_39_76 bitb_39_77 R_bl
Cb_39_76 bit_39_76 gnd C_bl
Cbb_39_76 bitb_39_76 gnd C_bl
Rb_39_77 bit_39_77 bit_39_78 R_bl
Rbb_39_77 bitb_39_77 bitb_39_78 R_bl
Cb_39_77 bit_39_77 gnd C_bl
Cbb_39_77 bitb_39_77 gnd C_bl
Rb_39_78 bit_39_78 bit_39_79 R_bl
Rbb_39_78 bitb_39_78 bitb_39_79 R_bl
Cb_39_78 bit_39_78 gnd C_bl
Cbb_39_78 bitb_39_78 gnd C_bl
Rb_39_79 bit_39_79 bit_39_80 R_bl
Rbb_39_79 bitb_39_79 bitb_39_80 R_bl
Cb_39_79 bit_39_79 gnd C_bl
Cbb_39_79 bitb_39_79 gnd C_bl
Rb_39_80 bit_39_80 bit_39_81 R_bl
Rbb_39_80 bitb_39_80 bitb_39_81 R_bl
Cb_39_80 bit_39_80 gnd C_bl
Cbb_39_80 bitb_39_80 gnd C_bl
Rb_39_81 bit_39_81 bit_39_82 R_bl
Rbb_39_81 bitb_39_81 bitb_39_82 R_bl
Cb_39_81 bit_39_81 gnd C_bl
Cbb_39_81 bitb_39_81 gnd C_bl
Rb_39_82 bit_39_82 bit_39_83 R_bl
Rbb_39_82 bitb_39_82 bitb_39_83 R_bl
Cb_39_82 bit_39_82 gnd C_bl
Cbb_39_82 bitb_39_82 gnd C_bl
Rb_39_83 bit_39_83 bit_39_84 R_bl
Rbb_39_83 bitb_39_83 bitb_39_84 R_bl
Cb_39_83 bit_39_83 gnd C_bl
Cbb_39_83 bitb_39_83 gnd C_bl
Rb_39_84 bit_39_84 bit_39_85 R_bl
Rbb_39_84 bitb_39_84 bitb_39_85 R_bl
Cb_39_84 bit_39_84 gnd C_bl
Cbb_39_84 bitb_39_84 gnd C_bl
Rb_39_85 bit_39_85 bit_39_86 R_bl
Rbb_39_85 bitb_39_85 bitb_39_86 R_bl
Cb_39_85 bit_39_85 gnd C_bl
Cbb_39_85 bitb_39_85 gnd C_bl
Rb_39_86 bit_39_86 bit_39_87 R_bl
Rbb_39_86 bitb_39_86 bitb_39_87 R_bl
Cb_39_86 bit_39_86 gnd C_bl
Cbb_39_86 bitb_39_86 gnd C_bl
Rb_39_87 bit_39_87 bit_39_88 R_bl
Rbb_39_87 bitb_39_87 bitb_39_88 R_bl
Cb_39_87 bit_39_87 gnd C_bl
Cbb_39_87 bitb_39_87 gnd C_bl
Rb_39_88 bit_39_88 bit_39_89 R_bl
Rbb_39_88 bitb_39_88 bitb_39_89 R_bl
Cb_39_88 bit_39_88 gnd C_bl
Cbb_39_88 bitb_39_88 gnd C_bl
Rb_39_89 bit_39_89 bit_39_90 R_bl
Rbb_39_89 bitb_39_89 bitb_39_90 R_bl
Cb_39_89 bit_39_89 gnd C_bl
Cbb_39_89 bitb_39_89 gnd C_bl
Rb_39_90 bit_39_90 bit_39_91 R_bl
Rbb_39_90 bitb_39_90 bitb_39_91 R_bl
Cb_39_90 bit_39_90 gnd C_bl
Cbb_39_90 bitb_39_90 gnd C_bl
Rb_39_91 bit_39_91 bit_39_92 R_bl
Rbb_39_91 bitb_39_91 bitb_39_92 R_bl
Cb_39_91 bit_39_91 gnd C_bl
Cbb_39_91 bitb_39_91 gnd C_bl
Rb_39_92 bit_39_92 bit_39_93 R_bl
Rbb_39_92 bitb_39_92 bitb_39_93 R_bl
Cb_39_92 bit_39_92 gnd C_bl
Cbb_39_92 bitb_39_92 gnd C_bl
Rb_39_93 bit_39_93 bit_39_94 R_bl
Rbb_39_93 bitb_39_93 bitb_39_94 R_bl
Cb_39_93 bit_39_93 gnd C_bl
Cbb_39_93 bitb_39_93 gnd C_bl
Rb_39_94 bit_39_94 bit_39_95 R_bl
Rbb_39_94 bitb_39_94 bitb_39_95 R_bl
Cb_39_94 bit_39_94 gnd C_bl
Cbb_39_94 bitb_39_94 gnd C_bl
Rb_39_95 bit_39_95 bit_39_96 R_bl
Rbb_39_95 bitb_39_95 bitb_39_96 R_bl
Cb_39_95 bit_39_95 gnd C_bl
Cbb_39_95 bitb_39_95 gnd C_bl
Rb_39_96 bit_39_96 bit_39_97 R_bl
Rbb_39_96 bitb_39_96 bitb_39_97 R_bl
Cb_39_96 bit_39_96 gnd C_bl
Cbb_39_96 bitb_39_96 gnd C_bl
Rb_39_97 bit_39_97 bit_39_98 R_bl
Rbb_39_97 bitb_39_97 bitb_39_98 R_bl
Cb_39_97 bit_39_97 gnd C_bl
Cbb_39_97 bitb_39_97 gnd C_bl
Rb_39_98 bit_39_98 bit_39_99 R_bl
Rbb_39_98 bitb_39_98 bitb_39_99 R_bl
Cb_39_98 bit_39_98 gnd C_bl
Cbb_39_98 bitb_39_98 gnd C_bl
Rb_39_99 bit_39_99 bit_39_100 R_bl
Rbb_39_99 bitb_39_99 bitb_39_100 R_bl
Cb_39_99 bit_39_99 gnd C_bl
Cbb_39_99 bitb_39_99 gnd C_bl
Rb_40_0 bit_40_0 bit_40_1 R_bl
Rbb_40_0 bitb_40_0 bitb_40_1 R_bl
Cb_40_0 bit_40_0 gnd C_bl
Cbb_40_0 bitb_40_0 gnd C_bl
Rb_40_1 bit_40_1 bit_40_2 R_bl
Rbb_40_1 bitb_40_1 bitb_40_2 R_bl
Cb_40_1 bit_40_1 gnd C_bl
Cbb_40_1 bitb_40_1 gnd C_bl
Rb_40_2 bit_40_2 bit_40_3 R_bl
Rbb_40_2 bitb_40_2 bitb_40_3 R_bl
Cb_40_2 bit_40_2 gnd C_bl
Cbb_40_2 bitb_40_2 gnd C_bl
Rb_40_3 bit_40_3 bit_40_4 R_bl
Rbb_40_3 bitb_40_3 bitb_40_4 R_bl
Cb_40_3 bit_40_3 gnd C_bl
Cbb_40_3 bitb_40_3 gnd C_bl
Rb_40_4 bit_40_4 bit_40_5 R_bl
Rbb_40_4 bitb_40_4 bitb_40_5 R_bl
Cb_40_4 bit_40_4 gnd C_bl
Cbb_40_4 bitb_40_4 gnd C_bl
Rb_40_5 bit_40_5 bit_40_6 R_bl
Rbb_40_5 bitb_40_5 bitb_40_6 R_bl
Cb_40_5 bit_40_5 gnd C_bl
Cbb_40_5 bitb_40_5 gnd C_bl
Rb_40_6 bit_40_6 bit_40_7 R_bl
Rbb_40_6 bitb_40_6 bitb_40_7 R_bl
Cb_40_6 bit_40_6 gnd C_bl
Cbb_40_6 bitb_40_6 gnd C_bl
Rb_40_7 bit_40_7 bit_40_8 R_bl
Rbb_40_7 bitb_40_7 bitb_40_8 R_bl
Cb_40_7 bit_40_7 gnd C_bl
Cbb_40_7 bitb_40_7 gnd C_bl
Rb_40_8 bit_40_8 bit_40_9 R_bl
Rbb_40_8 bitb_40_8 bitb_40_9 R_bl
Cb_40_8 bit_40_8 gnd C_bl
Cbb_40_8 bitb_40_8 gnd C_bl
Rb_40_9 bit_40_9 bit_40_10 R_bl
Rbb_40_9 bitb_40_9 bitb_40_10 R_bl
Cb_40_9 bit_40_9 gnd C_bl
Cbb_40_9 bitb_40_9 gnd C_bl
Rb_40_10 bit_40_10 bit_40_11 R_bl
Rbb_40_10 bitb_40_10 bitb_40_11 R_bl
Cb_40_10 bit_40_10 gnd C_bl
Cbb_40_10 bitb_40_10 gnd C_bl
Rb_40_11 bit_40_11 bit_40_12 R_bl
Rbb_40_11 bitb_40_11 bitb_40_12 R_bl
Cb_40_11 bit_40_11 gnd C_bl
Cbb_40_11 bitb_40_11 gnd C_bl
Rb_40_12 bit_40_12 bit_40_13 R_bl
Rbb_40_12 bitb_40_12 bitb_40_13 R_bl
Cb_40_12 bit_40_12 gnd C_bl
Cbb_40_12 bitb_40_12 gnd C_bl
Rb_40_13 bit_40_13 bit_40_14 R_bl
Rbb_40_13 bitb_40_13 bitb_40_14 R_bl
Cb_40_13 bit_40_13 gnd C_bl
Cbb_40_13 bitb_40_13 gnd C_bl
Rb_40_14 bit_40_14 bit_40_15 R_bl
Rbb_40_14 bitb_40_14 bitb_40_15 R_bl
Cb_40_14 bit_40_14 gnd C_bl
Cbb_40_14 bitb_40_14 gnd C_bl
Rb_40_15 bit_40_15 bit_40_16 R_bl
Rbb_40_15 bitb_40_15 bitb_40_16 R_bl
Cb_40_15 bit_40_15 gnd C_bl
Cbb_40_15 bitb_40_15 gnd C_bl
Rb_40_16 bit_40_16 bit_40_17 R_bl
Rbb_40_16 bitb_40_16 bitb_40_17 R_bl
Cb_40_16 bit_40_16 gnd C_bl
Cbb_40_16 bitb_40_16 gnd C_bl
Rb_40_17 bit_40_17 bit_40_18 R_bl
Rbb_40_17 bitb_40_17 bitb_40_18 R_bl
Cb_40_17 bit_40_17 gnd C_bl
Cbb_40_17 bitb_40_17 gnd C_bl
Rb_40_18 bit_40_18 bit_40_19 R_bl
Rbb_40_18 bitb_40_18 bitb_40_19 R_bl
Cb_40_18 bit_40_18 gnd C_bl
Cbb_40_18 bitb_40_18 gnd C_bl
Rb_40_19 bit_40_19 bit_40_20 R_bl
Rbb_40_19 bitb_40_19 bitb_40_20 R_bl
Cb_40_19 bit_40_19 gnd C_bl
Cbb_40_19 bitb_40_19 gnd C_bl
Rb_40_20 bit_40_20 bit_40_21 R_bl
Rbb_40_20 bitb_40_20 bitb_40_21 R_bl
Cb_40_20 bit_40_20 gnd C_bl
Cbb_40_20 bitb_40_20 gnd C_bl
Rb_40_21 bit_40_21 bit_40_22 R_bl
Rbb_40_21 bitb_40_21 bitb_40_22 R_bl
Cb_40_21 bit_40_21 gnd C_bl
Cbb_40_21 bitb_40_21 gnd C_bl
Rb_40_22 bit_40_22 bit_40_23 R_bl
Rbb_40_22 bitb_40_22 bitb_40_23 R_bl
Cb_40_22 bit_40_22 gnd C_bl
Cbb_40_22 bitb_40_22 gnd C_bl
Rb_40_23 bit_40_23 bit_40_24 R_bl
Rbb_40_23 bitb_40_23 bitb_40_24 R_bl
Cb_40_23 bit_40_23 gnd C_bl
Cbb_40_23 bitb_40_23 gnd C_bl
Rb_40_24 bit_40_24 bit_40_25 R_bl
Rbb_40_24 bitb_40_24 bitb_40_25 R_bl
Cb_40_24 bit_40_24 gnd C_bl
Cbb_40_24 bitb_40_24 gnd C_bl
Rb_40_25 bit_40_25 bit_40_26 R_bl
Rbb_40_25 bitb_40_25 bitb_40_26 R_bl
Cb_40_25 bit_40_25 gnd C_bl
Cbb_40_25 bitb_40_25 gnd C_bl
Rb_40_26 bit_40_26 bit_40_27 R_bl
Rbb_40_26 bitb_40_26 bitb_40_27 R_bl
Cb_40_26 bit_40_26 gnd C_bl
Cbb_40_26 bitb_40_26 gnd C_bl
Rb_40_27 bit_40_27 bit_40_28 R_bl
Rbb_40_27 bitb_40_27 bitb_40_28 R_bl
Cb_40_27 bit_40_27 gnd C_bl
Cbb_40_27 bitb_40_27 gnd C_bl
Rb_40_28 bit_40_28 bit_40_29 R_bl
Rbb_40_28 bitb_40_28 bitb_40_29 R_bl
Cb_40_28 bit_40_28 gnd C_bl
Cbb_40_28 bitb_40_28 gnd C_bl
Rb_40_29 bit_40_29 bit_40_30 R_bl
Rbb_40_29 bitb_40_29 bitb_40_30 R_bl
Cb_40_29 bit_40_29 gnd C_bl
Cbb_40_29 bitb_40_29 gnd C_bl
Rb_40_30 bit_40_30 bit_40_31 R_bl
Rbb_40_30 bitb_40_30 bitb_40_31 R_bl
Cb_40_30 bit_40_30 gnd C_bl
Cbb_40_30 bitb_40_30 gnd C_bl
Rb_40_31 bit_40_31 bit_40_32 R_bl
Rbb_40_31 bitb_40_31 bitb_40_32 R_bl
Cb_40_31 bit_40_31 gnd C_bl
Cbb_40_31 bitb_40_31 gnd C_bl
Rb_40_32 bit_40_32 bit_40_33 R_bl
Rbb_40_32 bitb_40_32 bitb_40_33 R_bl
Cb_40_32 bit_40_32 gnd C_bl
Cbb_40_32 bitb_40_32 gnd C_bl
Rb_40_33 bit_40_33 bit_40_34 R_bl
Rbb_40_33 bitb_40_33 bitb_40_34 R_bl
Cb_40_33 bit_40_33 gnd C_bl
Cbb_40_33 bitb_40_33 gnd C_bl
Rb_40_34 bit_40_34 bit_40_35 R_bl
Rbb_40_34 bitb_40_34 bitb_40_35 R_bl
Cb_40_34 bit_40_34 gnd C_bl
Cbb_40_34 bitb_40_34 gnd C_bl
Rb_40_35 bit_40_35 bit_40_36 R_bl
Rbb_40_35 bitb_40_35 bitb_40_36 R_bl
Cb_40_35 bit_40_35 gnd C_bl
Cbb_40_35 bitb_40_35 gnd C_bl
Rb_40_36 bit_40_36 bit_40_37 R_bl
Rbb_40_36 bitb_40_36 bitb_40_37 R_bl
Cb_40_36 bit_40_36 gnd C_bl
Cbb_40_36 bitb_40_36 gnd C_bl
Rb_40_37 bit_40_37 bit_40_38 R_bl
Rbb_40_37 bitb_40_37 bitb_40_38 R_bl
Cb_40_37 bit_40_37 gnd C_bl
Cbb_40_37 bitb_40_37 gnd C_bl
Rb_40_38 bit_40_38 bit_40_39 R_bl
Rbb_40_38 bitb_40_38 bitb_40_39 R_bl
Cb_40_38 bit_40_38 gnd C_bl
Cbb_40_38 bitb_40_38 gnd C_bl
Rb_40_39 bit_40_39 bit_40_40 R_bl
Rbb_40_39 bitb_40_39 bitb_40_40 R_bl
Cb_40_39 bit_40_39 gnd C_bl
Cbb_40_39 bitb_40_39 gnd C_bl
Rb_40_40 bit_40_40 bit_40_41 R_bl
Rbb_40_40 bitb_40_40 bitb_40_41 R_bl
Cb_40_40 bit_40_40 gnd C_bl
Cbb_40_40 bitb_40_40 gnd C_bl
Rb_40_41 bit_40_41 bit_40_42 R_bl
Rbb_40_41 bitb_40_41 bitb_40_42 R_bl
Cb_40_41 bit_40_41 gnd C_bl
Cbb_40_41 bitb_40_41 gnd C_bl
Rb_40_42 bit_40_42 bit_40_43 R_bl
Rbb_40_42 bitb_40_42 bitb_40_43 R_bl
Cb_40_42 bit_40_42 gnd C_bl
Cbb_40_42 bitb_40_42 gnd C_bl
Rb_40_43 bit_40_43 bit_40_44 R_bl
Rbb_40_43 bitb_40_43 bitb_40_44 R_bl
Cb_40_43 bit_40_43 gnd C_bl
Cbb_40_43 bitb_40_43 gnd C_bl
Rb_40_44 bit_40_44 bit_40_45 R_bl
Rbb_40_44 bitb_40_44 bitb_40_45 R_bl
Cb_40_44 bit_40_44 gnd C_bl
Cbb_40_44 bitb_40_44 gnd C_bl
Rb_40_45 bit_40_45 bit_40_46 R_bl
Rbb_40_45 bitb_40_45 bitb_40_46 R_bl
Cb_40_45 bit_40_45 gnd C_bl
Cbb_40_45 bitb_40_45 gnd C_bl
Rb_40_46 bit_40_46 bit_40_47 R_bl
Rbb_40_46 bitb_40_46 bitb_40_47 R_bl
Cb_40_46 bit_40_46 gnd C_bl
Cbb_40_46 bitb_40_46 gnd C_bl
Rb_40_47 bit_40_47 bit_40_48 R_bl
Rbb_40_47 bitb_40_47 bitb_40_48 R_bl
Cb_40_47 bit_40_47 gnd C_bl
Cbb_40_47 bitb_40_47 gnd C_bl
Rb_40_48 bit_40_48 bit_40_49 R_bl
Rbb_40_48 bitb_40_48 bitb_40_49 R_bl
Cb_40_48 bit_40_48 gnd C_bl
Cbb_40_48 bitb_40_48 gnd C_bl
Rb_40_49 bit_40_49 bit_40_50 R_bl
Rbb_40_49 bitb_40_49 bitb_40_50 R_bl
Cb_40_49 bit_40_49 gnd C_bl
Cbb_40_49 bitb_40_49 gnd C_bl
Rb_40_50 bit_40_50 bit_40_51 R_bl
Rbb_40_50 bitb_40_50 bitb_40_51 R_bl
Cb_40_50 bit_40_50 gnd C_bl
Cbb_40_50 bitb_40_50 gnd C_bl
Rb_40_51 bit_40_51 bit_40_52 R_bl
Rbb_40_51 bitb_40_51 bitb_40_52 R_bl
Cb_40_51 bit_40_51 gnd C_bl
Cbb_40_51 bitb_40_51 gnd C_bl
Rb_40_52 bit_40_52 bit_40_53 R_bl
Rbb_40_52 bitb_40_52 bitb_40_53 R_bl
Cb_40_52 bit_40_52 gnd C_bl
Cbb_40_52 bitb_40_52 gnd C_bl
Rb_40_53 bit_40_53 bit_40_54 R_bl
Rbb_40_53 bitb_40_53 bitb_40_54 R_bl
Cb_40_53 bit_40_53 gnd C_bl
Cbb_40_53 bitb_40_53 gnd C_bl
Rb_40_54 bit_40_54 bit_40_55 R_bl
Rbb_40_54 bitb_40_54 bitb_40_55 R_bl
Cb_40_54 bit_40_54 gnd C_bl
Cbb_40_54 bitb_40_54 gnd C_bl
Rb_40_55 bit_40_55 bit_40_56 R_bl
Rbb_40_55 bitb_40_55 bitb_40_56 R_bl
Cb_40_55 bit_40_55 gnd C_bl
Cbb_40_55 bitb_40_55 gnd C_bl
Rb_40_56 bit_40_56 bit_40_57 R_bl
Rbb_40_56 bitb_40_56 bitb_40_57 R_bl
Cb_40_56 bit_40_56 gnd C_bl
Cbb_40_56 bitb_40_56 gnd C_bl
Rb_40_57 bit_40_57 bit_40_58 R_bl
Rbb_40_57 bitb_40_57 bitb_40_58 R_bl
Cb_40_57 bit_40_57 gnd C_bl
Cbb_40_57 bitb_40_57 gnd C_bl
Rb_40_58 bit_40_58 bit_40_59 R_bl
Rbb_40_58 bitb_40_58 bitb_40_59 R_bl
Cb_40_58 bit_40_58 gnd C_bl
Cbb_40_58 bitb_40_58 gnd C_bl
Rb_40_59 bit_40_59 bit_40_60 R_bl
Rbb_40_59 bitb_40_59 bitb_40_60 R_bl
Cb_40_59 bit_40_59 gnd C_bl
Cbb_40_59 bitb_40_59 gnd C_bl
Rb_40_60 bit_40_60 bit_40_61 R_bl
Rbb_40_60 bitb_40_60 bitb_40_61 R_bl
Cb_40_60 bit_40_60 gnd C_bl
Cbb_40_60 bitb_40_60 gnd C_bl
Rb_40_61 bit_40_61 bit_40_62 R_bl
Rbb_40_61 bitb_40_61 bitb_40_62 R_bl
Cb_40_61 bit_40_61 gnd C_bl
Cbb_40_61 bitb_40_61 gnd C_bl
Rb_40_62 bit_40_62 bit_40_63 R_bl
Rbb_40_62 bitb_40_62 bitb_40_63 R_bl
Cb_40_62 bit_40_62 gnd C_bl
Cbb_40_62 bitb_40_62 gnd C_bl
Rb_40_63 bit_40_63 bit_40_64 R_bl
Rbb_40_63 bitb_40_63 bitb_40_64 R_bl
Cb_40_63 bit_40_63 gnd C_bl
Cbb_40_63 bitb_40_63 gnd C_bl
Rb_40_64 bit_40_64 bit_40_65 R_bl
Rbb_40_64 bitb_40_64 bitb_40_65 R_bl
Cb_40_64 bit_40_64 gnd C_bl
Cbb_40_64 bitb_40_64 gnd C_bl
Rb_40_65 bit_40_65 bit_40_66 R_bl
Rbb_40_65 bitb_40_65 bitb_40_66 R_bl
Cb_40_65 bit_40_65 gnd C_bl
Cbb_40_65 bitb_40_65 gnd C_bl
Rb_40_66 bit_40_66 bit_40_67 R_bl
Rbb_40_66 bitb_40_66 bitb_40_67 R_bl
Cb_40_66 bit_40_66 gnd C_bl
Cbb_40_66 bitb_40_66 gnd C_bl
Rb_40_67 bit_40_67 bit_40_68 R_bl
Rbb_40_67 bitb_40_67 bitb_40_68 R_bl
Cb_40_67 bit_40_67 gnd C_bl
Cbb_40_67 bitb_40_67 gnd C_bl
Rb_40_68 bit_40_68 bit_40_69 R_bl
Rbb_40_68 bitb_40_68 bitb_40_69 R_bl
Cb_40_68 bit_40_68 gnd C_bl
Cbb_40_68 bitb_40_68 gnd C_bl
Rb_40_69 bit_40_69 bit_40_70 R_bl
Rbb_40_69 bitb_40_69 bitb_40_70 R_bl
Cb_40_69 bit_40_69 gnd C_bl
Cbb_40_69 bitb_40_69 gnd C_bl
Rb_40_70 bit_40_70 bit_40_71 R_bl
Rbb_40_70 bitb_40_70 bitb_40_71 R_bl
Cb_40_70 bit_40_70 gnd C_bl
Cbb_40_70 bitb_40_70 gnd C_bl
Rb_40_71 bit_40_71 bit_40_72 R_bl
Rbb_40_71 bitb_40_71 bitb_40_72 R_bl
Cb_40_71 bit_40_71 gnd C_bl
Cbb_40_71 bitb_40_71 gnd C_bl
Rb_40_72 bit_40_72 bit_40_73 R_bl
Rbb_40_72 bitb_40_72 bitb_40_73 R_bl
Cb_40_72 bit_40_72 gnd C_bl
Cbb_40_72 bitb_40_72 gnd C_bl
Rb_40_73 bit_40_73 bit_40_74 R_bl
Rbb_40_73 bitb_40_73 bitb_40_74 R_bl
Cb_40_73 bit_40_73 gnd C_bl
Cbb_40_73 bitb_40_73 gnd C_bl
Rb_40_74 bit_40_74 bit_40_75 R_bl
Rbb_40_74 bitb_40_74 bitb_40_75 R_bl
Cb_40_74 bit_40_74 gnd C_bl
Cbb_40_74 bitb_40_74 gnd C_bl
Rb_40_75 bit_40_75 bit_40_76 R_bl
Rbb_40_75 bitb_40_75 bitb_40_76 R_bl
Cb_40_75 bit_40_75 gnd C_bl
Cbb_40_75 bitb_40_75 gnd C_bl
Rb_40_76 bit_40_76 bit_40_77 R_bl
Rbb_40_76 bitb_40_76 bitb_40_77 R_bl
Cb_40_76 bit_40_76 gnd C_bl
Cbb_40_76 bitb_40_76 gnd C_bl
Rb_40_77 bit_40_77 bit_40_78 R_bl
Rbb_40_77 bitb_40_77 bitb_40_78 R_bl
Cb_40_77 bit_40_77 gnd C_bl
Cbb_40_77 bitb_40_77 gnd C_bl
Rb_40_78 bit_40_78 bit_40_79 R_bl
Rbb_40_78 bitb_40_78 bitb_40_79 R_bl
Cb_40_78 bit_40_78 gnd C_bl
Cbb_40_78 bitb_40_78 gnd C_bl
Rb_40_79 bit_40_79 bit_40_80 R_bl
Rbb_40_79 bitb_40_79 bitb_40_80 R_bl
Cb_40_79 bit_40_79 gnd C_bl
Cbb_40_79 bitb_40_79 gnd C_bl
Rb_40_80 bit_40_80 bit_40_81 R_bl
Rbb_40_80 bitb_40_80 bitb_40_81 R_bl
Cb_40_80 bit_40_80 gnd C_bl
Cbb_40_80 bitb_40_80 gnd C_bl
Rb_40_81 bit_40_81 bit_40_82 R_bl
Rbb_40_81 bitb_40_81 bitb_40_82 R_bl
Cb_40_81 bit_40_81 gnd C_bl
Cbb_40_81 bitb_40_81 gnd C_bl
Rb_40_82 bit_40_82 bit_40_83 R_bl
Rbb_40_82 bitb_40_82 bitb_40_83 R_bl
Cb_40_82 bit_40_82 gnd C_bl
Cbb_40_82 bitb_40_82 gnd C_bl
Rb_40_83 bit_40_83 bit_40_84 R_bl
Rbb_40_83 bitb_40_83 bitb_40_84 R_bl
Cb_40_83 bit_40_83 gnd C_bl
Cbb_40_83 bitb_40_83 gnd C_bl
Rb_40_84 bit_40_84 bit_40_85 R_bl
Rbb_40_84 bitb_40_84 bitb_40_85 R_bl
Cb_40_84 bit_40_84 gnd C_bl
Cbb_40_84 bitb_40_84 gnd C_bl
Rb_40_85 bit_40_85 bit_40_86 R_bl
Rbb_40_85 bitb_40_85 bitb_40_86 R_bl
Cb_40_85 bit_40_85 gnd C_bl
Cbb_40_85 bitb_40_85 gnd C_bl
Rb_40_86 bit_40_86 bit_40_87 R_bl
Rbb_40_86 bitb_40_86 bitb_40_87 R_bl
Cb_40_86 bit_40_86 gnd C_bl
Cbb_40_86 bitb_40_86 gnd C_bl
Rb_40_87 bit_40_87 bit_40_88 R_bl
Rbb_40_87 bitb_40_87 bitb_40_88 R_bl
Cb_40_87 bit_40_87 gnd C_bl
Cbb_40_87 bitb_40_87 gnd C_bl
Rb_40_88 bit_40_88 bit_40_89 R_bl
Rbb_40_88 bitb_40_88 bitb_40_89 R_bl
Cb_40_88 bit_40_88 gnd C_bl
Cbb_40_88 bitb_40_88 gnd C_bl
Rb_40_89 bit_40_89 bit_40_90 R_bl
Rbb_40_89 bitb_40_89 bitb_40_90 R_bl
Cb_40_89 bit_40_89 gnd C_bl
Cbb_40_89 bitb_40_89 gnd C_bl
Rb_40_90 bit_40_90 bit_40_91 R_bl
Rbb_40_90 bitb_40_90 bitb_40_91 R_bl
Cb_40_90 bit_40_90 gnd C_bl
Cbb_40_90 bitb_40_90 gnd C_bl
Rb_40_91 bit_40_91 bit_40_92 R_bl
Rbb_40_91 bitb_40_91 bitb_40_92 R_bl
Cb_40_91 bit_40_91 gnd C_bl
Cbb_40_91 bitb_40_91 gnd C_bl
Rb_40_92 bit_40_92 bit_40_93 R_bl
Rbb_40_92 bitb_40_92 bitb_40_93 R_bl
Cb_40_92 bit_40_92 gnd C_bl
Cbb_40_92 bitb_40_92 gnd C_bl
Rb_40_93 bit_40_93 bit_40_94 R_bl
Rbb_40_93 bitb_40_93 bitb_40_94 R_bl
Cb_40_93 bit_40_93 gnd C_bl
Cbb_40_93 bitb_40_93 gnd C_bl
Rb_40_94 bit_40_94 bit_40_95 R_bl
Rbb_40_94 bitb_40_94 bitb_40_95 R_bl
Cb_40_94 bit_40_94 gnd C_bl
Cbb_40_94 bitb_40_94 gnd C_bl
Rb_40_95 bit_40_95 bit_40_96 R_bl
Rbb_40_95 bitb_40_95 bitb_40_96 R_bl
Cb_40_95 bit_40_95 gnd C_bl
Cbb_40_95 bitb_40_95 gnd C_bl
Rb_40_96 bit_40_96 bit_40_97 R_bl
Rbb_40_96 bitb_40_96 bitb_40_97 R_bl
Cb_40_96 bit_40_96 gnd C_bl
Cbb_40_96 bitb_40_96 gnd C_bl
Rb_40_97 bit_40_97 bit_40_98 R_bl
Rbb_40_97 bitb_40_97 bitb_40_98 R_bl
Cb_40_97 bit_40_97 gnd C_bl
Cbb_40_97 bitb_40_97 gnd C_bl
Rb_40_98 bit_40_98 bit_40_99 R_bl
Rbb_40_98 bitb_40_98 bitb_40_99 R_bl
Cb_40_98 bit_40_98 gnd C_bl
Cbb_40_98 bitb_40_98 gnd C_bl
Rb_40_99 bit_40_99 bit_40_100 R_bl
Rbb_40_99 bitb_40_99 bitb_40_100 R_bl
Cb_40_99 bit_40_99 gnd C_bl
Cbb_40_99 bitb_40_99 gnd C_bl
Rb_41_0 bit_41_0 bit_41_1 R_bl
Rbb_41_0 bitb_41_0 bitb_41_1 R_bl
Cb_41_0 bit_41_0 gnd C_bl
Cbb_41_0 bitb_41_0 gnd C_bl
Rb_41_1 bit_41_1 bit_41_2 R_bl
Rbb_41_1 bitb_41_1 bitb_41_2 R_bl
Cb_41_1 bit_41_1 gnd C_bl
Cbb_41_1 bitb_41_1 gnd C_bl
Rb_41_2 bit_41_2 bit_41_3 R_bl
Rbb_41_2 bitb_41_2 bitb_41_3 R_bl
Cb_41_2 bit_41_2 gnd C_bl
Cbb_41_2 bitb_41_2 gnd C_bl
Rb_41_3 bit_41_3 bit_41_4 R_bl
Rbb_41_3 bitb_41_3 bitb_41_4 R_bl
Cb_41_3 bit_41_3 gnd C_bl
Cbb_41_3 bitb_41_3 gnd C_bl
Rb_41_4 bit_41_4 bit_41_5 R_bl
Rbb_41_4 bitb_41_4 bitb_41_5 R_bl
Cb_41_4 bit_41_4 gnd C_bl
Cbb_41_4 bitb_41_4 gnd C_bl
Rb_41_5 bit_41_5 bit_41_6 R_bl
Rbb_41_5 bitb_41_5 bitb_41_6 R_bl
Cb_41_5 bit_41_5 gnd C_bl
Cbb_41_5 bitb_41_5 gnd C_bl
Rb_41_6 bit_41_6 bit_41_7 R_bl
Rbb_41_6 bitb_41_6 bitb_41_7 R_bl
Cb_41_6 bit_41_6 gnd C_bl
Cbb_41_6 bitb_41_6 gnd C_bl
Rb_41_7 bit_41_7 bit_41_8 R_bl
Rbb_41_7 bitb_41_7 bitb_41_8 R_bl
Cb_41_7 bit_41_7 gnd C_bl
Cbb_41_7 bitb_41_7 gnd C_bl
Rb_41_8 bit_41_8 bit_41_9 R_bl
Rbb_41_8 bitb_41_8 bitb_41_9 R_bl
Cb_41_8 bit_41_8 gnd C_bl
Cbb_41_8 bitb_41_8 gnd C_bl
Rb_41_9 bit_41_9 bit_41_10 R_bl
Rbb_41_9 bitb_41_9 bitb_41_10 R_bl
Cb_41_9 bit_41_9 gnd C_bl
Cbb_41_9 bitb_41_9 gnd C_bl
Rb_41_10 bit_41_10 bit_41_11 R_bl
Rbb_41_10 bitb_41_10 bitb_41_11 R_bl
Cb_41_10 bit_41_10 gnd C_bl
Cbb_41_10 bitb_41_10 gnd C_bl
Rb_41_11 bit_41_11 bit_41_12 R_bl
Rbb_41_11 bitb_41_11 bitb_41_12 R_bl
Cb_41_11 bit_41_11 gnd C_bl
Cbb_41_11 bitb_41_11 gnd C_bl
Rb_41_12 bit_41_12 bit_41_13 R_bl
Rbb_41_12 bitb_41_12 bitb_41_13 R_bl
Cb_41_12 bit_41_12 gnd C_bl
Cbb_41_12 bitb_41_12 gnd C_bl
Rb_41_13 bit_41_13 bit_41_14 R_bl
Rbb_41_13 bitb_41_13 bitb_41_14 R_bl
Cb_41_13 bit_41_13 gnd C_bl
Cbb_41_13 bitb_41_13 gnd C_bl
Rb_41_14 bit_41_14 bit_41_15 R_bl
Rbb_41_14 bitb_41_14 bitb_41_15 R_bl
Cb_41_14 bit_41_14 gnd C_bl
Cbb_41_14 bitb_41_14 gnd C_bl
Rb_41_15 bit_41_15 bit_41_16 R_bl
Rbb_41_15 bitb_41_15 bitb_41_16 R_bl
Cb_41_15 bit_41_15 gnd C_bl
Cbb_41_15 bitb_41_15 gnd C_bl
Rb_41_16 bit_41_16 bit_41_17 R_bl
Rbb_41_16 bitb_41_16 bitb_41_17 R_bl
Cb_41_16 bit_41_16 gnd C_bl
Cbb_41_16 bitb_41_16 gnd C_bl
Rb_41_17 bit_41_17 bit_41_18 R_bl
Rbb_41_17 bitb_41_17 bitb_41_18 R_bl
Cb_41_17 bit_41_17 gnd C_bl
Cbb_41_17 bitb_41_17 gnd C_bl
Rb_41_18 bit_41_18 bit_41_19 R_bl
Rbb_41_18 bitb_41_18 bitb_41_19 R_bl
Cb_41_18 bit_41_18 gnd C_bl
Cbb_41_18 bitb_41_18 gnd C_bl
Rb_41_19 bit_41_19 bit_41_20 R_bl
Rbb_41_19 bitb_41_19 bitb_41_20 R_bl
Cb_41_19 bit_41_19 gnd C_bl
Cbb_41_19 bitb_41_19 gnd C_bl
Rb_41_20 bit_41_20 bit_41_21 R_bl
Rbb_41_20 bitb_41_20 bitb_41_21 R_bl
Cb_41_20 bit_41_20 gnd C_bl
Cbb_41_20 bitb_41_20 gnd C_bl
Rb_41_21 bit_41_21 bit_41_22 R_bl
Rbb_41_21 bitb_41_21 bitb_41_22 R_bl
Cb_41_21 bit_41_21 gnd C_bl
Cbb_41_21 bitb_41_21 gnd C_bl
Rb_41_22 bit_41_22 bit_41_23 R_bl
Rbb_41_22 bitb_41_22 bitb_41_23 R_bl
Cb_41_22 bit_41_22 gnd C_bl
Cbb_41_22 bitb_41_22 gnd C_bl
Rb_41_23 bit_41_23 bit_41_24 R_bl
Rbb_41_23 bitb_41_23 bitb_41_24 R_bl
Cb_41_23 bit_41_23 gnd C_bl
Cbb_41_23 bitb_41_23 gnd C_bl
Rb_41_24 bit_41_24 bit_41_25 R_bl
Rbb_41_24 bitb_41_24 bitb_41_25 R_bl
Cb_41_24 bit_41_24 gnd C_bl
Cbb_41_24 bitb_41_24 gnd C_bl
Rb_41_25 bit_41_25 bit_41_26 R_bl
Rbb_41_25 bitb_41_25 bitb_41_26 R_bl
Cb_41_25 bit_41_25 gnd C_bl
Cbb_41_25 bitb_41_25 gnd C_bl
Rb_41_26 bit_41_26 bit_41_27 R_bl
Rbb_41_26 bitb_41_26 bitb_41_27 R_bl
Cb_41_26 bit_41_26 gnd C_bl
Cbb_41_26 bitb_41_26 gnd C_bl
Rb_41_27 bit_41_27 bit_41_28 R_bl
Rbb_41_27 bitb_41_27 bitb_41_28 R_bl
Cb_41_27 bit_41_27 gnd C_bl
Cbb_41_27 bitb_41_27 gnd C_bl
Rb_41_28 bit_41_28 bit_41_29 R_bl
Rbb_41_28 bitb_41_28 bitb_41_29 R_bl
Cb_41_28 bit_41_28 gnd C_bl
Cbb_41_28 bitb_41_28 gnd C_bl
Rb_41_29 bit_41_29 bit_41_30 R_bl
Rbb_41_29 bitb_41_29 bitb_41_30 R_bl
Cb_41_29 bit_41_29 gnd C_bl
Cbb_41_29 bitb_41_29 gnd C_bl
Rb_41_30 bit_41_30 bit_41_31 R_bl
Rbb_41_30 bitb_41_30 bitb_41_31 R_bl
Cb_41_30 bit_41_30 gnd C_bl
Cbb_41_30 bitb_41_30 gnd C_bl
Rb_41_31 bit_41_31 bit_41_32 R_bl
Rbb_41_31 bitb_41_31 bitb_41_32 R_bl
Cb_41_31 bit_41_31 gnd C_bl
Cbb_41_31 bitb_41_31 gnd C_bl
Rb_41_32 bit_41_32 bit_41_33 R_bl
Rbb_41_32 bitb_41_32 bitb_41_33 R_bl
Cb_41_32 bit_41_32 gnd C_bl
Cbb_41_32 bitb_41_32 gnd C_bl
Rb_41_33 bit_41_33 bit_41_34 R_bl
Rbb_41_33 bitb_41_33 bitb_41_34 R_bl
Cb_41_33 bit_41_33 gnd C_bl
Cbb_41_33 bitb_41_33 gnd C_bl
Rb_41_34 bit_41_34 bit_41_35 R_bl
Rbb_41_34 bitb_41_34 bitb_41_35 R_bl
Cb_41_34 bit_41_34 gnd C_bl
Cbb_41_34 bitb_41_34 gnd C_bl
Rb_41_35 bit_41_35 bit_41_36 R_bl
Rbb_41_35 bitb_41_35 bitb_41_36 R_bl
Cb_41_35 bit_41_35 gnd C_bl
Cbb_41_35 bitb_41_35 gnd C_bl
Rb_41_36 bit_41_36 bit_41_37 R_bl
Rbb_41_36 bitb_41_36 bitb_41_37 R_bl
Cb_41_36 bit_41_36 gnd C_bl
Cbb_41_36 bitb_41_36 gnd C_bl
Rb_41_37 bit_41_37 bit_41_38 R_bl
Rbb_41_37 bitb_41_37 bitb_41_38 R_bl
Cb_41_37 bit_41_37 gnd C_bl
Cbb_41_37 bitb_41_37 gnd C_bl
Rb_41_38 bit_41_38 bit_41_39 R_bl
Rbb_41_38 bitb_41_38 bitb_41_39 R_bl
Cb_41_38 bit_41_38 gnd C_bl
Cbb_41_38 bitb_41_38 gnd C_bl
Rb_41_39 bit_41_39 bit_41_40 R_bl
Rbb_41_39 bitb_41_39 bitb_41_40 R_bl
Cb_41_39 bit_41_39 gnd C_bl
Cbb_41_39 bitb_41_39 gnd C_bl
Rb_41_40 bit_41_40 bit_41_41 R_bl
Rbb_41_40 bitb_41_40 bitb_41_41 R_bl
Cb_41_40 bit_41_40 gnd C_bl
Cbb_41_40 bitb_41_40 gnd C_bl
Rb_41_41 bit_41_41 bit_41_42 R_bl
Rbb_41_41 bitb_41_41 bitb_41_42 R_bl
Cb_41_41 bit_41_41 gnd C_bl
Cbb_41_41 bitb_41_41 gnd C_bl
Rb_41_42 bit_41_42 bit_41_43 R_bl
Rbb_41_42 bitb_41_42 bitb_41_43 R_bl
Cb_41_42 bit_41_42 gnd C_bl
Cbb_41_42 bitb_41_42 gnd C_bl
Rb_41_43 bit_41_43 bit_41_44 R_bl
Rbb_41_43 bitb_41_43 bitb_41_44 R_bl
Cb_41_43 bit_41_43 gnd C_bl
Cbb_41_43 bitb_41_43 gnd C_bl
Rb_41_44 bit_41_44 bit_41_45 R_bl
Rbb_41_44 bitb_41_44 bitb_41_45 R_bl
Cb_41_44 bit_41_44 gnd C_bl
Cbb_41_44 bitb_41_44 gnd C_bl
Rb_41_45 bit_41_45 bit_41_46 R_bl
Rbb_41_45 bitb_41_45 bitb_41_46 R_bl
Cb_41_45 bit_41_45 gnd C_bl
Cbb_41_45 bitb_41_45 gnd C_bl
Rb_41_46 bit_41_46 bit_41_47 R_bl
Rbb_41_46 bitb_41_46 bitb_41_47 R_bl
Cb_41_46 bit_41_46 gnd C_bl
Cbb_41_46 bitb_41_46 gnd C_bl
Rb_41_47 bit_41_47 bit_41_48 R_bl
Rbb_41_47 bitb_41_47 bitb_41_48 R_bl
Cb_41_47 bit_41_47 gnd C_bl
Cbb_41_47 bitb_41_47 gnd C_bl
Rb_41_48 bit_41_48 bit_41_49 R_bl
Rbb_41_48 bitb_41_48 bitb_41_49 R_bl
Cb_41_48 bit_41_48 gnd C_bl
Cbb_41_48 bitb_41_48 gnd C_bl
Rb_41_49 bit_41_49 bit_41_50 R_bl
Rbb_41_49 bitb_41_49 bitb_41_50 R_bl
Cb_41_49 bit_41_49 gnd C_bl
Cbb_41_49 bitb_41_49 gnd C_bl
Rb_41_50 bit_41_50 bit_41_51 R_bl
Rbb_41_50 bitb_41_50 bitb_41_51 R_bl
Cb_41_50 bit_41_50 gnd C_bl
Cbb_41_50 bitb_41_50 gnd C_bl
Rb_41_51 bit_41_51 bit_41_52 R_bl
Rbb_41_51 bitb_41_51 bitb_41_52 R_bl
Cb_41_51 bit_41_51 gnd C_bl
Cbb_41_51 bitb_41_51 gnd C_bl
Rb_41_52 bit_41_52 bit_41_53 R_bl
Rbb_41_52 bitb_41_52 bitb_41_53 R_bl
Cb_41_52 bit_41_52 gnd C_bl
Cbb_41_52 bitb_41_52 gnd C_bl
Rb_41_53 bit_41_53 bit_41_54 R_bl
Rbb_41_53 bitb_41_53 bitb_41_54 R_bl
Cb_41_53 bit_41_53 gnd C_bl
Cbb_41_53 bitb_41_53 gnd C_bl
Rb_41_54 bit_41_54 bit_41_55 R_bl
Rbb_41_54 bitb_41_54 bitb_41_55 R_bl
Cb_41_54 bit_41_54 gnd C_bl
Cbb_41_54 bitb_41_54 gnd C_bl
Rb_41_55 bit_41_55 bit_41_56 R_bl
Rbb_41_55 bitb_41_55 bitb_41_56 R_bl
Cb_41_55 bit_41_55 gnd C_bl
Cbb_41_55 bitb_41_55 gnd C_bl
Rb_41_56 bit_41_56 bit_41_57 R_bl
Rbb_41_56 bitb_41_56 bitb_41_57 R_bl
Cb_41_56 bit_41_56 gnd C_bl
Cbb_41_56 bitb_41_56 gnd C_bl
Rb_41_57 bit_41_57 bit_41_58 R_bl
Rbb_41_57 bitb_41_57 bitb_41_58 R_bl
Cb_41_57 bit_41_57 gnd C_bl
Cbb_41_57 bitb_41_57 gnd C_bl
Rb_41_58 bit_41_58 bit_41_59 R_bl
Rbb_41_58 bitb_41_58 bitb_41_59 R_bl
Cb_41_58 bit_41_58 gnd C_bl
Cbb_41_58 bitb_41_58 gnd C_bl
Rb_41_59 bit_41_59 bit_41_60 R_bl
Rbb_41_59 bitb_41_59 bitb_41_60 R_bl
Cb_41_59 bit_41_59 gnd C_bl
Cbb_41_59 bitb_41_59 gnd C_bl
Rb_41_60 bit_41_60 bit_41_61 R_bl
Rbb_41_60 bitb_41_60 bitb_41_61 R_bl
Cb_41_60 bit_41_60 gnd C_bl
Cbb_41_60 bitb_41_60 gnd C_bl
Rb_41_61 bit_41_61 bit_41_62 R_bl
Rbb_41_61 bitb_41_61 bitb_41_62 R_bl
Cb_41_61 bit_41_61 gnd C_bl
Cbb_41_61 bitb_41_61 gnd C_bl
Rb_41_62 bit_41_62 bit_41_63 R_bl
Rbb_41_62 bitb_41_62 bitb_41_63 R_bl
Cb_41_62 bit_41_62 gnd C_bl
Cbb_41_62 bitb_41_62 gnd C_bl
Rb_41_63 bit_41_63 bit_41_64 R_bl
Rbb_41_63 bitb_41_63 bitb_41_64 R_bl
Cb_41_63 bit_41_63 gnd C_bl
Cbb_41_63 bitb_41_63 gnd C_bl
Rb_41_64 bit_41_64 bit_41_65 R_bl
Rbb_41_64 bitb_41_64 bitb_41_65 R_bl
Cb_41_64 bit_41_64 gnd C_bl
Cbb_41_64 bitb_41_64 gnd C_bl
Rb_41_65 bit_41_65 bit_41_66 R_bl
Rbb_41_65 bitb_41_65 bitb_41_66 R_bl
Cb_41_65 bit_41_65 gnd C_bl
Cbb_41_65 bitb_41_65 gnd C_bl
Rb_41_66 bit_41_66 bit_41_67 R_bl
Rbb_41_66 bitb_41_66 bitb_41_67 R_bl
Cb_41_66 bit_41_66 gnd C_bl
Cbb_41_66 bitb_41_66 gnd C_bl
Rb_41_67 bit_41_67 bit_41_68 R_bl
Rbb_41_67 bitb_41_67 bitb_41_68 R_bl
Cb_41_67 bit_41_67 gnd C_bl
Cbb_41_67 bitb_41_67 gnd C_bl
Rb_41_68 bit_41_68 bit_41_69 R_bl
Rbb_41_68 bitb_41_68 bitb_41_69 R_bl
Cb_41_68 bit_41_68 gnd C_bl
Cbb_41_68 bitb_41_68 gnd C_bl
Rb_41_69 bit_41_69 bit_41_70 R_bl
Rbb_41_69 bitb_41_69 bitb_41_70 R_bl
Cb_41_69 bit_41_69 gnd C_bl
Cbb_41_69 bitb_41_69 gnd C_bl
Rb_41_70 bit_41_70 bit_41_71 R_bl
Rbb_41_70 bitb_41_70 bitb_41_71 R_bl
Cb_41_70 bit_41_70 gnd C_bl
Cbb_41_70 bitb_41_70 gnd C_bl
Rb_41_71 bit_41_71 bit_41_72 R_bl
Rbb_41_71 bitb_41_71 bitb_41_72 R_bl
Cb_41_71 bit_41_71 gnd C_bl
Cbb_41_71 bitb_41_71 gnd C_bl
Rb_41_72 bit_41_72 bit_41_73 R_bl
Rbb_41_72 bitb_41_72 bitb_41_73 R_bl
Cb_41_72 bit_41_72 gnd C_bl
Cbb_41_72 bitb_41_72 gnd C_bl
Rb_41_73 bit_41_73 bit_41_74 R_bl
Rbb_41_73 bitb_41_73 bitb_41_74 R_bl
Cb_41_73 bit_41_73 gnd C_bl
Cbb_41_73 bitb_41_73 gnd C_bl
Rb_41_74 bit_41_74 bit_41_75 R_bl
Rbb_41_74 bitb_41_74 bitb_41_75 R_bl
Cb_41_74 bit_41_74 gnd C_bl
Cbb_41_74 bitb_41_74 gnd C_bl
Rb_41_75 bit_41_75 bit_41_76 R_bl
Rbb_41_75 bitb_41_75 bitb_41_76 R_bl
Cb_41_75 bit_41_75 gnd C_bl
Cbb_41_75 bitb_41_75 gnd C_bl
Rb_41_76 bit_41_76 bit_41_77 R_bl
Rbb_41_76 bitb_41_76 bitb_41_77 R_bl
Cb_41_76 bit_41_76 gnd C_bl
Cbb_41_76 bitb_41_76 gnd C_bl
Rb_41_77 bit_41_77 bit_41_78 R_bl
Rbb_41_77 bitb_41_77 bitb_41_78 R_bl
Cb_41_77 bit_41_77 gnd C_bl
Cbb_41_77 bitb_41_77 gnd C_bl
Rb_41_78 bit_41_78 bit_41_79 R_bl
Rbb_41_78 bitb_41_78 bitb_41_79 R_bl
Cb_41_78 bit_41_78 gnd C_bl
Cbb_41_78 bitb_41_78 gnd C_bl
Rb_41_79 bit_41_79 bit_41_80 R_bl
Rbb_41_79 bitb_41_79 bitb_41_80 R_bl
Cb_41_79 bit_41_79 gnd C_bl
Cbb_41_79 bitb_41_79 gnd C_bl
Rb_41_80 bit_41_80 bit_41_81 R_bl
Rbb_41_80 bitb_41_80 bitb_41_81 R_bl
Cb_41_80 bit_41_80 gnd C_bl
Cbb_41_80 bitb_41_80 gnd C_bl
Rb_41_81 bit_41_81 bit_41_82 R_bl
Rbb_41_81 bitb_41_81 bitb_41_82 R_bl
Cb_41_81 bit_41_81 gnd C_bl
Cbb_41_81 bitb_41_81 gnd C_bl
Rb_41_82 bit_41_82 bit_41_83 R_bl
Rbb_41_82 bitb_41_82 bitb_41_83 R_bl
Cb_41_82 bit_41_82 gnd C_bl
Cbb_41_82 bitb_41_82 gnd C_bl
Rb_41_83 bit_41_83 bit_41_84 R_bl
Rbb_41_83 bitb_41_83 bitb_41_84 R_bl
Cb_41_83 bit_41_83 gnd C_bl
Cbb_41_83 bitb_41_83 gnd C_bl
Rb_41_84 bit_41_84 bit_41_85 R_bl
Rbb_41_84 bitb_41_84 bitb_41_85 R_bl
Cb_41_84 bit_41_84 gnd C_bl
Cbb_41_84 bitb_41_84 gnd C_bl
Rb_41_85 bit_41_85 bit_41_86 R_bl
Rbb_41_85 bitb_41_85 bitb_41_86 R_bl
Cb_41_85 bit_41_85 gnd C_bl
Cbb_41_85 bitb_41_85 gnd C_bl
Rb_41_86 bit_41_86 bit_41_87 R_bl
Rbb_41_86 bitb_41_86 bitb_41_87 R_bl
Cb_41_86 bit_41_86 gnd C_bl
Cbb_41_86 bitb_41_86 gnd C_bl
Rb_41_87 bit_41_87 bit_41_88 R_bl
Rbb_41_87 bitb_41_87 bitb_41_88 R_bl
Cb_41_87 bit_41_87 gnd C_bl
Cbb_41_87 bitb_41_87 gnd C_bl
Rb_41_88 bit_41_88 bit_41_89 R_bl
Rbb_41_88 bitb_41_88 bitb_41_89 R_bl
Cb_41_88 bit_41_88 gnd C_bl
Cbb_41_88 bitb_41_88 gnd C_bl
Rb_41_89 bit_41_89 bit_41_90 R_bl
Rbb_41_89 bitb_41_89 bitb_41_90 R_bl
Cb_41_89 bit_41_89 gnd C_bl
Cbb_41_89 bitb_41_89 gnd C_bl
Rb_41_90 bit_41_90 bit_41_91 R_bl
Rbb_41_90 bitb_41_90 bitb_41_91 R_bl
Cb_41_90 bit_41_90 gnd C_bl
Cbb_41_90 bitb_41_90 gnd C_bl
Rb_41_91 bit_41_91 bit_41_92 R_bl
Rbb_41_91 bitb_41_91 bitb_41_92 R_bl
Cb_41_91 bit_41_91 gnd C_bl
Cbb_41_91 bitb_41_91 gnd C_bl
Rb_41_92 bit_41_92 bit_41_93 R_bl
Rbb_41_92 bitb_41_92 bitb_41_93 R_bl
Cb_41_92 bit_41_92 gnd C_bl
Cbb_41_92 bitb_41_92 gnd C_bl
Rb_41_93 bit_41_93 bit_41_94 R_bl
Rbb_41_93 bitb_41_93 bitb_41_94 R_bl
Cb_41_93 bit_41_93 gnd C_bl
Cbb_41_93 bitb_41_93 gnd C_bl
Rb_41_94 bit_41_94 bit_41_95 R_bl
Rbb_41_94 bitb_41_94 bitb_41_95 R_bl
Cb_41_94 bit_41_94 gnd C_bl
Cbb_41_94 bitb_41_94 gnd C_bl
Rb_41_95 bit_41_95 bit_41_96 R_bl
Rbb_41_95 bitb_41_95 bitb_41_96 R_bl
Cb_41_95 bit_41_95 gnd C_bl
Cbb_41_95 bitb_41_95 gnd C_bl
Rb_41_96 bit_41_96 bit_41_97 R_bl
Rbb_41_96 bitb_41_96 bitb_41_97 R_bl
Cb_41_96 bit_41_96 gnd C_bl
Cbb_41_96 bitb_41_96 gnd C_bl
Rb_41_97 bit_41_97 bit_41_98 R_bl
Rbb_41_97 bitb_41_97 bitb_41_98 R_bl
Cb_41_97 bit_41_97 gnd C_bl
Cbb_41_97 bitb_41_97 gnd C_bl
Rb_41_98 bit_41_98 bit_41_99 R_bl
Rbb_41_98 bitb_41_98 bitb_41_99 R_bl
Cb_41_98 bit_41_98 gnd C_bl
Cbb_41_98 bitb_41_98 gnd C_bl
Rb_41_99 bit_41_99 bit_41_100 R_bl
Rbb_41_99 bitb_41_99 bitb_41_100 R_bl
Cb_41_99 bit_41_99 gnd C_bl
Cbb_41_99 bitb_41_99 gnd C_bl
Rb_42_0 bit_42_0 bit_42_1 R_bl
Rbb_42_0 bitb_42_0 bitb_42_1 R_bl
Cb_42_0 bit_42_0 gnd C_bl
Cbb_42_0 bitb_42_0 gnd C_bl
Rb_42_1 bit_42_1 bit_42_2 R_bl
Rbb_42_1 bitb_42_1 bitb_42_2 R_bl
Cb_42_1 bit_42_1 gnd C_bl
Cbb_42_1 bitb_42_1 gnd C_bl
Rb_42_2 bit_42_2 bit_42_3 R_bl
Rbb_42_2 bitb_42_2 bitb_42_3 R_bl
Cb_42_2 bit_42_2 gnd C_bl
Cbb_42_2 bitb_42_2 gnd C_bl
Rb_42_3 bit_42_3 bit_42_4 R_bl
Rbb_42_3 bitb_42_3 bitb_42_4 R_bl
Cb_42_3 bit_42_3 gnd C_bl
Cbb_42_3 bitb_42_3 gnd C_bl
Rb_42_4 bit_42_4 bit_42_5 R_bl
Rbb_42_4 bitb_42_4 bitb_42_5 R_bl
Cb_42_4 bit_42_4 gnd C_bl
Cbb_42_4 bitb_42_4 gnd C_bl
Rb_42_5 bit_42_5 bit_42_6 R_bl
Rbb_42_5 bitb_42_5 bitb_42_6 R_bl
Cb_42_5 bit_42_5 gnd C_bl
Cbb_42_5 bitb_42_5 gnd C_bl
Rb_42_6 bit_42_6 bit_42_7 R_bl
Rbb_42_6 bitb_42_6 bitb_42_7 R_bl
Cb_42_6 bit_42_6 gnd C_bl
Cbb_42_6 bitb_42_6 gnd C_bl
Rb_42_7 bit_42_7 bit_42_8 R_bl
Rbb_42_7 bitb_42_7 bitb_42_8 R_bl
Cb_42_7 bit_42_7 gnd C_bl
Cbb_42_7 bitb_42_7 gnd C_bl
Rb_42_8 bit_42_8 bit_42_9 R_bl
Rbb_42_8 bitb_42_8 bitb_42_9 R_bl
Cb_42_8 bit_42_8 gnd C_bl
Cbb_42_8 bitb_42_8 gnd C_bl
Rb_42_9 bit_42_9 bit_42_10 R_bl
Rbb_42_9 bitb_42_9 bitb_42_10 R_bl
Cb_42_9 bit_42_9 gnd C_bl
Cbb_42_9 bitb_42_9 gnd C_bl
Rb_42_10 bit_42_10 bit_42_11 R_bl
Rbb_42_10 bitb_42_10 bitb_42_11 R_bl
Cb_42_10 bit_42_10 gnd C_bl
Cbb_42_10 bitb_42_10 gnd C_bl
Rb_42_11 bit_42_11 bit_42_12 R_bl
Rbb_42_11 bitb_42_11 bitb_42_12 R_bl
Cb_42_11 bit_42_11 gnd C_bl
Cbb_42_11 bitb_42_11 gnd C_bl
Rb_42_12 bit_42_12 bit_42_13 R_bl
Rbb_42_12 bitb_42_12 bitb_42_13 R_bl
Cb_42_12 bit_42_12 gnd C_bl
Cbb_42_12 bitb_42_12 gnd C_bl
Rb_42_13 bit_42_13 bit_42_14 R_bl
Rbb_42_13 bitb_42_13 bitb_42_14 R_bl
Cb_42_13 bit_42_13 gnd C_bl
Cbb_42_13 bitb_42_13 gnd C_bl
Rb_42_14 bit_42_14 bit_42_15 R_bl
Rbb_42_14 bitb_42_14 bitb_42_15 R_bl
Cb_42_14 bit_42_14 gnd C_bl
Cbb_42_14 bitb_42_14 gnd C_bl
Rb_42_15 bit_42_15 bit_42_16 R_bl
Rbb_42_15 bitb_42_15 bitb_42_16 R_bl
Cb_42_15 bit_42_15 gnd C_bl
Cbb_42_15 bitb_42_15 gnd C_bl
Rb_42_16 bit_42_16 bit_42_17 R_bl
Rbb_42_16 bitb_42_16 bitb_42_17 R_bl
Cb_42_16 bit_42_16 gnd C_bl
Cbb_42_16 bitb_42_16 gnd C_bl
Rb_42_17 bit_42_17 bit_42_18 R_bl
Rbb_42_17 bitb_42_17 bitb_42_18 R_bl
Cb_42_17 bit_42_17 gnd C_bl
Cbb_42_17 bitb_42_17 gnd C_bl
Rb_42_18 bit_42_18 bit_42_19 R_bl
Rbb_42_18 bitb_42_18 bitb_42_19 R_bl
Cb_42_18 bit_42_18 gnd C_bl
Cbb_42_18 bitb_42_18 gnd C_bl
Rb_42_19 bit_42_19 bit_42_20 R_bl
Rbb_42_19 bitb_42_19 bitb_42_20 R_bl
Cb_42_19 bit_42_19 gnd C_bl
Cbb_42_19 bitb_42_19 gnd C_bl
Rb_42_20 bit_42_20 bit_42_21 R_bl
Rbb_42_20 bitb_42_20 bitb_42_21 R_bl
Cb_42_20 bit_42_20 gnd C_bl
Cbb_42_20 bitb_42_20 gnd C_bl
Rb_42_21 bit_42_21 bit_42_22 R_bl
Rbb_42_21 bitb_42_21 bitb_42_22 R_bl
Cb_42_21 bit_42_21 gnd C_bl
Cbb_42_21 bitb_42_21 gnd C_bl
Rb_42_22 bit_42_22 bit_42_23 R_bl
Rbb_42_22 bitb_42_22 bitb_42_23 R_bl
Cb_42_22 bit_42_22 gnd C_bl
Cbb_42_22 bitb_42_22 gnd C_bl
Rb_42_23 bit_42_23 bit_42_24 R_bl
Rbb_42_23 bitb_42_23 bitb_42_24 R_bl
Cb_42_23 bit_42_23 gnd C_bl
Cbb_42_23 bitb_42_23 gnd C_bl
Rb_42_24 bit_42_24 bit_42_25 R_bl
Rbb_42_24 bitb_42_24 bitb_42_25 R_bl
Cb_42_24 bit_42_24 gnd C_bl
Cbb_42_24 bitb_42_24 gnd C_bl
Rb_42_25 bit_42_25 bit_42_26 R_bl
Rbb_42_25 bitb_42_25 bitb_42_26 R_bl
Cb_42_25 bit_42_25 gnd C_bl
Cbb_42_25 bitb_42_25 gnd C_bl
Rb_42_26 bit_42_26 bit_42_27 R_bl
Rbb_42_26 bitb_42_26 bitb_42_27 R_bl
Cb_42_26 bit_42_26 gnd C_bl
Cbb_42_26 bitb_42_26 gnd C_bl
Rb_42_27 bit_42_27 bit_42_28 R_bl
Rbb_42_27 bitb_42_27 bitb_42_28 R_bl
Cb_42_27 bit_42_27 gnd C_bl
Cbb_42_27 bitb_42_27 gnd C_bl
Rb_42_28 bit_42_28 bit_42_29 R_bl
Rbb_42_28 bitb_42_28 bitb_42_29 R_bl
Cb_42_28 bit_42_28 gnd C_bl
Cbb_42_28 bitb_42_28 gnd C_bl
Rb_42_29 bit_42_29 bit_42_30 R_bl
Rbb_42_29 bitb_42_29 bitb_42_30 R_bl
Cb_42_29 bit_42_29 gnd C_bl
Cbb_42_29 bitb_42_29 gnd C_bl
Rb_42_30 bit_42_30 bit_42_31 R_bl
Rbb_42_30 bitb_42_30 bitb_42_31 R_bl
Cb_42_30 bit_42_30 gnd C_bl
Cbb_42_30 bitb_42_30 gnd C_bl
Rb_42_31 bit_42_31 bit_42_32 R_bl
Rbb_42_31 bitb_42_31 bitb_42_32 R_bl
Cb_42_31 bit_42_31 gnd C_bl
Cbb_42_31 bitb_42_31 gnd C_bl
Rb_42_32 bit_42_32 bit_42_33 R_bl
Rbb_42_32 bitb_42_32 bitb_42_33 R_bl
Cb_42_32 bit_42_32 gnd C_bl
Cbb_42_32 bitb_42_32 gnd C_bl
Rb_42_33 bit_42_33 bit_42_34 R_bl
Rbb_42_33 bitb_42_33 bitb_42_34 R_bl
Cb_42_33 bit_42_33 gnd C_bl
Cbb_42_33 bitb_42_33 gnd C_bl
Rb_42_34 bit_42_34 bit_42_35 R_bl
Rbb_42_34 bitb_42_34 bitb_42_35 R_bl
Cb_42_34 bit_42_34 gnd C_bl
Cbb_42_34 bitb_42_34 gnd C_bl
Rb_42_35 bit_42_35 bit_42_36 R_bl
Rbb_42_35 bitb_42_35 bitb_42_36 R_bl
Cb_42_35 bit_42_35 gnd C_bl
Cbb_42_35 bitb_42_35 gnd C_bl
Rb_42_36 bit_42_36 bit_42_37 R_bl
Rbb_42_36 bitb_42_36 bitb_42_37 R_bl
Cb_42_36 bit_42_36 gnd C_bl
Cbb_42_36 bitb_42_36 gnd C_bl
Rb_42_37 bit_42_37 bit_42_38 R_bl
Rbb_42_37 bitb_42_37 bitb_42_38 R_bl
Cb_42_37 bit_42_37 gnd C_bl
Cbb_42_37 bitb_42_37 gnd C_bl
Rb_42_38 bit_42_38 bit_42_39 R_bl
Rbb_42_38 bitb_42_38 bitb_42_39 R_bl
Cb_42_38 bit_42_38 gnd C_bl
Cbb_42_38 bitb_42_38 gnd C_bl
Rb_42_39 bit_42_39 bit_42_40 R_bl
Rbb_42_39 bitb_42_39 bitb_42_40 R_bl
Cb_42_39 bit_42_39 gnd C_bl
Cbb_42_39 bitb_42_39 gnd C_bl
Rb_42_40 bit_42_40 bit_42_41 R_bl
Rbb_42_40 bitb_42_40 bitb_42_41 R_bl
Cb_42_40 bit_42_40 gnd C_bl
Cbb_42_40 bitb_42_40 gnd C_bl
Rb_42_41 bit_42_41 bit_42_42 R_bl
Rbb_42_41 bitb_42_41 bitb_42_42 R_bl
Cb_42_41 bit_42_41 gnd C_bl
Cbb_42_41 bitb_42_41 gnd C_bl
Rb_42_42 bit_42_42 bit_42_43 R_bl
Rbb_42_42 bitb_42_42 bitb_42_43 R_bl
Cb_42_42 bit_42_42 gnd C_bl
Cbb_42_42 bitb_42_42 gnd C_bl
Rb_42_43 bit_42_43 bit_42_44 R_bl
Rbb_42_43 bitb_42_43 bitb_42_44 R_bl
Cb_42_43 bit_42_43 gnd C_bl
Cbb_42_43 bitb_42_43 gnd C_bl
Rb_42_44 bit_42_44 bit_42_45 R_bl
Rbb_42_44 bitb_42_44 bitb_42_45 R_bl
Cb_42_44 bit_42_44 gnd C_bl
Cbb_42_44 bitb_42_44 gnd C_bl
Rb_42_45 bit_42_45 bit_42_46 R_bl
Rbb_42_45 bitb_42_45 bitb_42_46 R_bl
Cb_42_45 bit_42_45 gnd C_bl
Cbb_42_45 bitb_42_45 gnd C_bl
Rb_42_46 bit_42_46 bit_42_47 R_bl
Rbb_42_46 bitb_42_46 bitb_42_47 R_bl
Cb_42_46 bit_42_46 gnd C_bl
Cbb_42_46 bitb_42_46 gnd C_bl
Rb_42_47 bit_42_47 bit_42_48 R_bl
Rbb_42_47 bitb_42_47 bitb_42_48 R_bl
Cb_42_47 bit_42_47 gnd C_bl
Cbb_42_47 bitb_42_47 gnd C_bl
Rb_42_48 bit_42_48 bit_42_49 R_bl
Rbb_42_48 bitb_42_48 bitb_42_49 R_bl
Cb_42_48 bit_42_48 gnd C_bl
Cbb_42_48 bitb_42_48 gnd C_bl
Rb_42_49 bit_42_49 bit_42_50 R_bl
Rbb_42_49 bitb_42_49 bitb_42_50 R_bl
Cb_42_49 bit_42_49 gnd C_bl
Cbb_42_49 bitb_42_49 gnd C_bl
Rb_42_50 bit_42_50 bit_42_51 R_bl
Rbb_42_50 bitb_42_50 bitb_42_51 R_bl
Cb_42_50 bit_42_50 gnd C_bl
Cbb_42_50 bitb_42_50 gnd C_bl
Rb_42_51 bit_42_51 bit_42_52 R_bl
Rbb_42_51 bitb_42_51 bitb_42_52 R_bl
Cb_42_51 bit_42_51 gnd C_bl
Cbb_42_51 bitb_42_51 gnd C_bl
Rb_42_52 bit_42_52 bit_42_53 R_bl
Rbb_42_52 bitb_42_52 bitb_42_53 R_bl
Cb_42_52 bit_42_52 gnd C_bl
Cbb_42_52 bitb_42_52 gnd C_bl
Rb_42_53 bit_42_53 bit_42_54 R_bl
Rbb_42_53 bitb_42_53 bitb_42_54 R_bl
Cb_42_53 bit_42_53 gnd C_bl
Cbb_42_53 bitb_42_53 gnd C_bl
Rb_42_54 bit_42_54 bit_42_55 R_bl
Rbb_42_54 bitb_42_54 bitb_42_55 R_bl
Cb_42_54 bit_42_54 gnd C_bl
Cbb_42_54 bitb_42_54 gnd C_bl
Rb_42_55 bit_42_55 bit_42_56 R_bl
Rbb_42_55 bitb_42_55 bitb_42_56 R_bl
Cb_42_55 bit_42_55 gnd C_bl
Cbb_42_55 bitb_42_55 gnd C_bl
Rb_42_56 bit_42_56 bit_42_57 R_bl
Rbb_42_56 bitb_42_56 bitb_42_57 R_bl
Cb_42_56 bit_42_56 gnd C_bl
Cbb_42_56 bitb_42_56 gnd C_bl
Rb_42_57 bit_42_57 bit_42_58 R_bl
Rbb_42_57 bitb_42_57 bitb_42_58 R_bl
Cb_42_57 bit_42_57 gnd C_bl
Cbb_42_57 bitb_42_57 gnd C_bl
Rb_42_58 bit_42_58 bit_42_59 R_bl
Rbb_42_58 bitb_42_58 bitb_42_59 R_bl
Cb_42_58 bit_42_58 gnd C_bl
Cbb_42_58 bitb_42_58 gnd C_bl
Rb_42_59 bit_42_59 bit_42_60 R_bl
Rbb_42_59 bitb_42_59 bitb_42_60 R_bl
Cb_42_59 bit_42_59 gnd C_bl
Cbb_42_59 bitb_42_59 gnd C_bl
Rb_42_60 bit_42_60 bit_42_61 R_bl
Rbb_42_60 bitb_42_60 bitb_42_61 R_bl
Cb_42_60 bit_42_60 gnd C_bl
Cbb_42_60 bitb_42_60 gnd C_bl
Rb_42_61 bit_42_61 bit_42_62 R_bl
Rbb_42_61 bitb_42_61 bitb_42_62 R_bl
Cb_42_61 bit_42_61 gnd C_bl
Cbb_42_61 bitb_42_61 gnd C_bl
Rb_42_62 bit_42_62 bit_42_63 R_bl
Rbb_42_62 bitb_42_62 bitb_42_63 R_bl
Cb_42_62 bit_42_62 gnd C_bl
Cbb_42_62 bitb_42_62 gnd C_bl
Rb_42_63 bit_42_63 bit_42_64 R_bl
Rbb_42_63 bitb_42_63 bitb_42_64 R_bl
Cb_42_63 bit_42_63 gnd C_bl
Cbb_42_63 bitb_42_63 gnd C_bl
Rb_42_64 bit_42_64 bit_42_65 R_bl
Rbb_42_64 bitb_42_64 bitb_42_65 R_bl
Cb_42_64 bit_42_64 gnd C_bl
Cbb_42_64 bitb_42_64 gnd C_bl
Rb_42_65 bit_42_65 bit_42_66 R_bl
Rbb_42_65 bitb_42_65 bitb_42_66 R_bl
Cb_42_65 bit_42_65 gnd C_bl
Cbb_42_65 bitb_42_65 gnd C_bl
Rb_42_66 bit_42_66 bit_42_67 R_bl
Rbb_42_66 bitb_42_66 bitb_42_67 R_bl
Cb_42_66 bit_42_66 gnd C_bl
Cbb_42_66 bitb_42_66 gnd C_bl
Rb_42_67 bit_42_67 bit_42_68 R_bl
Rbb_42_67 bitb_42_67 bitb_42_68 R_bl
Cb_42_67 bit_42_67 gnd C_bl
Cbb_42_67 bitb_42_67 gnd C_bl
Rb_42_68 bit_42_68 bit_42_69 R_bl
Rbb_42_68 bitb_42_68 bitb_42_69 R_bl
Cb_42_68 bit_42_68 gnd C_bl
Cbb_42_68 bitb_42_68 gnd C_bl
Rb_42_69 bit_42_69 bit_42_70 R_bl
Rbb_42_69 bitb_42_69 bitb_42_70 R_bl
Cb_42_69 bit_42_69 gnd C_bl
Cbb_42_69 bitb_42_69 gnd C_bl
Rb_42_70 bit_42_70 bit_42_71 R_bl
Rbb_42_70 bitb_42_70 bitb_42_71 R_bl
Cb_42_70 bit_42_70 gnd C_bl
Cbb_42_70 bitb_42_70 gnd C_bl
Rb_42_71 bit_42_71 bit_42_72 R_bl
Rbb_42_71 bitb_42_71 bitb_42_72 R_bl
Cb_42_71 bit_42_71 gnd C_bl
Cbb_42_71 bitb_42_71 gnd C_bl
Rb_42_72 bit_42_72 bit_42_73 R_bl
Rbb_42_72 bitb_42_72 bitb_42_73 R_bl
Cb_42_72 bit_42_72 gnd C_bl
Cbb_42_72 bitb_42_72 gnd C_bl
Rb_42_73 bit_42_73 bit_42_74 R_bl
Rbb_42_73 bitb_42_73 bitb_42_74 R_bl
Cb_42_73 bit_42_73 gnd C_bl
Cbb_42_73 bitb_42_73 gnd C_bl
Rb_42_74 bit_42_74 bit_42_75 R_bl
Rbb_42_74 bitb_42_74 bitb_42_75 R_bl
Cb_42_74 bit_42_74 gnd C_bl
Cbb_42_74 bitb_42_74 gnd C_bl
Rb_42_75 bit_42_75 bit_42_76 R_bl
Rbb_42_75 bitb_42_75 bitb_42_76 R_bl
Cb_42_75 bit_42_75 gnd C_bl
Cbb_42_75 bitb_42_75 gnd C_bl
Rb_42_76 bit_42_76 bit_42_77 R_bl
Rbb_42_76 bitb_42_76 bitb_42_77 R_bl
Cb_42_76 bit_42_76 gnd C_bl
Cbb_42_76 bitb_42_76 gnd C_bl
Rb_42_77 bit_42_77 bit_42_78 R_bl
Rbb_42_77 bitb_42_77 bitb_42_78 R_bl
Cb_42_77 bit_42_77 gnd C_bl
Cbb_42_77 bitb_42_77 gnd C_bl
Rb_42_78 bit_42_78 bit_42_79 R_bl
Rbb_42_78 bitb_42_78 bitb_42_79 R_bl
Cb_42_78 bit_42_78 gnd C_bl
Cbb_42_78 bitb_42_78 gnd C_bl
Rb_42_79 bit_42_79 bit_42_80 R_bl
Rbb_42_79 bitb_42_79 bitb_42_80 R_bl
Cb_42_79 bit_42_79 gnd C_bl
Cbb_42_79 bitb_42_79 gnd C_bl
Rb_42_80 bit_42_80 bit_42_81 R_bl
Rbb_42_80 bitb_42_80 bitb_42_81 R_bl
Cb_42_80 bit_42_80 gnd C_bl
Cbb_42_80 bitb_42_80 gnd C_bl
Rb_42_81 bit_42_81 bit_42_82 R_bl
Rbb_42_81 bitb_42_81 bitb_42_82 R_bl
Cb_42_81 bit_42_81 gnd C_bl
Cbb_42_81 bitb_42_81 gnd C_bl
Rb_42_82 bit_42_82 bit_42_83 R_bl
Rbb_42_82 bitb_42_82 bitb_42_83 R_bl
Cb_42_82 bit_42_82 gnd C_bl
Cbb_42_82 bitb_42_82 gnd C_bl
Rb_42_83 bit_42_83 bit_42_84 R_bl
Rbb_42_83 bitb_42_83 bitb_42_84 R_bl
Cb_42_83 bit_42_83 gnd C_bl
Cbb_42_83 bitb_42_83 gnd C_bl
Rb_42_84 bit_42_84 bit_42_85 R_bl
Rbb_42_84 bitb_42_84 bitb_42_85 R_bl
Cb_42_84 bit_42_84 gnd C_bl
Cbb_42_84 bitb_42_84 gnd C_bl
Rb_42_85 bit_42_85 bit_42_86 R_bl
Rbb_42_85 bitb_42_85 bitb_42_86 R_bl
Cb_42_85 bit_42_85 gnd C_bl
Cbb_42_85 bitb_42_85 gnd C_bl
Rb_42_86 bit_42_86 bit_42_87 R_bl
Rbb_42_86 bitb_42_86 bitb_42_87 R_bl
Cb_42_86 bit_42_86 gnd C_bl
Cbb_42_86 bitb_42_86 gnd C_bl
Rb_42_87 bit_42_87 bit_42_88 R_bl
Rbb_42_87 bitb_42_87 bitb_42_88 R_bl
Cb_42_87 bit_42_87 gnd C_bl
Cbb_42_87 bitb_42_87 gnd C_bl
Rb_42_88 bit_42_88 bit_42_89 R_bl
Rbb_42_88 bitb_42_88 bitb_42_89 R_bl
Cb_42_88 bit_42_88 gnd C_bl
Cbb_42_88 bitb_42_88 gnd C_bl
Rb_42_89 bit_42_89 bit_42_90 R_bl
Rbb_42_89 bitb_42_89 bitb_42_90 R_bl
Cb_42_89 bit_42_89 gnd C_bl
Cbb_42_89 bitb_42_89 gnd C_bl
Rb_42_90 bit_42_90 bit_42_91 R_bl
Rbb_42_90 bitb_42_90 bitb_42_91 R_bl
Cb_42_90 bit_42_90 gnd C_bl
Cbb_42_90 bitb_42_90 gnd C_bl
Rb_42_91 bit_42_91 bit_42_92 R_bl
Rbb_42_91 bitb_42_91 bitb_42_92 R_bl
Cb_42_91 bit_42_91 gnd C_bl
Cbb_42_91 bitb_42_91 gnd C_bl
Rb_42_92 bit_42_92 bit_42_93 R_bl
Rbb_42_92 bitb_42_92 bitb_42_93 R_bl
Cb_42_92 bit_42_92 gnd C_bl
Cbb_42_92 bitb_42_92 gnd C_bl
Rb_42_93 bit_42_93 bit_42_94 R_bl
Rbb_42_93 bitb_42_93 bitb_42_94 R_bl
Cb_42_93 bit_42_93 gnd C_bl
Cbb_42_93 bitb_42_93 gnd C_bl
Rb_42_94 bit_42_94 bit_42_95 R_bl
Rbb_42_94 bitb_42_94 bitb_42_95 R_bl
Cb_42_94 bit_42_94 gnd C_bl
Cbb_42_94 bitb_42_94 gnd C_bl
Rb_42_95 bit_42_95 bit_42_96 R_bl
Rbb_42_95 bitb_42_95 bitb_42_96 R_bl
Cb_42_95 bit_42_95 gnd C_bl
Cbb_42_95 bitb_42_95 gnd C_bl
Rb_42_96 bit_42_96 bit_42_97 R_bl
Rbb_42_96 bitb_42_96 bitb_42_97 R_bl
Cb_42_96 bit_42_96 gnd C_bl
Cbb_42_96 bitb_42_96 gnd C_bl
Rb_42_97 bit_42_97 bit_42_98 R_bl
Rbb_42_97 bitb_42_97 bitb_42_98 R_bl
Cb_42_97 bit_42_97 gnd C_bl
Cbb_42_97 bitb_42_97 gnd C_bl
Rb_42_98 bit_42_98 bit_42_99 R_bl
Rbb_42_98 bitb_42_98 bitb_42_99 R_bl
Cb_42_98 bit_42_98 gnd C_bl
Cbb_42_98 bitb_42_98 gnd C_bl
Rb_42_99 bit_42_99 bit_42_100 R_bl
Rbb_42_99 bitb_42_99 bitb_42_100 R_bl
Cb_42_99 bit_42_99 gnd C_bl
Cbb_42_99 bitb_42_99 gnd C_bl
Rb_43_0 bit_43_0 bit_43_1 R_bl
Rbb_43_0 bitb_43_0 bitb_43_1 R_bl
Cb_43_0 bit_43_0 gnd C_bl
Cbb_43_0 bitb_43_0 gnd C_bl
Rb_43_1 bit_43_1 bit_43_2 R_bl
Rbb_43_1 bitb_43_1 bitb_43_2 R_bl
Cb_43_1 bit_43_1 gnd C_bl
Cbb_43_1 bitb_43_1 gnd C_bl
Rb_43_2 bit_43_2 bit_43_3 R_bl
Rbb_43_2 bitb_43_2 bitb_43_3 R_bl
Cb_43_2 bit_43_2 gnd C_bl
Cbb_43_2 bitb_43_2 gnd C_bl
Rb_43_3 bit_43_3 bit_43_4 R_bl
Rbb_43_3 bitb_43_3 bitb_43_4 R_bl
Cb_43_3 bit_43_3 gnd C_bl
Cbb_43_3 bitb_43_3 gnd C_bl
Rb_43_4 bit_43_4 bit_43_5 R_bl
Rbb_43_4 bitb_43_4 bitb_43_5 R_bl
Cb_43_4 bit_43_4 gnd C_bl
Cbb_43_4 bitb_43_4 gnd C_bl
Rb_43_5 bit_43_5 bit_43_6 R_bl
Rbb_43_5 bitb_43_5 bitb_43_6 R_bl
Cb_43_5 bit_43_5 gnd C_bl
Cbb_43_5 bitb_43_5 gnd C_bl
Rb_43_6 bit_43_6 bit_43_7 R_bl
Rbb_43_6 bitb_43_6 bitb_43_7 R_bl
Cb_43_6 bit_43_6 gnd C_bl
Cbb_43_6 bitb_43_6 gnd C_bl
Rb_43_7 bit_43_7 bit_43_8 R_bl
Rbb_43_7 bitb_43_7 bitb_43_8 R_bl
Cb_43_7 bit_43_7 gnd C_bl
Cbb_43_7 bitb_43_7 gnd C_bl
Rb_43_8 bit_43_8 bit_43_9 R_bl
Rbb_43_8 bitb_43_8 bitb_43_9 R_bl
Cb_43_8 bit_43_8 gnd C_bl
Cbb_43_8 bitb_43_8 gnd C_bl
Rb_43_9 bit_43_9 bit_43_10 R_bl
Rbb_43_9 bitb_43_9 bitb_43_10 R_bl
Cb_43_9 bit_43_9 gnd C_bl
Cbb_43_9 bitb_43_9 gnd C_bl
Rb_43_10 bit_43_10 bit_43_11 R_bl
Rbb_43_10 bitb_43_10 bitb_43_11 R_bl
Cb_43_10 bit_43_10 gnd C_bl
Cbb_43_10 bitb_43_10 gnd C_bl
Rb_43_11 bit_43_11 bit_43_12 R_bl
Rbb_43_11 bitb_43_11 bitb_43_12 R_bl
Cb_43_11 bit_43_11 gnd C_bl
Cbb_43_11 bitb_43_11 gnd C_bl
Rb_43_12 bit_43_12 bit_43_13 R_bl
Rbb_43_12 bitb_43_12 bitb_43_13 R_bl
Cb_43_12 bit_43_12 gnd C_bl
Cbb_43_12 bitb_43_12 gnd C_bl
Rb_43_13 bit_43_13 bit_43_14 R_bl
Rbb_43_13 bitb_43_13 bitb_43_14 R_bl
Cb_43_13 bit_43_13 gnd C_bl
Cbb_43_13 bitb_43_13 gnd C_bl
Rb_43_14 bit_43_14 bit_43_15 R_bl
Rbb_43_14 bitb_43_14 bitb_43_15 R_bl
Cb_43_14 bit_43_14 gnd C_bl
Cbb_43_14 bitb_43_14 gnd C_bl
Rb_43_15 bit_43_15 bit_43_16 R_bl
Rbb_43_15 bitb_43_15 bitb_43_16 R_bl
Cb_43_15 bit_43_15 gnd C_bl
Cbb_43_15 bitb_43_15 gnd C_bl
Rb_43_16 bit_43_16 bit_43_17 R_bl
Rbb_43_16 bitb_43_16 bitb_43_17 R_bl
Cb_43_16 bit_43_16 gnd C_bl
Cbb_43_16 bitb_43_16 gnd C_bl
Rb_43_17 bit_43_17 bit_43_18 R_bl
Rbb_43_17 bitb_43_17 bitb_43_18 R_bl
Cb_43_17 bit_43_17 gnd C_bl
Cbb_43_17 bitb_43_17 gnd C_bl
Rb_43_18 bit_43_18 bit_43_19 R_bl
Rbb_43_18 bitb_43_18 bitb_43_19 R_bl
Cb_43_18 bit_43_18 gnd C_bl
Cbb_43_18 bitb_43_18 gnd C_bl
Rb_43_19 bit_43_19 bit_43_20 R_bl
Rbb_43_19 bitb_43_19 bitb_43_20 R_bl
Cb_43_19 bit_43_19 gnd C_bl
Cbb_43_19 bitb_43_19 gnd C_bl
Rb_43_20 bit_43_20 bit_43_21 R_bl
Rbb_43_20 bitb_43_20 bitb_43_21 R_bl
Cb_43_20 bit_43_20 gnd C_bl
Cbb_43_20 bitb_43_20 gnd C_bl
Rb_43_21 bit_43_21 bit_43_22 R_bl
Rbb_43_21 bitb_43_21 bitb_43_22 R_bl
Cb_43_21 bit_43_21 gnd C_bl
Cbb_43_21 bitb_43_21 gnd C_bl
Rb_43_22 bit_43_22 bit_43_23 R_bl
Rbb_43_22 bitb_43_22 bitb_43_23 R_bl
Cb_43_22 bit_43_22 gnd C_bl
Cbb_43_22 bitb_43_22 gnd C_bl
Rb_43_23 bit_43_23 bit_43_24 R_bl
Rbb_43_23 bitb_43_23 bitb_43_24 R_bl
Cb_43_23 bit_43_23 gnd C_bl
Cbb_43_23 bitb_43_23 gnd C_bl
Rb_43_24 bit_43_24 bit_43_25 R_bl
Rbb_43_24 bitb_43_24 bitb_43_25 R_bl
Cb_43_24 bit_43_24 gnd C_bl
Cbb_43_24 bitb_43_24 gnd C_bl
Rb_43_25 bit_43_25 bit_43_26 R_bl
Rbb_43_25 bitb_43_25 bitb_43_26 R_bl
Cb_43_25 bit_43_25 gnd C_bl
Cbb_43_25 bitb_43_25 gnd C_bl
Rb_43_26 bit_43_26 bit_43_27 R_bl
Rbb_43_26 bitb_43_26 bitb_43_27 R_bl
Cb_43_26 bit_43_26 gnd C_bl
Cbb_43_26 bitb_43_26 gnd C_bl
Rb_43_27 bit_43_27 bit_43_28 R_bl
Rbb_43_27 bitb_43_27 bitb_43_28 R_bl
Cb_43_27 bit_43_27 gnd C_bl
Cbb_43_27 bitb_43_27 gnd C_bl
Rb_43_28 bit_43_28 bit_43_29 R_bl
Rbb_43_28 bitb_43_28 bitb_43_29 R_bl
Cb_43_28 bit_43_28 gnd C_bl
Cbb_43_28 bitb_43_28 gnd C_bl
Rb_43_29 bit_43_29 bit_43_30 R_bl
Rbb_43_29 bitb_43_29 bitb_43_30 R_bl
Cb_43_29 bit_43_29 gnd C_bl
Cbb_43_29 bitb_43_29 gnd C_bl
Rb_43_30 bit_43_30 bit_43_31 R_bl
Rbb_43_30 bitb_43_30 bitb_43_31 R_bl
Cb_43_30 bit_43_30 gnd C_bl
Cbb_43_30 bitb_43_30 gnd C_bl
Rb_43_31 bit_43_31 bit_43_32 R_bl
Rbb_43_31 bitb_43_31 bitb_43_32 R_bl
Cb_43_31 bit_43_31 gnd C_bl
Cbb_43_31 bitb_43_31 gnd C_bl
Rb_43_32 bit_43_32 bit_43_33 R_bl
Rbb_43_32 bitb_43_32 bitb_43_33 R_bl
Cb_43_32 bit_43_32 gnd C_bl
Cbb_43_32 bitb_43_32 gnd C_bl
Rb_43_33 bit_43_33 bit_43_34 R_bl
Rbb_43_33 bitb_43_33 bitb_43_34 R_bl
Cb_43_33 bit_43_33 gnd C_bl
Cbb_43_33 bitb_43_33 gnd C_bl
Rb_43_34 bit_43_34 bit_43_35 R_bl
Rbb_43_34 bitb_43_34 bitb_43_35 R_bl
Cb_43_34 bit_43_34 gnd C_bl
Cbb_43_34 bitb_43_34 gnd C_bl
Rb_43_35 bit_43_35 bit_43_36 R_bl
Rbb_43_35 bitb_43_35 bitb_43_36 R_bl
Cb_43_35 bit_43_35 gnd C_bl
Cbb_43_35 bitb_43_35 gnd C_bl
Rb_43_36 bit_43_36 bit_43_37 R_bl
Rbb_43_36 bitb_43_36 bitb_43_37 R_bl
Cb_43_36 bit_43_36 gnd C_bl
Cbb_43_36 bitb_43_36 gnd C_bl
Rb_43_37 bit_43_37 bit_43_38 R_bl
Rbb_43_37 bitb_43_37 bitb_43_38 R_bl
Cb_43_37 bit_43_37 gnd C_bl
Cbb_43_37 bitb_43_37 gnd C_bl
Rb_43_38 bit_43_38 bit_43_39 R_bl
Rbb_43_38 bitb_43_38 bitb_43_39 R_bl
Cb_43_38 bit_43_38 gnd C_bl
Cbb_43_38 bitb_43_38 gnd C_bl
Rb_43_39 bit_43_39 bit_43_40 R_bl
Rbb_43_39 bitb_43_39 bitb_43_40 R_bl
Cb_43_39 bit_43_39 gnd C_bl
Cbb_43_39 bitb_43_39 gnd C_bl
Rb_43_40 bit_43_40 bit_43_41 R_bl
Rbb_43_40 bitb_43_40 bitb_43_41 R_bl
Cb_43_40 bit_43_40 gnd C_bl
Cbb_43_40 bitb_43_40 gnd C_bl
Rb_43_41 bit_43_41 bit_43_42 R_bl
Rbb_43_41 bitb_43_41 bitb_43_42 R_bl
Cb_43_41 bit_43_41 gnd C_bl
Cbb_43_41 bitb_43_41 gnd C_bl
Rb_43_42 bit_43_42 bit_43_43 R_bl
Rbb_43_42 bitb_43_42 bitb_43_43 R_bl
Cb_43_42 bit_43_42 gnd C_bl
Cbb_43_42 bitb_43_42 gnd C_bl
Rb_43_43 bit_43_43 bit_43_44 R_bl
Rbb_43_43 bitb_43_43 bitb_43_44 R_bl
Cb_43_43 bit_43_43 gnd C_bl
Cbb_43_43 bitb_43_43 gnd C_bl
Rb_43_44 bit_43_44 bit_43_45 R_bl
Rbb_43_44 bitb_43_44 bitb_43_45 R_bl
Cb_43_44 bit_43_44 gnd C_bl
Cbb_43_44 bitb_43_44 gnd C_bl
Rb_43_45 bit_43_45 bit_43_46 R_bl
Rbb_43_45 bitb_43_45 bitb_43_46 R_bl
Cb_43_45 bit_43_45 gnd C_bl
Cbb_43_45 bitb_43_45 gnd C_bl
Rb_43_46 bit_43_46 bit_43_47 R_bl
Rbb_43_46 bitb_43_46 bitb_43_47 R_bl
Cb_43_46 bit_43_46 gnd C_bl
Cbb_43_46 bitb_43_46 gnd C_bl
Rb_43_47 bit_43_47 bit_43_48 R_bl
Rbb_43_47 bitb_43_47 bitb_43_48 R_bl
Cb_43_47 bit_43_47 gnd C_bl
Cbb_43_47 bitb_43_47 gnd C_bl
Rb_43_48 bit_43_48 bit_43_49 R_bl
Rbb_43_48 bitb_43_48 bitb_43_49 R_bl
Cb_43_48 bit_43_48 gnd C_bl
Cbb_43_48 bitb_43_48 gnd C_bl
Rb_43_49 bit_43_49 bit_43_50 R_bl
Rbb_43_49 bitb_43_49 bitb_43_50 R_bl
Cb_43_49 bit_43_49 gnd C_bl
Cbb_43_49 bitb_43_49 gnd C_bl
Rb_43_50 bit_43_50 bit_43_51 R_bl
Rbb_43_50 bitb_43_50 bitb_43_51 R_bl
Cb_43_50 bit_43_50 gnd C_bl
Cbb_43_50 bitb_43_50 gnd C_bl
Rb_43_51 bit_43_51 bit_43_52 R_bl
Rbb_43_51 bitb_43_51 bitb_43_52 R_bl
Cb_43_51 bit_43_51 gnd C_bl
Cbb_43_51 bitb_43_51 gnd C_bl
Rb_43_52 bit_43_52 bit_43_53 R_bl
Rbb_43_52 bitb_43_52 bitb_43_53 R_bl
Cb_43_52 bit_43_52 gnd C_bl
Cbb_43_52 bitb_43_52 gnd C_bl
Rb_43_53 bit_43_53 bit_43_54 R_bl
Rbb_43_53 bitb_43_53 bitb_43_54 R_bl
Cb_43_53 bit_43_53 gnd C_bl
Cbb_43_53 bitb_43_53 gnd C_bl
Rb_43_54 bit_43_54 bit_43_55 R_bl
Rbb_43_54 bitb_43_54 bitb_43_55 R_bl
Cb_43_54 bit_43_54 gnd C_bl
Cbb_43_54 bitb_43_54 gnd C_bl
Rb_43_55 bit_43_55 bit_43_56 R_bl
Rbb_43_55 bitb_43_55 bitb_43_56 R_bl
Cb_43_55 bit_43_55 gnd C_bl
Cbb_43_55 bitb_43_55 gnd C_bl
Rb_43_56 bit_43_56 bit_43_57 R_bl
Rbb_43_56 bitb_43_56 bitb_43_57 R_bl
Cb_43_56 bit_43_56 gnd C_bl
Cbb_43_56 bitb_43_56 gnd C_bl
Rb_43_57 bit_43_57 bit_43_58 R_bl
Rbb_43_57 bitb_43_57 bitb_43_58 R_bl
Cb_43_57 bit_43_57 gnd C_bl
Cbb_43_57 bitb_43_57 gnd C_bl
Rb_43_58 bit_43_58 bit_43_59 R_bl
Rbb_43_58 bitb_43_58 bitb_43_59 R_bl
Cb_43_58 bit_43_58 gnd C_bl
Cbb_43_58 bitb_43_58 gnd C_bl
Rb_43_59 bit_43_59 bit_43_60 R_bl
Rbb_43_59 bitb_43_59 bitb_43_60 R_bl
Cb_43_59 bit_43_59 gnd C_bl
Cbb_43_59 bitb_43_59 gnd C_bl
Rb_43_60 bit_43_60 bit_43_61 R_bl
Rbb_43_60 bitb_43_60 bitb_43_61 R_bl
Cb_43_60 bit_43_60 gnd C_bl
Cbb_43_60 bitb_43_60 gnd C_bl
Rb_43_61 bit_43_61 bit_43_62 R_bl
Rbb_43_61 bitb_43_61 bitb_43_62 R_bl
Cb_43_61 bit_43_61 gnd C_bl
Cbb_43_61 bitb_43_61 gnd C_bl
Rb_43_62 bit_43_62 bit_43_63 R_bl
Rbb_43_62 bitb_43_62 bitb_43_63 R_bl
Cb_43_62 bit_43_62 gnd C_bl
Cbb_43_62 bitb_43_62 gnd C_bl
Rb_43_63 bit_43_63 bit_43_64 R_bl
Rbb_43_63 bitb_43_63 bitb_43_64 R_bl
Cb_43_63 bit_43_63 gnd C_bl
Cbb_43_63 bitb_43_63 gnd C_bl
Rb_43_64 bit_43_64 bit_43_65 R_bl
Rbb_43_64 bitb_43_64 bitb_43_65 R_bl
Cb_43_64 bit_43_64 gnd C_bl
Cbb_43_64 bitb_43_64 gnd C_bl
Rb_43_65 bit_43_65 bit_43_66 R_bl
Rbb_43_65 bitb_43_65 bitb_43_66 R_bl
Cb_43_65 bit_43_65 gnd C_bl
Cbb_43_65 bitb_43_65 gnd C_bl
Rb_43_66 bit_43_66 bit_43_67 R_bl
Rbb_43_66 bitb_43_66 bitb_43_67 R_bl
Cb_43_66 bit_43_66 gnd C_bl
Cbb_43_66 bitb_43_66 gnd C_bl
Rb_43_67 bit_43_67 bit_43_68 R_bl
Rbb_43_67 bitb_43_67 bitb_43_68 R_bl
Cb_43_67 bit_43_67 gnd C_bl
Cbb_43_67 bitb_43_67 gnd C_bl
Rb_43_68 bit_43_68 bit_43_69 R_bl
Rbb_43_68 bitb_43_68 bitb_43_69 R_bl
Cb_43_68 bit_43_68 gnd C_bl
Cbb_43_68 bitb_43_68 gnd C_bl
Rb_43_69 bit_43_69 bit_43_70 R_bl
Rbb_43_69 bitb_43_69 bitb_43_70 R_bl
Cb_43_69 bit_43_69 gnd C_bl
Cbb_43_69 bitb_43_69 gnd C_bl
Rb_43_70 bit_43_70 bit_43_71 R_bl
Rbb_43_70 bitb_43_70 bitb_43_71 R_bl
Cb_43_70 bit_43_70 gnd C_bl
Cbb_43_70 bitb_43_70 gnd C_bl
Rb_43_71 bit_43_71 bit_43_72 R_bl
Rbb_43_71 bitb_43_71 bitb_43_72 R_bl
Cb_43_71 bit_43_71 gnd C_bl
Cbb_43_71 bitb_43_71 gnd C_bl
Rb_43_72 bit_43_72 bit_43_73 R_bl
Rbb_43_72 bitb_43_72 bitb_43_73 R_bl
Cb_43_72 bit_43_72 gnd C_bl
Cbb_43_72 bitb_43_72 gnd C_bl
Rb_43_73 bit_43_73 bit_43_74 R_bl
Rbb_43_73 bitb_43_73 bitb_43_74 R_bl
Cb_43_73 bit_43_73 gnd C_bl
Cbb_43_73 bitb_43_73 gnd C_bl
Rb_43_74 bit_43_74 bit_43_75 R_bl
Rbb_43_74 bitb_43_74 bitb_43_75 R_bl
Cb_43_74 bit_43_74 gnd C_bl
Cbb_43_74 bitb_43_74 gnd C_bl
Rb_43_75 bit_43_75 bit_43_76 R_bl
Rbb_43_75 bitb_43_75 bitb_43_76 R_bl
Cb_43_75 bit_43_75 gnd C_bl
Cbb_43_75 bitb_43_75 gnd C_bl
Rb_43_76 bit_43_76 bit_43_77 R_bl
Rbb_43_76 bitb_43_76 bitb_43_77 R_bl
Cb_43_76 bit_43_76 gnd C_bl
Cbb_43_76 bitb_43_76 gnd C_bl
Rb_43_77 bit_43_77 bit_43_78 R_bl
Rbb_43_77 bitb_43_77 bitb_43_78 R_bl
Cb_43_77 bit_43_77 gnd C_bl
Cbb_43_77 bitb_43_77 gnd C_bl
Rb_43_78 bit_43_78 bit_43_79 R_bl
Rbb_43_78 bitb_43_78 bitb_43_79 R_bl
Cb_43_78 bit_43_78 gnd C_bl
Cbb_43_78 bitb_43_78 gnd C_bl
Rb_43_79 bit_43_79 bit_43_80 R_bl
Rbb_43_79 bitb_43_79 bitb_43_80 R_bl
Cb_43_79 bit_43_79 gnd C_bl
Cbb_43_79 bitb_43_79 gnd C_bl
Rb_43_80 bit_43_80 bit_43_81 R_bl
Rbb_43_80 bitb_43_80 bitb_43_81 R_bl
Cb_43_80 bit_43_80 gnd C_bl
Cbb_43_80 bitb_43_80 gnd C_bl
Rb_43_81 bit_43_81 bit_43_82 R_bl
Rbb_43_81 bitb_43_81 bitb_43_82 R_bl
Cb_43_81 bit_43_81 gnd C_bl
Cbb_43_81 bitb_43_81 gnd C_bl
Rb_43_82 bit_43_82 bit_43_83 R_bl
Rbb_43_82 bitb_43_82 bitb_43_83 R_bl
Cb_43_82 bit_43_82 gnd C_bl
Cbb_43_82 bitb_43_82 gnd C_bl
Rb_43_83 bit_43_83 bit_43_84 R_bl
Rbb_43_83 bitb_43_83 bitb_43_84 R_bl
Cb_43_83 bit_43_83 gnd C_bl
Cbb_43_83 bitb_43_83 gnd C_bl
Rb_43_84 bit_43_84 bit_43_85 R_bl
Rbb_43_84 bitb_43_84 bitb_43_85 R_bl
Cb_43_84 bit_43_84 gnd C_bl
Cbb_43_84 bitb_43_84 gnd C_bl
Rb_43_85 bit_43_85 bit_43_86 R_bl
Rbb_43_85 bitb_43_85 bitb_43_86 R_bl
Cb_43_85 bit_43_85 gnd C_bl
Cbb_43_85 bitb_43_85 gnd C_bl
Rb_43_86 bit_43_86 bit_43_87 R_bl
Rbb_43_86 bitb_43_86 bitb_43_87 R_bl
Cb_43_86 bit_43_86 gnd C_bl
Cbb_43_86 bitb_43_86 gnd C_bl
Rb_43_87 bit_43_87 bit_43_88 R_bl
Rbb_43_87 bitb_43_87 bitb_43_88 R_bl
Cb_43_87 bit_43_87 gnd C_bl
Cbb_43_87 bitb_43_87 gnd C_bl
Rb_43_88 bit_43_88 bit_43_89 R_bl
Rbb_43_88 bitb_43_88 bitb_43_89 R_bl
Cb_43_88 bit_43_88 gnd C_bl
Cbb_43_88 bitb_43_88 gnd C_bl
Rb_43_89 bit_43_89 bit_43_90 R_bl
Rbb_43_89 bitb_43_89 bitb_43_90 R_bl
Cb_43_89 bit_43_89 gnd C_bl
Cbb_43_89 bitb_43_89 gnd C_bl
Rb_43_90 bit_43_90 bit_43_91 R_bl
Rbb_43_90 bitb_43_90 bitb_43_91 R_bl
Cb_43_90 bit_43_90 gnd C_bl
Cbb_43_90 bitb_43_90 gnd C_bl
Rb_43_91 bit_43_91 bit_43_92 R_bl
Rbb_43_91 bitb_43_91 bitb_43_92 R_bl
Cb_43_91 bit_43_91 gnd C_bl
Cbb_43_91 bitb_43_91 gnd C_bl
Rb_43_92 bit_43_92 bit_43_93 R_bl
Rbb_43_92 bitb_43_92 bitb_43_93 R_bl
Cb_43_92 bit_43_92 gnd C_bl
Cbb_43_92 bitb_43_92 gnd C_bl
Rb_43_93 bit_43_93 bit_43_94 R_bl
Rbb_43_93 bitb_43_93 bitb_43_94 R_bl
Cb_43_93 bit_43_93 gnd C_bl
Cbb_43_93 bitb_43_93 gnd C_bl
Rb_43_94 bit_43_94 bit_43_95 R_bl
Rbb_43_94 bitb_43_94 bitb_43_95 R_bl
Cb_43_94 bit_43_94 gnd C_bl
Cbb_43_94 bitb_43_94 gnd C_bl
Rb_43_95 bit_43_95 bit_43_96 R_bl
Rbb_43_95 bitb_43_95 bitb_43_96 R_bl
Cb_43_95 bit_43_95 gnd C_bl
Cbb_43_95 bitb_43_95 gnd C_bl
Rb_43_96 bit_43_96 bit_43_97 R_bl
Rbb_43_96 bitb_43_96 bitb_43_97 R_bl
Cb_43_96 bit_43_96 gnd C_bl
Cbb_43_96 bitb_43_96 gnd C_bl
Rb_43_97 bit_43_97 bit_43_98 R_bl
Rbb_43_97 bitb_43_97 bitb_43_98 R_bl
Cb_43_97 bit_43_97 gnd C_bl
Cbb_43_97 bitb_43_97 gnd C_bl
Rb_43_98 bit_43_98 bit_43_99 R_bl
Rbb_43_98 bitb_43_98 bitb_43_99 R_bl
Cb_43_98 bit_43_98 gnd C_bl
Cbb_43_98 bitb_43_98 gnd C_bl
Rb_43_99 bit_43_99 bit_43_100 R_bl
Rbb_43_99 bitb_43_99 bitb_43_100 R_bl
Cb_43_99 bit_43_99 gnd C_bl
Cbb_43_99 bitb_43_99 gnd C_bl
Rb_44_0 bit_44_0 bit_44_1 R_bl
Rbb_44_0 bitb_44_0 bitb_44_1 R_bl
Cb_44_0 bit_44_0 gnd C_bl
Cbb_44_0 bitb_44_0 gnd C_bl
Rb_44_1 bit_44_1 bit_44_2 R_bl
Rbb_44_1 bitb_44_1 bitb_44_2 R_bl
Cb_44_1 bit_44_1 gnd C_bl
Cbb_44_1 bitb_44_1 gnd C_bl
Rb_44_2 bit_44_2 bit_44_3 R_bl
Rbb_44_2 bitb_44_2 bitb_44_3 R_bl
Cb_44_2 bit_44_2 gnd C_bl
Cbb_44_2 bitb_44_2 gnd C_bl
Rb_44_3 bit_44_3 bit_44_4 R_bl
Rbb_44_3 bitb_44_3 bitb_44_4 R_bl
Cb_44_3 bit_44_3 gnd C_bl
Cbb_44_3 bitb_44_3 gnd C_bl
Rb_44_4 bit_44_4 bit_44_5 R_bl
Rbb_44_4 bitb_44_4 bitb_44_5 R_bl
Cb_44_4 bit_44_4 gnd C_bl
Cbb_44_4 bitb_44_4 gnd C_bl
Rb_44_5 bit_44_5 bit_44_6 R_bl
Rbb_44_5 bitb_44_5 bitb_44_6 R_bl
Cb_44_5 bit_44_5 gnd C_bl
Cbb_44_5 bitb_44_5 gnd C_bl
Rb_44_6 bit_44_6 bit_44_7 R_bl
Rbb_44_6 bitb_44_6 bitb_44_7 R_bl
Cb_44_6 bit_44_6 gnd C_bl
Cbb_44_6 bitb_44_6 gnd C_bl
Rb_44_7 bit_44_7 bit_44_8 R_bl
Rbb_44_7 bitb_44_7 bitb_44_8 R_bl
Cb_44_7 bit_44_7 gnd C_bl
Cbb_44_7 bitb_44_7 gnd C_bl
Rb_44_8 bit_44_8 bit_44_9 R_bl
Rbb_44_8 bitb_44_8 bitb_44_9 R_bl
Cb_44_8 bit_44_8 gnd C_bl
Cbb_44_8 bitb_44_8 gnd C_bl
Rb_44_9 bit_44_9 bit_44_10 R_bl
Rbb_44_9 bitb_44_9 bitb_44_10 R_bl
Cb_44_9 bit_44_9 gnd C_bl
Cbb_44_9 bitb_44_9 gnd C_bl
Rb_44_10 bit_44_10 bit_44_11 R_bl
Rbb_44_10 bitb_44_10 bitb_44_11 R_bl
Cb_44_10 bit_44_10 gnd C_bl
Cbb_44_10 bitb_44_10 gnd C_bl
Rb_44_11 bit_44_11 bit_44_12 R_bl
Rbb_44_11 bitb_44_11 bitb_44_12 R_bl
Cb_44_11 bit_44_11 gnd C_bl
Cbb_44_11 bitb_44_11 gnd C_bl
Rb_44_12 bit_44_12 bit_44_13 R_bl
Rbb_44_12 bitb_44_12 bitb_44_13 R_bl
Cb_44_12 bit_44_12 gnd C_bl
Cbb_44_12 bitb_44_12 gnd C_bl
Rb_44_13 bit_44_13 bit_44_14 R_bl
Rbb_44_13 bitb_44_13 bitb_44_14 R_bl
Cb_44_13 bit_44_13 gnd C_bl
Cbb_44_13 bitb_44_13 gnd C_bl
Rb_44_14 bit_44_14 bit_44_15 R_bl
Rbb_44_14 bitb_44_14 bitb_44_15 R_bl
Cb_44_14 bit_44_14 gnd C_bl
Cbb_44_14 bitb_44_14 gnd C_bl
Rb_44_15 bit_44_15 bit_44_16 R_bl
Rbb_44_15 bitb_44_15 bitb_44_16 R_bl
Cb_44_15 bit_44_15 gnd C_bl
Cbb_44_15 bitb_44_15 gnd C_bl
Rb_44_16 bit_44_16 bit_44_17 R_bl
Rbb_44_16 bitb_44_16 bitb_44_17 R_bl
Cb_44_16 bit_44_16 gnd C_bl
Cbb_44_16 bitb_44_16 gnd C_bl
Rb_44_17 bit_44_17 bit_44_18 R_bl
Rbb_44_17 bitb_44_17 bitb_44_18 R_bl
Cb_44_17 bit_44_17 gnd C_bl
Cbb_44_17 bitb_44_17 gnd C_bl
Rb_44_18 bit_44_18 bit_44_19 R_bl
Rbb_44_18 bitb_44_18 bitb_44_19 R_bl
Cb_44_18 bit_44_18 gnd C_bl
Cbb_44_18 bitb_44_18 gnd C_bl
Rb_44_19 bit_44_19 bit_44_20 R_bl
Rbb_44_19 bitb_44_19 bitb_44_20 R_bl
Cb_44_19 bit_44_19 gnd C_bl
Cbb_44_19 bitb_44_19 gnd C_bl
Rb_44_20 bit_44_20 bit_44_21 R_bl
Rbb_44_20 bitb_44_20 bitb_44_21 R_bl
Cb_44_20 bit_44_20 gnd C_bl
Cbb_44_20 bitb_44_20 gnd C_bl
Rb_44_21 bit_44_21 bit_44_22 R_bl
Rbb_44_21 bitb_44_21 bitb_44_22 R_bl
Cb_44_21 bit_44_21 gnd C_bl
Cbb_44_21 bitb_44_21 gnd C_bl
Rb_44_22 bit_44_22 bit_44_23 R_bl
Rbb_44_22 bitb_44_22 bitb_44_23 R_bl
Cb_44_22 bit_44_22 gnd C_bl
Cbb_44_22 bitb_44_22 gnd C_bl
Rb_44_23 bit_44_23 bit_44_24 R_bl
Rbb_44_23 bitb_44_23 bitb_44_24 R_bl
Cb_44_23 bit_44_23 gnd C_bl
Cbb_44_23 bitb_44_23 gnd C_bl
Rb_44_24 bit_44_24 bit_44_25 R_bl
Rbb_44_24 bitb_44_24 bitb_44_25 R_bl
Cb_44_24 bit_44_24 gnd C_bl
Cbb_44_24 bitb_44_24 gnd C_bl
Rb_44_25 bit_44_25 bit_44_26 R_bl
Rbb_44_25 bitb_44_25 bitb_44_26 R_bl
Cb_44_25 bit_44_25 gnd C_bl
Cbb_44_25 bitb_44_25 gnd C_bl
Rb_44_26 bit_44_26 bit_44_27 R_bl
Rbb_44_26 bitb_44_26 bitb_44_27 R_bl
Cb_44_26 bit_44_26 gnd C_bl
Cbb_44_26 bitb_44_26 gnd C_bl
Rb_44_27 bit_44_27 bit_44_28 R_bl
Rbb_44_27 bitb_44_27 bitb_44_28 R_bl
Cb_44_27 bit_44_27 gnd C_bl
Cbb_44_27 bitb_44_27 gnd C_bl
Rb_44_28 bit_44_28 bit_44_29 R_bl
Rbb_44_28 bitb_44_28 bitb_44_29 R_bl
Cb_44_28 bit_44_28 gnd C_bl
Cbb_44_28 bitb_44_28 gnd C_bl
Rb_44_29 bit_44_29 bit_44_30 R_bl
Rbb_44_29 bitb_44_29 bitb_44_30 R_bl
Cb_44_29 bit_44_29 gnd C_bl
Cbb_44_29 bitb_44_29 gnd C_bl
Rb_44_30 bit_44_30 bit_44_31 R_bl
Rbb_44_30 bitb_44_30 bitb_44_31 R_bl
Cb_44_30 bit_44_30 gnd C_bl
Cbb_44_30 bitb_44_30 gnd C_bl
Rb_44_31 bit_44_31 bit_44_32 R_bl
Rbb_44_31 bitb_44_31 bitb_44_32 R_bl
Cb_44_31 bit_44_31 gnd C_bl
Cbb_44_31 bitb_44_31 gnd C_bl
Rb_44_32 bit_44_32 bit_44_33 R_bl
Rbb_44_32 bitb_44_32 bitb_44_33 R_bl
Cb_44_32 bit_44_32 gnd C_bl
Cbb_44_32 bitb_44_32 gnd C_bl
Rb_44_33 bit_44_33 bit_44_34 R_bl
Rbb_44_33 bitb_44_33 bitb_44_34 R_bl
Cb_44_33 bit_44_33 gnd C_bl
Cbb_44_33 bitb_44_33 gnd C_bl
Rb_44_34 bit_44_34 bit_44_35 R_bl
Rbb_44_34 bitb_44_34 bitb_44_35 R_bl
Cb_44_34 bit_44_34 gnd C_bl
Cbb_44_34 bitb_44_34 gnd C_bl
Rb_44_35 bit_44_35 bit_44_36 R_bl
Rbb_44_35 bitb_44_35 bitb_44_36 R_bl
Cb_44_35 bit_44_35 gnd C_bl
Cbb_44_35 bitb_44_35 gnd C_bl
Rb_44_36 bit_44_36 bit_44_37 R_bl
Rbb_44_36 bitb_44_36 bitb_44_37 R_bl
Cb_44_36 bit_44_36 gnd C_bl
Cbb_44_36 bitb_44_36 gnd C_bl
Rb_44_37 bit_44_37 bit_44_38 R_bl
Rbb_44_37 bitb_44_37 bitb_44_38 R_bl
Cb_44_37 bit_44_37 gnd C_bl
Cbb_44_37 bitb_44_37 gnd C_bl
Rb_44_38 bit_44_38 bit_44_39 R_bl
Rbb_44_38 bitb_44_38 bitb_44_39 R_bl
Cb_44_38 bit_44_38 gnd C_bl
Cbb_44_38 bitb_44_38 gnd C_bl
Rb_44_39 bit_44_39 bit_44_40 R_bl
Rbb_44_39 bitb_44_39 bitb_44_40 R_bl
Cb_44_39 bit_44_39 gnd C_bl
Cbb_44_39 bitb_44_39 gnd C_bl
Rb_44_40 bit_44_40 bit_44_41 R_bl
Rbb_44_40 bitb_44_40 bitb_44_41 R_bl
Cb_44_40 bit_44_40 gnd C_bl
Cbb_44_40 bitb_44_40 gnd C_bl
Rb_44_41 bit_44_41 bit_44_42 R_bl
Rbb_44_41 bitb_44_41 bitb_44_42 R_bl
Cb_44_41 bit_44_41 gnd C_bl
Cbb_44_41 bitb_44_41 gnd C_bl
Rb_44_42 bit_44_42 bit_44_43 R_bl
Rbb_44_42 bitb_44_42 bitb_44_43 R_bl
Cb_44_42 bit_44_42 gnd C_bl
Cbb_44_42 bitb_44_42 gnd C_bl
Rb_44_43 bit_44_43 bit_44_44 R_bl
Rbb_44_43 bitb_44_43 bitb_44_44 R_bl
Cb_44_43 bit_44_43 gnd C_bl
Cbb_44_43 bitb_44_43 gnd C_bl
Rb_44_44 bit_44_44 bit_44_45 R_bl
Rbb_44_44 bitb_44_44 bitb_44_45 R_bl
Cb_44_44 bit_44_44 gnd C_bl
Cbb_44_44 bitb_44_44 gnd C_bl
Rb_44_45 bit_44_45 bit_44_46 R_bl
Rbb_44_45 bitb_44_45 bitb_44_46 R_bl
Cb_44_45 bit_44_45 gnd C_bl
Cbb_44_45 bitb_44_45 gnd C_bl
Rb_44_46 bit_44_46 bit_44_47 R_bl
Rbb_44_46 bitb_44_46 bitb_44_47 R_bl
Cb_44_46 bit_44_46 gnd C_bl
Cbb_44_46 bitb_44_46 gnd C_bl
Rb_44_47 bit_44_47 bit_44_48 R_bl
Rbb_44_47 bitb_44_47 bitb_44_48 R_bl
Cb_44_47 bit_44_47 gnd C_bl
Cbb_44_47 bitb_44_47 gnd C_bl
Rb_44_48 bit_44_48 bit_44_49 R_bl
Rbb_44_48 bitb_44_48 bitb_44_49 R_bl
Cb_44_48 bit_44_48 gnd C_bl
Cbb_44_48 bitb_44_48 gnd C_bl
Rb_44_49 bit_44_49 bit_44_50 R_bl
Rbb_44_49 bitb_44_49 bitb_44_50 R_bl
Cb_44_49 bit_44_49 gnd C_bl
Cbb_44_49 bitb_44_49 gnd C_bl
Rb_44_50 bit_44_50 bit_44_51 R_bl
Rbb_44_50 bitb_44_50 bitb_44_51 R_bl
Cb_44_50 bit_44_50 gnd C_bl
Cbb_44_50 bitb_44_50 gnd C_bl
Rb_44_51 bit_44_51 bit_44_52 R_bl
Rbb_44_51 bitb_44_51 bitb_44_52 R_bl
Cb_44_51 bit_44_51 gnd C_bl
Cbb_44_51 bitb_44_51 gnd C_bl
Rb_44_52 bit_44_52 bit_44_53 R_bl
Rbb_44_52 bitb_44_52 bitb_44_53 R_bl
Cb_44_52 bit_44_52 gnd C_bl
Cbb_44_52 bitb_44_52 gnd C_bl
Rb_44_53 bit_44_53 bit_44_54 R_bl
Rbb_44_53 bitb_44_53 bitb_44_54 R_bl
Cb_44_53 bit_44_53 gnd C_bl
Cbb_44_53 bitb_44_53 gnd C_bl
Rb_44_54 bit_44_54 bit_44_55 R_bl
Rbb_44_54 bitb_44_54 bitb_44_55 R_bl
Cb_44_54 bit_44_54 gnd C_bl
Cbb_44_54 bitb_44_54 gnd C_bl
Rb_44_55 bit_44_55 bit_44_56 R_bl
Rbb_44_55 bitb_44_55 bitb_44_56 R_bl
Cb_44_55 bit_44_55 gnd C_bl
Cbb_44_55 bitb_44_55 gnd C_bl
Rb_44_56 bit_44_56 bit_44_57 R_bl
Rbb_44_56 bitb_44_56 bitb_44_57 R_bl
Cb_44_56 bit_44_56 gnd C_bl
Cbb_44_56 bitb_44_56 gnd C_bl
Rb_44_57 bit_44_57 bit_44_58 R_bl
Rbb_44_57 bitb_44_57 bitb_44_58 R_bl
Cb_44_57 bit_44_57 gnd C_bl
Cbb_44_57 bitb_44_57 gnd C_bl
Rb_44_58 bit_44_58 bit_44_59 R_bl
Rbb_44_58 bitb_44_58 bitb_44_59 R_bl
Cb_44_58 bit_44_58 gnd C_bl
Cbb_44_58 bitb_44_58 gnd C_bl
Rb_44_59 bit_44_59 bit_44_60 R_bl
Rbb_44_59 bitb_44_59 bitb_44_60 R_bl
Cb_44_59 bit_44_59 gnd C_bl
Cbb_44_59 bitb_44_59 gnd C_bl
Rb_44_60 bit_44_60 bit_44_61 R_bl
Rbb_44_60 bitb_44_60 bitb_44_61 R_bl
Cb_44_60 bit_44_60 gnd C_bl
Cbb_44_60 bitb_44_60 gnd C_bl
Rb_44_61 bit_44_61 bit_44_62 R_bl
Rbb_44_61 bitb_44_61 bitb_44_62 R_bl
Cb_44_61 bit_44_61 gnd C_bl
Cbb_44_61 bitb_44_61 gnd C_bl
Rb_44_62 bit_44_62 bit_44_63 R_bl
Rbb_44_62 bitb_44_62 bitb_44_63 R_bl
Cb_44_62 bit_44_62 gnd C_bl
Cbb_44_62 bitb_44_62 gnd C_bl
Rb_44_63 bit_44_63 bit_44_64 R_bl
Rbb_44_63 bitb_44_63 bitb_44_64 R_bl
Cb_44_63 bit_44_63 gnd C_bl
Cbb_44_63 bitb_44_63 gnd C_bl
Rb_44_64 bit_44_64 bit_44_65 R_bl
Rbb_44_64 bitb_44_64 bitb_44_65 R_bl
Cb_44_64 bit_44_64 gnd C_bl
Cbb_44_64 bitb_44_64 gnd C_bl
Rb_44_65 bit_44_65 bit_44_66 R_bl
Rbb_44_65 bitb_44_65 bitb_44_66 R_bl
Cb_44_65 bit_44_65 gnd C_bl
Cbb_44_65 bitb_44_65 gnd C_bl
Rb_44_66 bit_44_66 bit_44_67 R_bl
Rbb_44_66 bitb_44_66 bitb_44_67 R_bl
Cb_44_66 bit_44_66 gnd C_bl
Cbb_44_66 bitb_44_66 gnd C_bl
Rb_44_67 bit_44_67 bit_44_68 R_bl
Rbb_44_67 bitb_44_67 bitb_44_68 R_bl
Cb_44_67 bit_44_67 gnd C_bl
Cbb_44_67 bitb_44_67 gnd C_bl
Rb_44_68 bit_44_68 bit_44_69 R_bl
Rbb_44_68 bitb_44_68 bitb_44_69 R_bl
Cb_44_68 bit_44_68 gnd C_bl
Cbb_44_68 bitb_44_68 gnd C_bl
Rb_44_69 bit_44_69 bit_44_70 R_bl
Rbb_44_69 bitb_44_69 bitb_44_70 R_bl
Cb_44_69 bit_44_69 gnd C_bl
Cbb_44_69 bitb_44_69 gnd C_bl
Rb_44_70 bit_44_70 bit_44_71 R_bl
Rbb_44_70 bitb_44_70 bitb_44_71 R_bl
Cb_44_70 bit_44_70 gnd C_bl
Cbb_44_70 bitb_44_70 gnd C_bl
Rb_44_71 bit_44_71 bit_44_72 R_bl
Rbb_44_71 bitb_44_71 bitb_44_72 R_bl
Cb_44_71 bit_44_71 gnd C_bl
Cbb_44_71 bitb_44_71 gnd C_bl
Rb_44_72 bit_44_72 bit_44_73 R_bl
Rbb_44_72 bitb_44_72 bitb_44_73 R_bl
Cb_44_72 bit_44_72 gnd C_bl
Cbb_44_72 bitb_44_72 gnd C_bl
Rb_44_73 bit_44_73 bit_44_74 R_bl
Rbb_44_73 bitb_44_73 bitb_44_74 R_bl
Cb_44_73 bit_44_73 gnd C_bl
Cbb_44_73 bitb_44_73 gnd C_bl
Rb_44_74 bit_44_74 bit_44_75 R_bl
Rbb_44_74 bitb_44_74 bitb_44_75 R_bl
Cb_44_74 bit_44_74 gnd C_bl
Cbb_44_74 bitb_44_74 gnd C_bl
Rb_44_75 bit_44_75 bit_44_76 R_bl
Rbb_44_75 bitb_44_75 bitb_44_76 R_bl
Cb_44_75 bit_44_75 gnd C_bl
Cbb_44_75 bitb_44_75 gnd C_bl
Rb_44_76 bit_44_76 bit_44_77 R_bl
Rbb_44_76 bitb_44_76 bitb_44_77 R_bl
Cb_44_76 bit_44_76 gnd C_bl
Cbb_44_76 bitb_44_76 gnd C_bl
Rb_44_77 bit_44_77 bit_44_78 R_bl
Rbb_44_77 bitb_44_77 bitb_44_78 R_bl
Cb_44_77 bit_44_77 gnd C_bl
Cbb_44_77 bitb_44_77 gnd C_bl
Rb_44_78 bit_44_78 bit_44_79 R_bl
Rbb_44_78 bitb_44_78 bitb_44_79 R_bl
Cb_44_78 bit_44_78 gnd C_bl
Cbb_44_78 bitb_44_78 gnd C_bl
Rb_44_79 bit_44_79 bit_44_80 R_bl
Rbb_44_79 bitb_44_79 bitb_44_80 R_bl
Cb_44_79 bit_44_79 gnd C_bl
Cbb_44_79 bitb_44_79 gnd C_bl
Rb_44_80 bit_44_80 bit_44_81 R_bl
Rbb_44_80 bitb_44_80 bitb_44_81 R_bl
Cb_44_80 bit_44_80 gnd C_bl
Cbb_44_80 bitb_44_80 gnd C_bl
Rb_44_81 bit_44_81 bit_44_82 R_bl
Rbb_44_81 bitb_44_81 bitb_44_82 R_bl
Cb_44_81 bit_44_81 gnd C_bl
Cbb_44_81 bitb_44_81 gnd C_bl
Rb_44_82 bit_44_82 bit_44_83 R_bl
Rbb_44_82 bitb_44_82 bitb_44_83 R_bl
Cb_44_82 bit_44_82 gnd C_bl
Cbb_44_82 bitb_44_82 gnd C_bl
Rb_44_83 bit_44_83 bit_44_84 R_bl
Rbb_44_83 bitb_44_83 bitb_44_84 R_bl
Cb_44_83 bit_44_83 gnd C_bl
Cbb_44_83 bitb_44_83 gnd C_bl
Rb_44_84 bit_44_84 bit_44_85 R_bl
Rbb_44_84 bitb_44_84 bitb_44_85 R_bl
Cb_44_84 bit_44_84 gnd C_bl
Cbb_44_84 bitb_44_84 gnd C_bl
Rb_44_85 bit_44_85 bit_44_86 R_bl
Rbb_44_85 bitb_44_85 bitb_44_86 R_bl
Cb_44_85 bit_44_85 gnd C_bl
Cbb_44_85 bitb_44_85 gnd C_bl
Rb_44_86 bit_44_86 bit_44_87 R_bl
Rbb_44_86 bitb_44_86 bitb_44_87 R_bl
Cb_44_86 bit_44_86 gnd C_bl
Cbb_44_86 bitb_44_86 gnd C_bl
Rb_44_87 bit_44_87 bit_44_88 R_bl
Rbb_44_87 bitb_44_87 bitb_44_88 R_bl
Cb_44_87 bit_44_87 gnd C_bl
Cbb_44_87 bitb_44_87 gnd C_bl
Rb_44_88 bit_44_88 bit_44_89 R_bl
Rbb_44_88 bitb_44_88 bitb_44_89 R_bl
Cb_44_88 bit_44_88 gnd C_bl
Cbb_44_88 bitb_44_88 gnd C_bl
Rb_44_89 bit_44_89 bit_44_90 R_bl
Rbb_44_89 bitb_44_89 bitb_44_90 R_bl
Cb_44_89 bit_44_89 gnd C_bl
Cbb_44_89 bitb_44_89 gnd C_bl
Rb_44_90 bit_44_90 bit_44_91 R_bl
Rbb_44_90 bitb_44_90 bitb_44_91 R_bl
Cb_44_90 bit_44_90 gnd C_bl
Cbb_44_90 bitb_44_90 gnd C_bl
Rb_44_91 bit_44_91 bit_44_92 R_bl
Rbb_44_91 bitb_44_91 bitb_44_92 R_bl
Cb_44_91 bit_44_91 gnd C_bl
Cbb_44_91 bitb_44_91 gnd C_bl
Rb_44_92 bit_44_92 bit_44_93 R_bl
Rbb_44_92 bitb_44_92 bitb_44_93 R_bl
Cb_44_92 bit_44_92 gnd C_bl
Cbb_44_92 bitb_44_92 gnd C_bl
Rb_44_93 bit_44_93 bit_44_94 R_bl
Rbb_44_93 bitb_44_93 bitb_44_94 R_bl
Cb_44_93 bit_44_93 gnd C_bl
Cbb_44_93 bitb_44_93 gnd C_bl
Rb_44_94 bit_44_94 bit_44_95 R_bl
Rbb_44_94 bitb_44_94 bitb_44_95 R_bl
Cb_44_94 bit_44_94 gnd C_bl
Cbb_44_94 bitb_44_94 gnd C_bl
Rb_44_95 bit_44_95 bit_44_96 R_bl
Rbb_44_95 bitb_44_95 bitb_44_96 R_bl
Cb_44_95 bit_44_95 gnd C_bl
Cbb_44_95 bitb_44_95 gnd C_bl
Rb_44_96 bit_44_96 bit_44_97 R_bl
Rbb_44_96 bitb_44_96 bitb_44_97 R_bl
Cb_44_96 bit_44_96 gnd C_bl
Cbb_44_96 bitb_44_96 gnd C_bl
Rb_44_97 bit_44_97 bit_44_98 R_bl
Rbb_44_97 bitb_44_97 bitb_44_98 R_bl
Cb_44_97 bit_44_97 gnd C_bl
Cbb_44_97 bitb_44_97 gnd C_bl
Rb_44_98 bit_44_98 bit_44_99 R_bl
Rbb_44_98 bitb_44_98 bitb_44_99 R_bl
Cb_44_98 bit_44_98 gnd C_bl
Cbb_44_98 bitb_44_98 gnd C_bl
Rb_44_99 bit_44_99 bit_44_100 R_bl
Rbb_44_99 bitb_44_99 bitb_44_100 R_bl
Cb_44_99 bit_44_99 gnd C_bl
Cbb_44_99 bitb_44_99 gnd C_bl
Rb_45_0 bit_45_0 bit_45_1 R_bl
Rbb_45_0 bitb_45_0 bitb_45_1 R_bl
Cb_45_0 bit_45_0 gnd C_bl
Cbb_45_0 bitb_45_0 gnd C_bl
Rb_45_1 bit_45_1 bit_45_2 R_bl
Rbb_45_1 bitb_45_1 bitb_45_2 R_bl
Cb_45_1 bit_45_1 gnd C_bl
Cbb_45_1 bitb_45_1 gnd C_bl
Rb_45_2 bit_45_2 bit_45_3 R_bl
Rbb_45_2 bitb_45_2 bitb_45_3 R_bl
Cb_45_2 bit_45_2 gnd C_bl
Cbb_45_2 bitb_45_2 gnd C_bl
Rb_45_3 bit_45_3 bit_45_4 R_bl
Rbb_45_3 bitb_45_3 bitb_45_4 R_bl
Cb_45_3 bit_45_3 gnd C_bl
Cbb_45_3 bitb_45_3 gnd C_bl
Rb_45_4 bit_45_4 bit_45_5 R_bl
Rbb_45_4 bitb_45_4 bitb_45_5 R_bl
Cb_45_4 bit_45_4 gnd C_bl
Cbb_45_4 bitb_45_4 gnd C_bl
Rb_45_5 bit_45_5 bit_45_6 R_bl
Rbb_45_5 bitb_45_5 bitb_45_6 R_bl
Cb_45_5 bit_45_5 gnd C_bl
Cbb_45_5 bitb_45_5 gnd C_bl
Rb_45_6 bit_45_6 bit_45_7 R_bl
Rbb_45_6 bitb_45_6 bitb_45_7 R_bl
Cb_45_6 bit_45_6 gnd C_bl
Cbb_45_6 bitb_45_6 gnd C_bl
Rb_45_7 bit_45_7 bit_45_8 R_bl
Rbb_45_7 bitb_45_7 bitb_45_8 R_bl
Cb_45_7 bit_45_7 gnd C_bl
Cbb_45_7 bitb_45_7 gnd C_bl
Rb_45_8 bit_45_8 bit_45_9 R_bl
Rbb_45_8 bitb_45_8 bitb_45_9 R_bl
Cb_45_8 bit_45_8 gnd C_bl
Cbb_45_8 bitb_45_8 gnd C_bl
Rb_45_9 bit_45_9 bit_45_10 R_bl
Rbb_45_9 bitb_45_9 bitb_45_10 R_bl
Cb_45_9 bit_45_9 gnd C_bl
Cbb_45_9 bitb_45_9 gnd C_bl
Rb_45_10 bit_45_10 bit_45_11 R_bl
Rbb_45_10 bitb_45_10 bitb_45_11 R_bl
Cb_45_10 bit_45_10 gnd C_bl
Cbb_45_10 bitb_45_10 gnd C_bl
Rb_45_11 bit_45_11 bit_45_12 R_bl
Rbb_45_11 bitb_45_11 bitb_45_12 R_bl
Cb_45_11 bit_45_11 gnd C_bl
Cbb_45_11 bitb_45_11 gnd C_bl
Rb_45_12 bit_45_12 bit_45_13 R_bl
Rbb_45_12 bitb_45_12 bitb_45_13 R_bl
Cb_45_12 bit_45_12 gnd C_bl
Cbb_45_12 bitb_45_12 gnd C_bl
Rb_45_13 bit_45_13 bit_45_14 R_bl
Rbb_45_13 bitb_45_13 bitb_45_14 R_bl
Cb_45_13 bit_45_13 gnd C_bl
Cbb_45_13 bitb_45_13 gnd C_bl
Rb_45_14 bit_45_14 bit_45_15 R_bl
Rbb_45_14 bitb_45_14 bitb_45_15 R_bl
Cb_45_14 bit_45_14 gnd C_bl
Cbb_45_14 bitb_45_14 gnd C_bl
Rb_45_15 bit_45_15 bit_45_16 R_bl
Rbb_45_15 bitb_45_15 bitb_45_16 R_bl
Cb_45_15 bit_45_15 gnd C_bl
Cbb_45_15 bitb_45_15 gnd C_bl
Rb_45_16 bit_45_16 bit_45_17 R_bl
Rbb_45_16 bitb_45_16 bitb_45_17 R_bl
Cb_45_16 bit_45_16 gnd C_bl
Cbb_45_16 bitb_45_16 gnd C_bl
Rb_45_17 bit_45_17 bit_45_18 R_bl
Rbb_45_17 bitb_45_17 bitb_45_18 R_bl
Cb_45_17 bit_45_17 gnd C_bl
Cbb_45_17 bitb_45_17 gnd C_bl
Rb_45_18 bit_45_18 bit_45_19 R_bl
Rbb_45_18 bitb_45_18 bitb_45_19 R_bl
Cb_45_18 bit_45_18 gnd C_bl
Cbb_45_18 bitb_45_18 gnd C_bl
Rb_45_19 bit_45_19 bit_45_20 R_bl
Rbb_45_19 bitb_45_19 bitb_45_20 R_bl
Cb_45_19 bit_45_19 gnd C_bl
Cbb_45_19 bitb_45_19 gnd C_bl
Rb_45_20 bit_45_20 bit_45_21 R_bl
Rbb_45_20 bitb_45_20 bitb_45_21 R_bl
Cb_45_20 bit_45_20 gnd C_bl
Cbb_45_20 bitb_45_20 gnd C_bl
Rb_45_21 bit_45_21 bit_45_22 R_bl
Rbb_45_21 bitb_45_21 bitb_45_22 R_bl
Cb_45_21 bit_45_21 gnd C_bl
Cbb_45_21 bitb_45_21 gnd C_bl
Rb_45_22 bit_45_22 bit_45_23 R_bl
Rbb_45_22 bitb_45_22 bitb_45_23 R_bl
Cb_45_22 bit_45_22 gnd C_bl
Cbb_45_22 bitb_45_22 gnd C_bl
Rb_45_23 bit_45_23 bit_45_24 R_bl
Rbb_45_23 bitb_45_23 bitb_45_24 R_bl
Cb_45_23 bit_45_23 gnd C_bl
Cbb_45_23 bitb_45_23 gnd C_bl
Rb_45_24 bit_45_24 bit_45_25 R_bl
Rbb_45_24 bitb_45_24 bitb_45_25 R_bl
Cb_45_24 bit_45_24 gnd C_bl
Cbb_45_24 bitb_45_24 gnd C_bl
Rb_45_25 bit_45_25 bit_45_26 R_bl
Rbb_45_25 bitb_45_25 bitb_45_26 R_bl
Cb_45_25 bit_45_25 gnd C_bl
Cbb_45_25 bitb_45_25 gnd C_bl
Rb_45_26 bit_45_26 bit_45_27 R_bl
Rbb_45_26 bitb_45_26 bitb_45_27 R_bl
Cb_45_26 bit_45_26 gnd C_bl
Cbb_45_26 bitb_45_26 gnd C_bl
Rb_45_27 bit_45_27 bit_45_28 R_bl
Rbb_45_27 bitb_45_27 bitb_45_28 R_bl
Cb_45_27 bit_45_27 gnd C_bl
Cbb_45_27 bitb_45_27 gnd C_bl
Rb_45_28 bit_45_28 bit_45_29 R_bl
Rbb_45_28 bitb_45_28 bitb_45_29 R_bl
Cb_45_28 bit_45_28 gnd C_bl
Cbb_45_28 bitb_45_28 gnd C_bl
Rb_45_29 bit_45_29 bit_45_30 R_bl
Rbb_45_29 bitb_45_29 bitb_45_30 R_bl
Cb_45_29 bit_45_29 gnd C_bl
Cbb_45_29 bitb_45_29 gnd C_bl
Rb_45_30 bit_45_30 bit_45_31 R_bl
Rbb_45_30 bitb_45_30 bitb_45_31 R_bl
Cb_45_30 bit_45_30 gnd C_bl
Cbb_45_30 bitb_45_30 gnd C_bl
Rb_45_31 bit_45_31 bit_45_32 R_bl
Rbb_45_31 bitb_45_31 bitb_45_32 R_bl
Cb_45_31 bit_45_31 gnd C_bl
Cbb_45_31 bitb_45_31 gnd C_bl
Rb_45_32 bit_45_32 bit_45_33 R_bl
Rbb_45_32 bitb_45_32 bitb_45_33 R_bl
Cb_45_32 bit_45_32 gnd C_bl
Cbb_45_32 bitb_45_32 gnd C_bl
Rb_45_33 bit_45_33 bit_45_34 R_bl
Rbb_45_33 bitb_45_33 bitb_45_34 R_bl
Cb_45_33 bit_45_33 gnd C_bl
Cbb_45_33 bitb_45_33 gnd C_bl
Rb_45_34 bit_45_34 bit_45_35 R_bl
Rbb_45_34 bitb_45_34 bitb_45_35 R_bl
Cb_45_34 bit_45_34 gnd C_bl
Cbb_45_34 bitb_45_34 gnd C_bl
Rb_45_35 bit_45_35 bit_45_36 R_bl
Rbb_45_35 bitb_45_35 bitb_45_36 R_bl
Cb_45_35 bit_45_35 gnd C_bl
Cbb_45_35 bitb_45_35 gnd C_bl
Rb_45_36 bit_45_36 bit_45_37 R_bl
Rbb_45_36 bitb_45_36 bitb_45_37 R_bl
Cb_45_36 bit_45_36 gnd C_bl
Cbb_45_36 bitb_45_36 gnd C_bl
Rb_45_37 bit_45_37 bit_45_38 R_bl
Rbb_45_37 bitb_45_37 bitb_45_38 R_bl
Cb_45_37 bit_45_37 gnd C_bl
Cbb_45_37 bitb_45_37 gnd C_bl
Rb_45_38 bit_45_38 bit_45_39 R_bl
Rbb_45_38 bitb_45_38 bitb_45_39 R_bl
Cb_45_38 bit_45_38 gnd C_bl
Cbb_45_38 bitb_45_38 gnd C_bl
Rb_45_39 bit_45_39 bit_45_40 R_bl
Rbb_45_39 bitb_45_39 bitb_45_40 R_bl
Cb_45_39 bit_45_39 gnd C_bl
Cbb_45_39 bitb_45_39 gnd C_bl
Rb_45_40 bit_45_40 bit_45_41 R_bl
Rbb_45_40 bitb_45_40 bitb_45_41 R_bl
Cb_45_40 bit_45_40 gnd C_bl
Cbb_45_40 bitb_45_40 gnd C_bl
Rb_45_41 bit_45_41 bit_45_42 R_bl
Rbb_45_41 bitb_45_41 bitb_45_42 R_bl
Cb_45_41 bit_45_41 gnd C_bl
Cbb_45_41 bitb_45_41 gnd C_bl
Rb_45_42 bit_45_42 bit_45_43 R_bl
Rbb_45_42 bitb_45_42 bitb_45_43 R_bl
Cb_45_42 bit_45_42 gnd C_bl
Cbb_45_42 bitb_45_42 gnd C_bl
Rb_45_43 bit_45_43 bit_45_44 R_bl
Rbb_45_43 bitb_45_43 bitb_45_44 R_bl
Cb_45_43 bit_45_43 gnd C_bl
Cbb_45_43 bitb_45_43 gnd C_bl
Rb_45_44 bit_45_44 bit_45_45 R_bl
Rbb_45_44 bitb_45_44 bitb_45_45 R_bl
Cb_45_44 bit_45_44 gnd C_bl
Cbb_45_44 bitb_45_44 gnd C_bl
Rb_45_45 bit_45_45 bit_45_46 R_bl
Rbb_45_45 bitb_45_45 bitb_45_46 R_bl
Cb_45_45 bit_45_45 gnd C_bl
Cbb_45_45 bitb_45_45 gnd C_bl
Rb_45_46 bit_45_46 bit_45_47 R_bl
Rbb_45_46 bitb_45_46 bitb_45_47 R_bl
Cb_45_46 bit_45_46 gnd C_bl
Cbb_45_46 bitb_45_46 gnd C_bl
Rb_45_47 bit_45_47 bit_45_48 R_bl
Rbb_45_47 bitb_45_47 bitb_45_48 R_bl
Cb_45_47 bit_45_47 gnd C_bl
Cbb_45_47 bitb_45_47 gnd C_bl
Rb_45_48 bit_45_48 bit_45_49 R_bl
Rbb_45_48 bitb_45_48 bitb_45_49 R_bl
Cb_45_48 bit_45_48 gnd C_bl
Cbb_45_48 bitb_45_48 gnd C_bl
Rb_45_49 bit_45_49 bit_45_50 R_bl
Rbb_45_49 bitb_45_49 bitb_45_50 R_bl
Cb_45_49 bit_45_49 gnd C_bl
Cbb_45_49 bitb_45_49 gnd C_bl
Rb_45_50 bit_45_50 bit_45_51 R_bl
Rbb_45_50 bitb_45_50 bitb_45_51 R_bl
Cb_45_50 bit_45_50 gnd C_bl
Cbb_45_50 bitb_45_50 gnd C_bl
Rb_45_51 bit_45_51 bit_45_52 R_bl
Rbb_45_51 bitb_45_51 bitb_45_52 R_bl
Cb_45_51 bit_45_51 gnd C_bl
Cbb_45_51 bitb_45_51 gnd C_bl
Rb_45_52 bit_45_52 bit_45_53 R_bl
Rbb_45_52 bitb_45_52 bitb_45_53 R_bl
Cb_45_52 bit_45_52 gnd C_bl
Cbb_45_52 bitb_45_52 gnd C_bl
Rb_45_53 bit_45_53 bit_45_54 R_bl
Rbb_45_53 bitb_45_53 bitb_45_54 R_bl
Cb_45_53 bit_45_53 gnd C_bl
Cbb_45_53 bitb_45_53 gnd C_bl
Rb_45_54 bit_45_54 bit_45_55 R_bl
Rbb_45_54 bitb_45_54 bitb_45_55 R_bl
Cb_45_54 bit_45_54 gnd C_bl
Cbb_45_54 bitb_45_54 gnd C_bl
Rb_45_55 bit_45_55 bit_45_56 R_bl
Rbb_45_55 bitb_45_55 bitb_45_56 R_bl
Cb_45_55 bit_45_55 gnd C_bl
Cbb_45_55 bitb_45_55 gnd C_bl
Rb_45_56 bit_45_56 bit_45_57 R_bl
Rbb_45_56 bitb_45_56 bitb_45_57 R_bl
Cb_45_56 bit_45_56 gnd C_bl
Cbb_45_56 bitb_45_56 gnd C_bl
Rb_45_57 bit_45_57 bit_45_58 R_bl
Rbb_45_57 bitb_45_57 bitb_45_58 R_bl
Cb_45_57 bit_45_57 gnd C_bl
Cbb_45_57 bitb_45_57 gnd C_bl
Rb_45_58 bit_45_58 bit_45_59 R_bl
Rbb_45_58 bitb_45_58 bitb_45_59 R_bl
Cb_45_58 bit_45_58 gnd C_bl
Cbb_45_58 bitb_45_58 gnd C_bl
Rb_45_59 bit_45_59 bit_45_60 R_bl
Rbb_45_59 bitb_45_59 bitb_45_60 R_bl
Cb_45_59 bit_45_59 gnd C_bl
Cbb_45_59 bitb_45_59 gnd C_bl
Rb_45_60 bit_45_60 bit_45_61 R_bl
Rbb_45_60 bitb_45_60 bitb_45_61 R_bl
Cb_45_60 bit_45_60 gnd C_bl
Cbb_45_60 bitb_45_60 gnd C_bl
Rb_45_61 bit_45_61 bit_45_62 R_bl
Rbb_45_61 bitb_45_61 bitb_45_62 R_bl
Cb_45_61 bit_45_61 gnd C_bl
Cbb_45_61 bitb_45_61 gnd C_bl
Rb_45_62 bit_45_62 bit_45_63 R_bl
Rbb_45_62 bitb_45_62 bitb_45_63 R_bl
Cb_45_62 bit_45_62 gnd C_bl
Cbb_45_62 bitb_45_62 gnd C_bl
Rb_45_63 bit_45_63 bit_45_64 R_bl
Rbb_45_63 bitb_45_63 bitb_45_64 R_bl
Cb_45_63 bit_45_63 gnd C_bl
Cbb_45_63 bitb_45_63 gnd C_bl
Rb_45_64 bit_45_64 bit_45_65 R_bl
Rbb_45_64 bitb_45_64 bitb_45_65 R_bl
Cb_45_64 bit_45_64 gnd C_bl
Cbb_45_64 bitb_45_64 gnd C_bl
Rb_45_65 bit_45_65 bit_45_66 R_bl
Rbb_45_65 bitb_45_65 bitb_45_66 R_bl
Cb_45_65 bit_45_65 gnd C_bl
Cbb_45_65 bitb_45_65 gnd C_bl
Rb_45_66 bit_45_66 bit_45_67 R_bl
Rbb_45_66 bitb_45_66 bitb_45_67 R_bl
Cb_45_66 bit_45_66 gnd C_bl
Cbb_45_66 bitb_45_66 gnd C_bl
Rb_45_67 bit_45_67 bit_45_68 R_bl
Rbb_45_67 bitb_45_67 bitb_45_68 R_bl
Cb_45_67 bit_45_67 gnd C_bl
Cbb_45_67 bitb_45_67 gnd C_bl
Rb_45_68 bit_45_68 bit_45_69 R_bl
Rbb_45_68 bitb_45_68 bitb_45_69 R_bl
Cb_45_68 bit_45_68 gnd C_bl
Cbb_45_68 bitb_45_68 gnd C_bl
Rb_45_69 bit_45_69 bit_45_70 R_bl
Rbb_45_69 bitb_45_69 bitb_45_70 R_bl
Cb_45_69 bit_45_69 gnd C_bl
Cbb_45_69 bitb_45_69 gnd C_bl
Rb_45_70 bit_45_70 bit_45_71 R_bl
Rbb_45_70 bitb_45_70 bitb_45_71 R_bl
Cb_45_70 bit_45_70 gnd C_bl
Cbb_45_70 bitb_45_70 gnd C_bl
Rb_45_71 bit_45_71 bit_45_72 R_bl
Rbb_45_71 bitb_45_71 bitb_45_72 R_bl
Cb_45_71 bit_45_71 gnd C_bl
Cbb_45_71 bitb_45_71 gnd C_bl
Rb_45_72 bit_45_72 bit_45_73 R_bl
Rbb_45_72 bitb_45_72 bitb_45_73 R_bl
Cb_45_72 bit_45_72 gnd C_bl
Cbb_45_72 bitb_45_72 gnd C_bl
Rb_45_73 bit_45_73 bit_45_74 R_bl
Rbb_45_73 bitb_45_73 bitb_45_74 R_bl
Cb_45_73 bit_45_73 gnd C_bl
Cbb_45_73 bitb_45_73 gnd C_bl
Rb_45_74 bit_45_74 bit_45_75 R_bl
Rbb_45_74 bitb_45_74 bitb_45_75 R_bl
Cb_45_74 bit_45_74 gnd C_bl
Cbb_45_74 bitb_45_74 gnd C_bl
Rb_45_75 bit_45_75 bit_45_76 R_bl
Rbb_45_75 bitb_45_75 bitb_45_76 R_bl
Cb_45_75 bit_45_75 gnd C_bl
Cbb_45_75 bitb_45_75 gnd C_bl
Rb_45_76 bit_45_76 bit_45_77 R_bl
Rbb_45_76 bitb_45_76 bitb_45_77 R_bl
Cb_45_76 bit_45_76 gnd C_bl
Cbb_45_76 bitb_45_76 gnd C_bl
Rb_45_77 bit_45_77 bit_45_78 R_bl
Rbb_45_77 bitb_45_77 bitb_45_78 R_bl
Cb_45_77 bit_45_77 gnd C_bl
Cbb_45_77 bitb_45_77 gnd C_bl
Rb_45_78 bit_45_78 bit_45_79 R_bl
Rbb_45_78 bitb_45_78 bitb_45_79 R_bl
Cb_45_78 bit_45_78 gnd C_bl
Cbb_45_78 bitb_45_78 gnd C_bl
Rb_45_79 bit_45_79 bit_45_80 R_bl
Rbb_45_79 bitb_45_79 bitb_45_80 R_bl
Cb_45_79 bit_45_79 gnd C_bl
Cbb_45_79 bitb_45_79 gnd C_bl
Rb_45_80 bit_45_80 bit_45_81 R_bl
Rbb_45_80 bitb_45_80 bitb_45_81 R_bl
Cb_45_80 bit_45_80 gnd C_bl
Cbb_45_80 bitb_45_80 gnd C_bl
Rb_45_81 bit_45_81 bit_45_82 R_bl
Rbb_45_81 bitb_45_81 bitb_45_82 R_bl
Cb_45_81 bit_45_81 gnd C_bl
Cbb_45_81 bitb_45_81 gnd C_bl
Rb_45_82 bit_45_82 bit_45_83 R_bl
Rbb_45_82 bitb_45_82 bitb_45_83 R_bl
Cb_45_82 bit_45_82 gnd C_bl
Cbb_45_82 bitb_45_82 gnd C_bl
Rb_45_83 bit_45_83 bit_45_84 R_bl
Rbb_45_83 bitb_45_83 bitb_45_84 R_bl
Cb_45_83 bit_45_83 gnd C_bl
Cbb_45_83 bitb_45_83 gnd C_bl
Rb_45_84 bit_45_84 bit_45_85 R_bl
Rbb_45_84 bitb_45_84 bitb_45_85 R_bl
Cb_45_84 bit_45_84 gnd C_bl
Cbb_45_84 bitb_45_84 gnd C_bl
Rb_45_85 bit_45_85 bit_45_86 R_bl
Rbb_45_85 bitb_45_85 bitb_45_86 R_bl
Cb_45_85 bit_45_85 gnd C_bl
Cbb_45_85 bitb_45_85 gnd C_bl
Rb_45_86 bit_45_86 bit_45_87 R_bl
Rbb_45_86 bitb_45_86 bitb_45_87 R_bl
Cb_45_86 bit_45_86 gnd C_bl
Cbb_45_86 bitb_45_86 gnd C_bl
Rb_45_87 bit_45_87 bit_45_88 R_bl
Rbb_45_87 bitb_45_87 bitb_45_88 R_bl
Cb_45_87 bit_45_87 gnd C_bl
Cbb_45_87 bitb_45_87 gnd C_bl
Rb_45_88 bit_45_88 bit_45_89 R_bl
Rbb_45_88 bitb_45_88 bitb_45_89 R_bl
Cb_45_88 bit_45_88 gnd C_bl
Cbb_45_88 bitb_45_88 gnd C_bl
Rb_45_89 bit_45_89 bit_45_90 R_bl
Rbb_45_89 bitb_45_89 bitb_45_90 R_bl
Cb_45_89 bit_45_89 gnd C_bl
Cbb_45_89 bitb_45_89 gnd C_bl
Rb_45_90 bit_45_90 bit_45_91 R_bl
Rbb_45_90 bitb_45_90 bitb_45_91 R_bl
Cb_45_90 bit_45_90 gnd C_bl
Cbb_45_90 bitb_45_90 gnd C_bl
Rb_45_91 bit_45_91 bit_45_92 R_bl
Rbb_45_91 bitb_45_91 bitb_45_92 R_bl
Cb_45_91 bit_45_91 gnd C_bl
Cbb_45_91 bitb_45_91 gnd C_bl
Rb_45_92 bit_45_92 bit_45_93 R_bl
Rbb_45_92 bitb_45_92 bitb_45_93 R_bl
Cb_45_92 bit_45_92 gnd C_bl
Cbb_45_92 bitb_45_92 gnd C_bl
Rb_45_93 bit_45_93 bit_45_94 R_bl
Rbb_45_93 bitb_45_93 bitb_45_94 R_bl
Cb_45_93 bit_45_93 gnd C_bl
Cbb_45_93 bitb_45_93 gnd C_bl
Rb_45_94 bit_45_94 bit_45_95 R_bl
Rbb_45_94 bitb_45_94 bitb_45_95 R_bl
Cb_45_94 bit_45_94 gnd C_bl
Cbb_45_94 bitb_45_94 gnd C_bl
Rb_45_95 bit_45_95 bit_45_96 R_bl
Rbb_45_95 bitb_45_95 bitb_45_96 R_bl
Cb_45_95 bit_45_95 gnd C_bl
Cbb_45_95 bitb_45_95 gnd C_bl
Rb_45_96 bit_45_96 bit_45_97 R_bl
Rbb_45_96 bitb_45_96 bitb_45_97 R_bl
Cb_45_96 bit_45_96 gnd C_bl
Cbb_45_96 bitb_45_96 gnd C_bl
Rb_45_97 bit_45_97 bit_45_98 R_bl
Rbb_45_97 bitb_45_97 bitb_45_98 R_bl
Cb_45_97 bit_45_97 gnd C_bl
Cbb_45_97 bitb_45_97 gnd C_bl
Rb_45_98 bit_45_98 bit_45_99 R_bl
Rbb_45_98 bitb_45_98 bitb_45_99 R_bl
Cb_45_98 bit_45_98 gnd C_bl
Cbb_45_98 bitb_45_98 gnd C_bl
Rb_45_99 bit_45_99 bit_45_100 R_bl
Rbb_45_99 bitb_45_99 bitb_45_100 R_bl
Cb_45_99 bit_45_99 gnd C_bl
Cbb_45_99 bitb_45_99 gnd C_bl
Rb_46_0 bit_46_0 bit_46_1 R_bl
Rbb_46_0 bitb_46_0 bitb_46_1 R_bl
Cb_46_0 bit_46_0 gnd C_bl
Cbb_46_0 bitb_46_0 gnd C_bl
Rb_46_1 bit_46_1 bit_46_2 R_bl
Rbb_46_1 bitb_46_1 bitb_46_2 R_bl
Cb_46_1 bit_46_1 gnd C_bl
Cbb_46_1 bitb_46_1 gnd C_bl
Rb_46_2 bit_46_2 bit_46_3 R_bl
Rbb_46_2 bitb_46_2 bitb_46_3 R_bl
Cb_46_2 bit_46_2 gnd C_bl
Cbb_46_2 bitb_46_2 gnd C_bl
Rb_46_3 bit_46_3 bit_46_4 R_bl
Rbb_46_3 bitb_46_3 bitb_46_4 R_bl
Cb_46_3 bit_46_3 gnd C_bl
Cbb_46_3 bitb_46_3 gnd C_bl
Rb_46_4 bit_46_4 bit_46_5 R_bl
Rbb_46_4 bitb_46_4 bitb_46_5 R_bl
Cb_46_4 bit_46_4 gnd C_bl
Cbb_46_4 bitb_46_4 gnd C_bl
Rb_46_5 bit_46_5 bit_46_6 R_bl
Rbb_46_5 bitb_46_5 bitb_46_6 R_bl
Cb_46_5 bit_46_5 gnd C_bl
Cbb_46_5 bitb_46_5 gnd C_bl
Rb_46_6 bit_46_6 bit_46_7 R_bl
Rbb_46_6 bitb_46_6 bitb_46_7 R_bl
Cb_46_6 bit_46_6 gnd C_bl
Cbb_46_6 bitb_46_6 gnd C_bl
Rb_46_7 bit_46_7 bit_46_8 R_bl
Rbb_46_7 bitb_46_7 bitb_46_8 R_bl
Cb_46_7 bit_46_7 gnd C_bl
Cbb_46_7 bitb_46_7 gnd C_bl
Rb_46_8 bit_46_8 bit_46_9 R_bl
Rbb_46_8 bitb_46_8 bitb_46_9 R_bl
Cb_46_8 bit_46_8 gnd C_bl
Cbb_46_8 bitb_46_8 gnd C_bl
Rb_46_9 bit_46_9 bit_46_10 R_bl
Rbb_46_9 bitb_46_9 bitb_46_10 R_bl
Cb_46_9 bit_46_9 gnd C_bl
Cbb_46_9 bitb_46_9 gnd C_bl
Rb_46_10 bit_46_10 bit_46_11 R_bl
Rbb_46_10 bitb_46_10 bitb_46_11 R_bl
Cb_46_10 bit_46_10 gnd C_bl
Cbb_46_10 bitb_46_10 gnd C_bl
Rb_46_11 bit_46_11 bit_46_12 R_bl
Rbb_46_11 bitb_46_11 bitb_46_12 R_bl
Cb_46_11 bit_46_11 gnd C_bl
Cbb_46_11 bitb_46_11 gnd C_bl
Rb_46_12 bit_46_12 bit_46_13 R_bl
Rbb_46_12 bitb_46_12 bitb_46_13 R_bl
Cb_46_12 bit_46_12 gnd C_bl
Cbb_46_12 bitb_46_12 gnd C_bl
Rb_46_13 bit_46_13 bit_46_14 R_bl
Rbb_46_13 bitb_46_13 bitb_46_14 R_bl
Cb_46_13 bit_46_13 gnd C_bl
Cbb_46_13 bitb_46_13 gnd C_bl
Rb_46_14 bit_46_14 bit_46_15 R_bl
Rbb_46_14 bitb_46_14 bitb_46_15 R_bl
Cb_46_14 bit_46_14 gnd C_bl
Cbb_46_14 bitb_46_14 gnd C_bl
Rb_46_15 bit_46_15 bit_46_16 R_bl
Rbb_46_15 bitb_46_15 bitb_46_16 R_bl
Cb_46_15 bit_46_15 gnd C_bl
Cbb_46_15 bitb_46_15 gnd C_bl
Rb_46_16 bit_46_16 bit_46_17 R_bl
Rbb_46_16 bitb_46_16 bitb_46_17 R_bl
Cb_46_16 bit_46_16 gnd C_bl
Cbb_46_16 bitb_46_16 gnd C_bl
Rb_46_17 bit_46_17 bit_46_18 R_bl
Rbb_46_17 bitb_46_17 bitb_46_18 R_bl
Cb_46_17 bit_46_17 gnd C_bl
Cbb_46_17 bitb_46_17 gnd C_bl
Rb_46_18 bit_46_18 bit_46_19 R_bl
Rbb_46_18 bitb_46_18 bitb_46_19 R_bl
Cb_46_18 bit_46_18 gnd C_bl
Cbb_46_18 bitb_46_18 gnd C_bl
Rb_46_19 bit_46_19 bit_46_20 R_bl
Rbb_46_19 bitb_46_19 bitb_46_20 R_bl
Cb_46_19 bit_46_19 gnd C_bl
Cbb_46_19 bitb_46_19 gnd C_bl
Rb_46_20 bit_46_20 bit_46_21 R_bl
Rbb_46_20 bitb_46_20 bitb_46_21 R_bl
Cb_46_20 bit_46_20 gnd C_bl
Cbb_46_20 bitb_46_20 gnd C_bl
Rb_46_21 bit_46_21 bit_46_22 R_bl
Rbb_46_21 bitb_46_21 bitb_46_22 R_bl
Cb_46_21 bit_46_21 gnd C_bl
Cbb_46_21 bitb_46_21 gnd C_bl
Rb_46_22 bit_46_22 bit_46_23 R_bl
Rbb_46_22 bitb_46_22 bitb_46_23 R_bl
Cb_46_22 bit_46_22 gnd C_bl
Cbb_46_22 bitb_46_22 gnd C_bl
Rb_46_23 bit_46_23 bit_46_24 R_bl
Rbb_46_23 bitb_46_23 bitb_46_24 R_bl
Cb_46_23 bit_46_23 gnd C_bl
Cbb_46_23 bitb_46_23 gnd C_bl
Rb_46_24 bit_46_24 bit_46_25 R_bl
Rbb_46_24 bitb_46_24 bitb_46_25 R_bl
Cb_46_24 bit_46_24 gnd C_bl
Cbb_46_24 bitb_46_24 gnd C_bl
Rb_46_25 bit_46_25 bit_46_26 R_bl
Rbb_46_25 bitb_46_25 bitb_46_26 R_bl
Cb_46_25 bit_46_25 gnd C_bl
Cbb_46_25 bitb_46_25 gnd C_bl
Rb_46_26 bit_46_26 bit_46_27 R_bl
Rbb_46_26 bitb_46_26 bitb_46_27 R_bl
Cb_46_26 bit_46_26 gnd C_bl
Cbb_46_26 bitb_46_26 gnd C_bl
Rb_46_27 bit_46_27 bit_46_28 R_bl
Rbb_46_27 bitb_46_27 bitb_46_28 R_bl
Cb_46_27 bit_46_27 gnd C_bl
Cbb_46_27 bitb_46_27 gnd C_bl
Rb_46_28 bit_46_28 bit_46_29 R_bl
Rbb_46_28 bitb_46_28 bitb_46_29 R_bl
Cb_46_28 bit_46_28 gnd C_bl
Cbb_46_28 bitb_46_28 gnd C_bl
Rb_46_29 bit_46_29 bit_46_30 R_bl
Rbb_46_29 bitb_46_29 bitb_46_30 R_bl
Cb_46_29 bit_46_29 gnd C_bl
Cbb_46_29 bitb_46_29 gnd C_bl
Rb_46_30 bit_46_30 bit_46_31 R_bl
Rbb_46_30 bitb_46_30 bitb_46_31 R_bl
Cb_46_30 bit_46_30 gnd C_bl
Cbb_46_30 bitb_46_30 gnd C_bl
Rb_46_31 bit_46_31 bit_46_32 R_bl
Rbb_46_31 bitb_46_31 bitb_46_32 R_bl
Cb_46_31 bit_46_31 gnd C_bl
Cbb_46_31 bitb_46_31 gnd C_bl
Rb_46_32 bit_46_32 bit_46_33 R_bl
Rbb_46_32 bitb_46_32 bitb_46_33 R_bl
Cb_46_32 bit_46_32 gnd C_bl
Cbb_46_32 bitb_46_32 gnd C_bl
Rb_46_33 bit_46_33 bit_46_34 R_bl
Rbb_46_33 bitb_46_33 bitb_46_34 R_bl
Cb_46_33 bit_46_33 gnd C_bl
Cbb_46_33 bitb_46_33 gnd C_bl
Rb_46_34 bit_46_34 bit_46_35 R_bl
Rbb_46_34 bitb_46_34 bitb_46_35 R_bl
Cb_46_34 bit_46_34 gnd C_bl
Cbb_46_34 bitb_46_34 gnd C_bl
Rb_46_35 bit_46_35 bit_46_36 R_bl
Rbb_46_35 bitb_46_35 bitb_46_36 R_bl
Cb_46_35 bit_46_35 gnd C_bl
Cbb_46_35 bitb_46_35 gnd C_bl
Rb_46_36 bit_46_36 bit_46_37 R_bl
Rbb_46_36 bitb_46_36 bitb_46_37 R_bl
Cb_46_36 bit_46_36 gnd C_bl
Cbb_46_36 bitb_46_36 gnd C_bl
Rb_46_37 bit_46_37 bit_46_38 R_bl
Rbb_46_37 bitb_46_37 bitb_46_38 R_bl
Cb_46_37 bit_46_37 gnd C_bl
Cbb_46_37 bitb_46_37 gnd C_bl
Rb_46_38 bit_46_38 bit_46_39 R_bl
Rbb_46_38 bitb_46_38 bitb_46_39 R_bl
Cb_46_38 bit_46_38 gnd C_bl
Cbb_46_38 bitb_46_38 gnd C_bl
Rb_46_39 bit_46_39 bit_46_40 R_bl
Rbb_46_39 bitb_46_39 bitb_46_40 R_bl
Cb_46_39 bit_46_39 gnd C_bl
Cbb_46_39 bitb_46_39 gnd C_bl
Rb_46_40 bit_46_40 bit_46_41 R_bl
Rbb_46_40 bitb_46_40 bitb_46_41 R_bl
Cb_46_40 bit_46_40 gnd C_bl
Cbb_46_40 bitb_46_40 gnd C_bl
Rb_46_41 bit_46_41 bit_46_42 R_bl
Rbb_46_41 bitb_46_41 bitb_46_42 R_bl
Cb_46_41 bit_46_41 gnd C_bl
Cbb_46_41 bitb_46_41 gnd C_bl
Rb_46_42 bit_46_42 bit_46_43 R_bl
Rbb_46_42 bitb_46_42 bitb_46_43 R_bl
Cb_46_42 bit_46_42 gnd C_bl
Cbb_46_42 bitb_46_42 gnd C_bl
Rb_46_43 bit_46_43 bit_46_44 R_bl
Rbb_46_43 bitb_46_43 bitb_46_44 R_bl
Cb_46_43 bit_46_43 gnd C_bl
Cbb_46_43 bitb_46_43 gnd C_bl
Rb_46_44 bit_46_44 bit_46_45 R_bl
Rbb_46_44 bitb_46_44 bitb_46_45 R_bl
Cb_46_44 bit_46_44 gnd C_bl
Cbb_46_44 bitb_46_44 gnd C_bl
Rb_46_45 bit_46_45 bit_46_46 R_bl
Rbb_46_45 bitb_46_45 bitb_46_46 R_bl
Cb_46_45 bit_46_45 gnd C_bl
Cbb_46_45 bitb_46_45 gnd C_bl
Rb_46_46 bit_46_46 bit_46_47 R_bl
Rbb_46_46 bitb_46_46 bitb_46_47 R_bl
Cb_46_46 bit_46_46 gnd C_bl
Cbb_46_46 bitb_46_46 gnd C_bl
Rb_46_47 bit_46_47 bit_46_48 R_bl
Rbb_46_47 bitb_46_47 bitb_46_48 R_bl
Cb_46_47 bit_46_47 gnd C_bl
Cbb_46_47 bitb_46_47 gnd C_bl
Rb_46_48 bit_46_48 bit_46_49 R_bl
Rbb_46_48 bitb_46_48 bitb_46_49 R_bl
Cb_46_48 bit_46_48 gnd C_bl
Cbb_46_48 bitb_46_48 gnd C_bl
Rb_46_49 bit_46_49 bit_46_50 R_bl
Rbb_46_49 bitb_46_49 bitb_46_50 R_bl
Cb_46_49 bit_46_49 gnd C_bl
Cbb_46_49 bitb_46_49 gnd C_bl
Rb_46_50 bit_46_50 bit_46_51 R_bl
Rbb_46_50 bitb_46_50 bitb_46_51 R_bl
Cb_46_50 bit_46_50 gnd C_bl
Cbb_46_50 bitb_46_50 gnd C_bl
Rb_46_51 bit_46_51 bit_46_52 R_bl
Rbb_46_51 bitb_46_51 bitb_46_52 R_bl
Cb_46_51 bit_46_51 gnd C_bl
Cbb_46_51 bitb_46_51 gnd C_bl
Rb_46_52 bit_46_52 bit_46_53 R_bl
Rbb_46_52 bitb_46_52 bitb_46_53 R_bl
Cb_46_52 bit_46_52 gnd C_bl
Cbb_46_52 bitb_46_52 gnd C_bl
Rb_46_53 bit_46_53 bit_46_54 R_bl
Rbb_46_53 bitb_46_53 bitb_46_54 R_bl
Cb_46_53 bit_46_53 gnd C_bl
Cbb_46_53 bitb_46_53 gnd C_bl
Rb_46_54 bit_46_54 bit_46_55 R_bl
Rbb_46_54 bitb_46_54 bitb_46_55 R_bl
Cb_46_54 bit_46_54 gnd C_bl
Cbb_46_54 bitb_46_54 gnd C_bl
Rb_46_55 bit_46_55 bit_46_56 R_bl
Rbb_46_55 bitb_46_55 bitb_46_56 R_bl
Cb_46_55 bit_46_55 gnd C_bl
Cbb_46_55 bitb_46_55 gnd C_bl
Rb_46_56 bit_46_56 bit_46_57 R_bl
Rbb_46_56 bitb_46_56 bitb_46_57 R_bl
Cb_46_56 bit_46_56 gnd C_bl
Cbb_46_56 bitb_46_56 gnd C_bl
Rb_46_57 bit_46_57 bit_46_58 R_bl
Rbb_46_57 bitb_46_57 bitb_46_58 R_bl
Cb_46_57 bit_46_57 gnd C_bl
Cbb_46_57 bitb_46_57 gnd C_bl
Rb_46_58 bit_46_58 bit_46_59 R_bl
Rbb_46_58 bitb_46_58 bitb_46_59 R_bl
Cb_46_58 bit_46_58 gnd C_bl
Cbb_46_58 bitb_46_58 gnd C_bl
Rb_46_59 bit_46_59 bit_46_60 R_bl
Rbb_46_59 bitb_46_59 bitb_46_60 R_bl
Cb_46_59 bit_46_59 gnd C_bl
Cbb_46_59 bitb_46_59 gnd C_bl
Rb_46_60 bit_46_60 bit_46_61 R_bl
Rbb_46_60 bitb_46_60 bitb_46_61 R_bl
Cb_46_60 bit_46_60 gnd C_bl
Cbb_46_60 bitb_46_60 gnd C_bl
Rb_46_61 bit_46_61 bit_46_62 R_bl
Rbb_46_61 bitb_46_61 bitb_46_62 R_bl
Cb_46_61 bit_46_61 gnd C_bl
Cbb_46_61 bitb_46_61 gnd C_bl
Rb_46_62 bit_46_62 bit_46_63 R_bl
Rbb_46_62 bitb_46_62 bitb_46_63 R_bl
Cb_46_62 bit_46_62 gnd C_bl
Cbb_46_62 bitb_46_62 gnd C_bl
Rb_46_63 bit_46_63 bit_46_64 R_bl
Rbb_46_63 bitb_46_63 bitb_46_64 R_bl
Cb_46_63 bit_46_63 gnd C_bl
Cbb_46_63 bitb_46_63 gnd C_bl
Rb_46_64 bit_46_64 bit_46_65 R_bl
Rbb_46_64 bitb_46_64 bitb_46_65 R_bl
Cb_46_64 bit_46_64 gnd C_bl
Cbb_46_64 bitb_46_64 gnd C_bl
Rb_46_65 bit_46_65 bit_46_66 R_bl
Rbb_46_65 bitb_46_65 bitb_46_66 R_bl
Cb_46_65 bit_46_65 gnd C_bl
Cbb_46_65 bitb_46_65 gnd C_bl
Rb_46_66 bit_46_66 bit_46_67 R_bl
Rbb_46_66 bitb_46_66 bitb_46_67 R_bl
Cb_46_66 bit_46_66 gnd C_bl
Cbb_46_66 bitb_46_66 gnd C_bl
Rb_46_67 bit_46_67 bit_46_68 R_bl
Rbb_46_67 bitb_46_67 bitb_46_68 R_bl
Cb_46_67 bit_46_67 gnd C_bl
Cbb_46_67 bitb_46_67 gnd C_bl
Rb_46_68 bit_46_68 bit_46_69 R_bl
Rbb_46_68 bitb_46_68 bitb_46_69 R_bl
Cb_46_68 bit_46_68 gnd C_bl
Cbb_46_68 bitb_46_68 gnd C_bl
Rb_46_69 bit_46_69 bit_46_70 R_bl
Rbb_46_69 bitb_46_69 bitb_46_70 R_bl
Cb_46_69 bit_46_69 gnd C_bl
Cbb_46_69 bitb_46_69 gnd C_bl
Rb_46_70 bit_46_70 bit_46_71 R_bl
Rbb_46_70 bitb_46_70 bitb_46_71 R_bl
Cb_46_70 bit_46_70 gnd C_bl
Cbb_46_70 bitb_46_70 gnd C_bl
Rb_46_71 bit_46_71 bit_46_72 R_bl
Rbb_46_71 bitb_46_71 bitb_46_72 R_bl
Cb_46_71 bit_46_71 gnd C_bl
Cbb_46_71 bitb_46_71 gnd C_bl
Rb_46_72 bit_46_72 bit_46_73 R_bl
Rbb_46_72 bitb_46_72 bitb_46_73 R_bl
Cb_46_72 bit_46_72 gnd C_bl
Cbb_46_72 bitb_46_72 gnd C_bl
Rb_46_73 bit_46_73 bit_46_74 R_bl
Rbb_46_73 bitb_46_73 bitb_46_74 R_bl
Cb_46_73 bit_46_73 gnd C_bl
Cbb_46_73 bitb_46_73 gnd C_bl
Rb_46_74 bit_46_74 bit_46_75 R_bl
Rbb_46_74 bitb_46_74 bitb_46_75 R_bl
Cb_46_74 bit_46_74 gnd C_bl
Cbb_46_74 bitb_46_74 gnd C_bl
Rb_46_75 bit_46_75 bit_46_76 R_bl
Rbb_46_75 bitb_46_75 bitb_46_76 R_bl
Cb_46_75 bit_46_75 gnd C_bl
Cbb_46_75 bitb_46_75 gnd C_bl
Rb_46_76 bit_46_76 bit_46_77 R_bl
Rbb_46_76 bitb_46_76 bitb_46_77 R_bl
Cb_46_76 bit_46_76 gnd C_bl
Cbb_46_76 bitb_46_76 gnd C_bl
Rb_46_77 bit_46_77 bit_46_78 R_bl
Rbb_46_77 bitb_46_77 bitb_46_78 R_bl
Cb_46_77 bit_46_77 gnd C_bl
Cbb_46_77 bitb_46_77 gnd C_bl
Rb_46_78 bit_46_78 bit_46_79 R_bl
Rbb_46_78 bitb_46_78 bitb_46_79 R_bl
Cb_46_78 bit_46_78 gnd C_bl
Cbb_46_78 bitb_46_78 gnd C_bl
Rb_46_79 bit_46_79 bit_46_80 R_bl
Rbb_46_79 bitb_46_79 bitb_46_80 R_bl
Cb_46_79 bit_46_79 gnd C_bl
Cbb_46_79 bitb_46_79 gnd C_bl
Rb_46_80 bit_46_80 bit_46_81 R_bl
Rbb_46_80 bitb_46_80 bitb_46_81 R_bl
Cb_46_80 bit_46_80 gnd C_bl
Cbb_46_80 bitb_46_80 gnd C_bl
Rb_46_81 bit_46_81 bit_46_82 R_bl
Rbb_46_81 bitb_46_81 bitb_46_82 R_bl
Cb_46_81 bit_46_81 gnd C_bl
Cbb_46_81 bitb_46_81 gnd C_bl
Rb_46_82 bit_46_82 bit_46_83 R_bl
Rbb_46_82 bitb_46_82 bitb_46_83 R_bl
Cb_46_82 bit_46_82 gnd C_bl
Cbb_46_82 bitb_46_82 gnd C_bl
Rb_46_83 bit_46_83 bit_46_84 R_bl
Rbb_46_83 bitb_46_83 bitb_46_84 R_bl
Cb_46_83 bit_46_83 gnd C_bl
Cbb_46_83 bitb_46_83 gnd C_bl
Rb_46_84 bit_46_84 bit_46_85 R_bl
Rbb_46_84 bitb_46_84 bitb_46_85 R_bl
Cb_46_84 bit_46_84 gnd C_bl
Cbb_46_84 bitb_46_84 gnd C_bl
Rb_46_85 bit_46_85 bit_46_86 R_bl
Rbb_46_85 bitb_46_85 bitb_46_86 R_bl
Cb_46_85 bit_46_85 gnd C_bl
Cbb_46_85 bitb_46_85 gnd C_bl
Rb_46_86 bit_46_86 bit_46_87 R_bl
Rbb_46_86 bitb_46_86 bitb_46_87 R_bl
Cb_46_86 bit_46_86 gnd C_bl
Cbb_46_86 bitb_46_86 gnd C_bl
Rb_46_87 bit_46_87 bit_46_88 R_bl
Rbb_46_87 bitb_46_87 bitb_46_88 R_bl
Cb_46_87 bit_46_87 gnd C_bl
Cbb_46_87 bitb_46_87 gnd C_bl
Rb_46_88 bit_46_88 bit_46_89 R_bl
Rbb_46_88 bitb_46_88 bitb_46_89 R_bl
Cb_46_88 bit_46_88 gnd C_bl
Cbb_46_88 bitb_46_88 gnd C_bl
Rb_46_89 bit_46_89 bit_46_90 R_bl
Rbb_46_89 bitb_46_89 bitb_46_90 R_bl
Cb_46_89 bit_46_89 gnd C_bl
Cbb_46_89 bitb_46_89 gnd C_bl
Rb_46_90 bit_46_90 bit_46_91 R_bl
Rbb_46_90 bitb_46_90 bitb_46_91 R_bl
Cb_46_90 bit_46_90 gnd C_bl
Cbb_46_90 bitb_46_90 gnd C_bl
Rb_46_91 bit_46_91 bit_46_92 R_bl
Rbb_46_91 bitb_46_91 bitb_46_92 R_bl
Cb_46_91 bit_46_91 gnd C_bl
Cbb_46_91 bitb_46_91 gnd C_bl
Rb_46_92 bit_46_92 bit_46_93 R_bl
Rbb_46_92 bitb_46_92 bitb_46_93 R_bl
Cb_46_92 bit_46_92 gnd C_bl
Cbb_46_92 bitb_46_92 gnd C_bl
Rb_46_93 bit_46_93 bit_46_94 R_bl
Rbb_46_93 bitb_46_93 bitb_46_94 R_bl
Cb_46_93 bit_46_93 gnd C_bl
Cbb_46_93 bitb_46_93 gnd C_bl
Rb_46_94 bit_46_94 bit_46_95 R_bl
Rbb_46_94 bitb_46_94 bitb_46_95 R_bl
Cb_46_94 bit_46_94 gnd C_bl
Cbb_46_94 bitb_46_94 gnd C_bl
Rb_46_95 bit_46_95 bit_46_96 R_bl
Rbb_46_95 bitb_46_95 bitb_46_96 R_bl
Cb_46_95 bit_46_95 gnd C_bl
Cbb_46_95 bitb_46_95 gnd C_bl
Rb_46_96 bit_46_96 bit_46_97 R_bl
Rbb_46_96 bitb_46_96 bitb_46_97 R_bl
Cb_46_96 bit_46_96 gnd C_bl
Cbb_46_96 bitb_46_96 gnd C_bl
Rb_46_97 bit_46_97 bit_46_98 R_bl
Rbb_46_97 bitb_46_97 bitb_46_98 R_bl
Cb_46_97 bit_46_97 gnd C_bl
Cbb_46_97 bitb_46_97 gnd C_bl
Rb_46_98 bit_46_98 bit_46_99 R_bl
Rbb_46_98 bitb_46_98 bitb_46_99 R_bl
Cb_46_98 bit_46_98 gnd C_bl
Cbb_46_98 bitb_46_98 gnd C_bl
Rb_46_99 bit_46_99 bit_46_100 R_bl
Rbb_46_99 bitb_46_99 bitb_46_100 R_bl
Cb_46_99 bit_46_99 gnd C_bl
Cbb_46_99 bitb_46_99 gnd C_bl
Rb_47_0 bit_47_0 bit_47_1 R_bl
Rbb_47_0 bitb_47_0 bitb_47_1 R_bl
Cb_47_0 bit_47_0 gnd C_bl
Cbb_47_0 bitb_47_0 gnd C_bl
Rb_47_1 bit_47_1 bit_47_2 R_bl
Rbb_47_1 bitb_47_1 bitb_47_2 R_bl
Cb_47_1 bit_47_1 gnd C_bl
Cbb_47_1 bitb_47_1 gnd C_bl
Rb_47_2 bit_47_2 bit_47_3 R_bl
Rbb_47_2 bitb_47_2 bitb_47_3 R_bl
Cb_47_2 bit_47_2 gnd C_bl
Cbb_47_2 bitb_47_2 gnd C_bl
Rb_47_3 bit_47_3 bit_47_4 R_bl
Rbb_47_3 bitb_47_3 bitb_47_4 R_bl
Cb_47_3 bit_47_3 gnd C_bl
Cbb_47_3 bitb_47_3 gnd C_bl
Rb_47_4 bit_47_4 bit_47_5 R_bl
Rbb_47_4 bitb_47_4 bitb_47_5 R_bl
Cb_47_4 bit_47_4 gnd C_bl
Cbb_47_4 bitb_47_4 gnd C_bl
Rb_47_5 bit_47_5 bit_47_6 R_bl
Rbb_47_5 bitb_47_5 bitb_47_6 R_bl
Cb_47_5 bit_47_5 gnd C_bl
Cbb_47_5 bitb_47_5 gnd C_bl
Rb_47_6 bit_47_6 bit_47_7 R_bl
Rbb_47_6 bitb_47_6 bitb_47_7 R_bl
Cb_47_6 bit_47_6 gnd C_bl
Cbb_47_6 bitb_47_6 gnd C_bl
Rb_47_7 bit_47_7 bit_47_8 R_bl
Rbb_47_7 bitb_47_7 bitb_47_8 R_bl
Cb_47_7 bit_47_7 gnd C_bl
Cbb_47_7 bitb_47_7 gnd C_bl
Rb_47_8 bit_47_8 bit_47_9 R_bl
Rbb_47_8 bitb_47_8 bitb_47_9 R_bl
Cb_47_8 bit_47_8 gnd C_bl
Cbb_47_8 bitb_47_8 gnd C_bl
Rb_47_9 bit_47_9 bit_47_10 R_bl
Rbb_47_9 bitb_47_9 bitb_47_10 R_bl
Cb_47_9 bit_47_9 gnd C_bl
Cbb_47_9 bitb_47_9 gnd C_bl
Rb_47_10 bit_47_10 bit_47_11 R_bl
Rbb_47_10 bitb_47_10 bitb_47_11 R_bl
Cb_47_10 bit_47_10 gnd C_bl
Cbb_47_10 bitb_47_10 gnd C_bl
Rb_47_11 bit_47_11 bit_47_12 R_bl
Rbb_47_11 bitb_47_11 bitb_47_12 R_bl
Cb_47_11 bit_47_11 gnd C_bl
Cbb_47_11 bitb_47_11 gnd C_bl
Rb_47_12 bit_47_12 bit_47_13 R_bl
Rbb_47_12 bitb_47_12 bitb_47_13 R_bl
Cb_47_12 bit_47_12 gnd C_bl
Cbb_47_12 bitb_47_12 gnd C_bl
Rb_47_13 bit_47_13 bit_47_14 R_bl
Rbb_47_13 bitb_47_13 bitb_47_14 R_bl
Cb_47_13 bit_47_13 gnd C_bl
Cbb_47_13 bitb_47_13 gnd C_bl
Rb_47_14 bit_47_14 bit_47_15 R_bl
Rbb_47_14 bitb_47_14 bitb_47_15 R_bl
Cb_47_14 bit_47_14 gnd C_bl
Cbb_47_14 bitb_47_14 gnd C_bl
Rb_47_15 bit_47_15 bit_47_16 R_bl
Rbb_47_15 bitb_47_15 bitb_47_16 R_bl
Cb_47_15 bit_47_15 gnd C_bl
Cbb_47_15 bitb_47_15 gnd C_bl
Rb_47_16 bit_47_16 bit_47_17 R_bl
Rbb_47_16 bitb_47_16 bitb_47_17 R_bl
Cb_47_16 bit_47_16 gnd C_bl
Cbb_47_16 bitb_47_16 gnd C_bl
Rb_47_17 bit_47_17 bit_47_18 R_bl
Rbb_47_17 bitb_47_17 bitb_47_18 R_bl
Cb_47_17 bit_47_17 gnd C_bl
Cbb_47_17 bitb_47_17 gnd C_bl
Rb_47_18 bit_47_18 bit_47_19 R_bl
Rbb_47_18 bitb_47_18 bitb_47_19 R_bl
Cb_47_18 bit_47_18 gnd C_bl
Cbb_47_18 bitb_47_18 gnd C_bl
Rb_47_19 bit_47_19 bit_47_20 R_bl
Rbb_47_19 bitb_47_19 bitb_47_20 R_bl
Cb_47_19 bit_47_19 gnd C_bl
Cbb_47_19 bitb_47_19 gnd C_bl
Rb_47_20 bit_47_20 bit_47_21 R_bl
Rbb_47_20 bitb_47_20 bitb_47_21 R_bl
Cb_47_20 bit_47_20 gnd C_bl
Cbb_47_20 bitb_47_20 gnd C_bl
Rb_47_21 bit_47_21 bit_47_22 R_bl
Rbb_47_21 bitb_47_21 bitb_47_22 R_bl
Cb_47_21 bit_47_21 gnd C_bl
Cbb_47_21 bitb_47_21 gnd C_bl
Rb_47_22 bit_47_22 bit_47_23 R_bl
Rbb_47_22 bitb_47_22 bitb_47_23 R_bl
Cb_47_22 bit_47_22 gnd C_bl
Cbb_47_22 bitb_47_22 gnd C_bl
Rb_47_23 bit_47_23 bit_47_24 R_bl
Rbb_47_23 bitb_47_23 bitb_47_24 R_bl
Cb_47_23 bit_47_23 gnd C_bl
Cbb_47_23 bitb_47_23 gnd C_bl
Rb_47_24 bit_47_24 bit_47_25 R_bl
Rbb_47_24 bitb_47_24 bitb_47_25 R_bl
Cb_47_24 bit_47_24 gnd C_bl
Cbb_47_24 bitb_47_24 gnd C_bl
Rb_47_25 bit_47_25 bit_47_26 R_bl
Rbb_47_25 bitb_47_25 bitb_47_26 R_bl
Cb_47_25 bit_47_25 gnd C_bl
Cbb_47_25 bitb_47_25 gnd C_bl
Rb_47_26 bit_47_26 bit_47_27 R_bl
Rbb_47_26 bitb_47_26 bitb_47_27 R_bl
Cb_47_26 bit_47_26 gnd C_bl
Cbb_47_26 bitb_47_26 gnd C_bl
Rb_47_27 bit_47_27 bit_47_28 R_bl
Rbb_47_27 bitb_47_27 bitb_47_28 R_bl
Cb_47_27 bit_47_27 gnd C_bl
Cbb_47_27 bitb_47_27 gnd C_bl
Rb_47_28 bit_47_28 bit_47_29 R_bl
Rbb_47_28 bitb_47_28 bitb_47_29 R_bl
Cb_47_28 bit_47_28 gnd C_bl
Cbb_47_28 bitb_47_28 gnd C_bl
Rb_47_29 bit_47_29 bit_47_30 R_bl
Rbb_47_29 bitb_47_29 bitb_47_30 R_bl
Cb_47_29 bit_47_29 gnd C_bl
Cbb_47_29 bitb_47_29 gnd C_bl
Rb_47_30 bit_47_30 bit_47_31 R_bl
Rbb_47_30 bitb_47_30 bitb_47_31 R_bl
Cb_47_30 bit_47_30 gnd C_bl
Cbb_47_30 bitb_47_30 gnd C_bl
Rb_47_31 bit_47_31 bit_47_32 R_bl
Rbb_47_31 bitb_47_31 bitb_47_32 R_bl
Cb_47_31 bit_47_31 gnd C_bl
Cbb_47_31 bitb_47_31 gnd C_bl
Rb_47_32 bit_47_32 bit_47_33 R_bl
Rbb_47_32 bitb_47_32 bitb_47_33 R_bl
Cb_47_32 bit_47_32 gnd C_bl
Cbb_47_32 bitb_47_32 gnd C_bl
Rb_47_33 bit_47_33 bit_47_34 R_bl
Rbb_47_33 bitb_47_33 bitb_47_34 R_bl
Cb_47_33 bit_47_33 gnd C_bl
Cbb_47_33 bitb_47_33 gnd C_bl
Rb_47_34 bit_47_34 bit_47_35 R_bl
Rbb_47_34 bitb_47_34 bitb_47_35 R_bl
Cb_47_34 bit_47_34 gnd C_bl
Cbb_47_34 bitb_47_34 gnd C_bl
Rb_47_35 bit_47_35 bit_47_36 R_bl
Rbb_47_35 bitb_47_35 bitb_47_36 R_bl
Cb_47_35 bit_47_35 gnd C_bl
Cbb_47_35 bitb_47_35 gnd C_bl
Rb_47_36 bit_47_36 bit_47_37 R_bl
Rbb_47_36 bitb_47_36 bitb_47_37 R_bl
Cb_47_36 bit_47_36 gnd C_bl
Cbb_47_36 bitb_47_36 gnd C_bl
Rb_47_37 bit_47_37 bit_47_38 R_bl
Rbb_47_37 bitb_47_37 bitb_47_38 R_bl
Cb_47_37 bit_47_37 gnd C_bl
Cbb_47_37 bitb_47_37 gnd C_bl
Rb_47_38 bit_47_38 bit_47_39 R_bl
Rbb_47_38 bitb_47_38 bitb_47_39 R_bl
Cb_47_38 bit_47_38 gnd C_bl
Cbb_47_38 bitb_47_38 gnd C_bl
Rb_47_39 bit_47_39 bit_47_40 R_bl
Rbb_47_39 bitb_47_39 bitb_47_40 R_bl
Cb_47_39 bit_47_39 gnd C_bl
Cbb_47_39 bitb_47_39 gnd C_bl
Rb_47_40 bit_47_40 bit_47_41 R_bl
Rbb_47_40 bitb_47_40 bitb_47_41 R_bl
Cb_47_40 bit_47_40 gnd C_bl
Cbb_47_40 bitb_47_40 gnd C_bl
Rb_47_41 bit_47_41 bit_47_42 R_bl
Rbb_47_41 bitb_47_41 bitb_47_42 R_bl
Cb_47_41 bit_47_41 gnd C_bl
Cbb_47_41 bitb_47_41 gnd C_bl
Rb_47_42 bit_47_42 bit_47_43 R_bl
Rbb_47_42 bitb_47_42 bitb_47_43 R_bl
Cb_47_42 bit_47_42 gnd C_bl
Cbb_47_42 bitb_47_42 gnd C_bl
Rb_47_43 bit_47_43 bit_47_44 R_bl
Rbb_47_43 bitb_47_43 bitb_47_44 R_bl
Cb_47_43 bit_47_43 gnd C_bl
Cbb_47_43 bitb_47_43 gnd C_bl
Rb_47_44 bit_47_44 bit_47_45 R_bl
Rbb_47_44 bitb_47_44 bitb_47_45 R_bl
Cb_47_44 bit_47_44 gnd C_bl
Cbb_47_44 bitb_47_44 gnd C_bl
Rb_47_45 bit_47_45 bit_47_46 R_bl
Rbb_47_45 bitb_47_45 bitb_47_46 R_bl
Cb_47_45 bit_47_45 gnd C_bl
Cbb_47_45 bitb_47_45 gnd C_bl
Rb_47_46 bit_47_46 bit_47_47 R_bl
Rbb_47_46 bitb_47_46 bitb_47_47 R_bl
Cb_47_46 bit_47_46 gnd C_bl
Cbb_47_46 bitb_47_46 gnd C_bl
Rb_47_47 bit_47_47 bit_47_48 R_bl
Rbb_47_47 bitb_47_47 bitb_47_48 R_bl
Cb_47_47 bit_47_47 gnd C_bl
Cbb_47_47 bitb_47_47 gnd C_bl
Rb_47_48 bit_47_48 bit_47_49 R_bl
Rbb_47_48 bitb_47_48 bitb_47_49 R_bl
Cb_47_48 bit_47_48 gnd C_bl
Cbb_47_48 bitb_47_48 gnd C_bl
Rb_47_49 bit_47_49 bit_47_50 R_bl
Rbb_47_49 bitb_47_49 bitb_47_50 R_bl
Cb_47_49 bit_47_49 gnd C_bl
Cbb_47_49 bitb_47_49 gnd C_bl
Rb_47_50 bit_47_50 bit_47_51 R_bl
Rbb_47_50 bitb_47_50 bitb_47_51 R_bl
Cb_47_50 bit_47_50 gnd C_bl
Cbb_47_50 bitb_47_50 gnd C_bl
Rb_47_51 bit_47_51 bit_47_52 R_bl
Rbb_47_51 bitb_47_51 bitb_47_52 R_bl
Cb_47_51 bit_47_51 gnd C_bl
Cbb_47_51 bitb_47_51 gnd C_bl
Rb_47_52 bit_47_52 bit_47_53 R_bl
Rbb_47_52 bitb_47_52 bitb_47_53 R_bl
Cb_47_52 bit_47_52 gnd C_bl
Cbb_47_52 bitb_47_52 gnd C_bl
Rb_47_53 bit_47_53 bit_47_54 R_bl
Rbb_47_53 bitb_47_53 bitb_47_54 R_bl
Cb_47_53 bit_47_53 gnd C_bl
Cbb_47_53 bitb_47_53 gnd C_bl
Rb_47_54 bit_47_54 bit_47_55 R_bl
Rbb_47_54 bitb_47_54 bitb_47_55 R_bl
Cb_47_54 bit_47_54 gnd C_bl
Cbb_47_54 bitb_47_54 gnd C_bl
Rb_47_55 bit_47_55 bit_47_56 R_bl
Rbb_47_55 bitb_47_55 bitb_47_56 R_bl
Cb_47_55 bit_47_55 gnd C_bl
Cbb_47_55 bitb_47_55 gnd C_bl
Rb_47_56 bit_47_56 bit_47_57 R_bl
Rbb_47_56 bitb_47_56 bitb_47_57 R_bl
Cb_47_56 bit_47_56 gnd C_bl
Cbb_47_56 bitb_47_56 gnd C_bl
Rb_47_57 bit_47_57 bit_47_58 R_bl
Rbb_47_57 bitb_47_57 bitb_47_58 R_bl
Cb_47_57 bit_47_57 gnd C_bl
Cbb_47_57 bitb_47_57 gnd C_bl
Rb_47_58 bit_47_58 bit_47_59 R_bl
Rbb_47_58 bitb_47_58 bitb_47_59 R_bl
Cb_47_58 bit_47_58 gnd C_bl
Cbb_47_58 bitb_47_58 gnd C_bl
Rb_47_59 bit_47_59 bit_47_60 R_bl
Rbb_47_59 bitb_47_59 bitb_47_60 R_bl
Cb_47_59 bit_47_59 gnd C_bl
Cbb_47_59 bitb_47_59 gnd C_bl
Rb_47_60 bit_47_60 bit_47_61 R_bl
Rbb_47_60 bitb_47_60 bitb_47_61 R_bl
Cb_47_60 bit_47_60 gnd C_bl
Cbb_47_60 bitb_47_60 gnd C_bl
Rb_47_61 bit_47_61 bit_47_62 R_bl
Rbb_47_61 bitb_47_61 bitb_47_62 R_bl
Cb_47_61 bit_47_61 gnd C_bl
Cbb_47_61 bitb_47_61 gnd C_bl
Rb_47_62 bit_47_62 bit_47_63 R_bl
Rbb_47_62 bitb_47_62 bitb_47_63 R_bl
Cb_47_62 bit_47_62 gnd C_bl
Cbb_47_62 bitb_47_62 gnd C_bl
Rb_47_63 bit_47_63 bit_47_64 R_bl
Rbb_47_63 bitb_47_63 bitb_47_64 R_bl
Cb_47_63 bit_47_63 gnd C_bl
Cbb_47_63 bitb_47_63 gnd C_bl
Rb_47_64 bit_47_64 bit_47_65 R_bl
Rbb_47_64 bitb_47_64 bitb_47_65 R_bl
Cb_47_64 bit_47_64 gnd C_bl
Cbb_47_64 bitb_47_64 gnd C_bl
Rb_47_65 bit_47_65 bit_47_66 R_bl
Rbb_47_65 bitb_47_65 bitb_47_66 R_bl
Cb_47_65 bit_47_65 gnd C_bl
Cbb_47_65 bitb_47_65 gnd C_bl
Rb_47_66 bit_47_66 bit_47_67 R_bl
Rbb_47_66 bitb_47_66 bitb_47_67 R_bl
Cb_47_66 bit_47_66 gnd C_bl
Cbb_47_66 bitb_47_66 gnd C_bl
Rb_47_67 bit_47_67 bit_47_68 R_bl
Rbb_47_67 bitb_47_67 bitb_47_68 R_bl
Cb_47_67 bit_47_67 gnd C_bl
Cbb_47_67 bitb_47_67 gnd C_bl
Rb_47_68 bit_47_68 bit_47_69 R_bl
Rbb_47_68 bitb_47_68 bitb_47_69 R_bl
Cb_47_68 bit_47_68 gnd C_bl
Cbb_47_68 bitb_47_68 gnd C_bl
Rb_47_69 bit_47_69 bit_47_70 R_bl
Rbb_47_69 bitb_47_69 bitb_47_70 R_bl
Cb_47_69 bit_47_69 gnd C_bl
Cbb_47_69 bitb_47_69 gnd C_bl
Rb_47_70 bit_47_70 bit_47_71 R_bl
Rbb_47_70 bitb_47_70 bitb_47_71 R_bl
Cb_47_70 bit_47_70 gnd C_bl
Cbb_47_70 bitb_47_70 gnd C_bl
Rb_47_71 bit_47_71 bit_47_72 R_bl
Rbb_47_71 bitb_47_71 bitb_47_72 R_bl
Cb_47_71 bit_47_71 gnd C_bl
Cbb_47_71 bitb_47_71 gnd C_bl
Rb_47_72 bit_47_72 bit_47_73 R_bl
Rbb_47_72 bitb_47_72 bitb_47_73 R_bl
Cb_47_72 bit_47_72 gnd C_bl
Cbb_47_72 bitb_47_72 gnd C_bl
Rb_47_73 bit_47_73 bit_47_74 R_bl
Rbb_47_73 bitb_47_73 bitb_47_74 R_bl
Cb_47_73 bit_47_73 gnd C_bl
Cbb_47_73 bitb_47_73 gnd C_bl
Rb_47_74 bit_47_74 bit_47_75 R_bl
Rbb_47_74 bitb_47_74 bitb_47_75 R_bl
Cb_47_74 bit_47_74 gnd C_bl
Cbb_47_74 bitb_47_74 gnd C_bl
Rb_47_75 bit_47_75 bit_47_76 R_bl
Rbb_47_75 bitb_47_75 bitb_47_76 R_bl
Cb_47_75 bit_47_75 gnd C_bl
Cbb_47_75 bitb_47_75 gnd C_bl
Rb_47_76 bit_47_76 bit_47_77 R_bl
Rbb_47_76 bitb_47_76 bitb_47_77 R_bl
Cb_47_76 bit_47_76 gnd C_bl
Cbb_47_76 bitb_47_76 gnd C_bl
Rb_47_77 bit_47_77 bit_47_78 R_bl
Rbb_47_77 bitb_47_77 bitb_47_78 R_bl
Cb_47_77 bit_47_77 gnd C_bl
Cbb_47_77 bitb_47_77 gnd C_bl
Rb_47_78 bit_47_78 bit_47_79 R_bl
Rbb_47_78 bitb_47_78 bitb_47_79 R_bl
Cb_47_78 bit_47_78 gnd C_bl
Cbb_47_78 bitb_47_78 gnd C_bl
Rb_47_79 bit_47_79 bit_47_80 R_bl
Rbb_47_79 bitb_47_79 bitb_47_80 R_bl
Cb_47_79 bit_47_79 gnd C_bl
Cbb_47_79 bitb_47_79 gnd C_bl
Rb_47_80 bit_47_80 bit_47_81 R_bl
Rbb_47_80 bitb_47_80 bitb_47_81 R_bl
Cb_47_80 bit_47_80 gnd C_bl
Cbb_47_80 bitb_47_80 gnd C_bl
Rb_47_81 bit_47_81 bit_47_82 R_bl
Rbb_47_81 bitb_47_81 bitb_47_82 R_bl
Cb_47_81 bit_47_81 gnd C_bl
Cbb_47_81 bitb_47_81 gnd C_bl
Rb_47_82 bit_47_82 bit_47_83 R_bl
Rbb_47_82 bitb_47_82 bitb_47_83 R_bl
Cb_47_82 bit_47_82 gnd C_bl
Cbb_47_82 bitb_47_82 gnd C_bl
Rb_47_83 bit_47_83 bit_47_84 R_bl
Rbb_47_83 bitb_47_83 bitb_47_84 R_bl
Cb_47_83 bit_47_83 gnd C_bl
Cbb_47_83 bitb_47_83 gnd C_bl
Rb_47_84 bit_47_84 bit_47_85 R_bl
Rbb_47_84 bitb_47_84 bitb_47_85 R_bl
Cb_47_84 bit_47_84 gnd C_bl
Cbb_47_84 bitb_47_84 gnd C_bl
Rb_47_85 bit_47_85 bit_47_86 R_bl
Rbb_47_85 bitb_47_85 bitb_47_86 R_bl
Cb_47_85 bit_47_85 gnd C_bl
Cbb_47_85 bitb_47_85 gnd C_bl
Rb_47_86 bit_47_86 bit_47_87 R_bl
Rbb_47_86 bitb_47_86 bitb_47_87 R_bl
Cb_47_86 bit_47_86 gnd C_bl
Cbb_47_86 bitb_47_86 gnd C_bl
Rb_47_87 bit_47_87 bit_47_88 R_bl
Rbb_47_87 bitb_47_87 bitb_47_88 R_bl
Cb_47_87 bit_47_87 gnd C_bl
Cbb_47_87 bitb_47_87 gnd C_bl
Rb_47_88 bit_47_88 bit_47_89 R_bl
Rbb_47_88 bitb_47_88 bitb_47_89 R_bl
Cb_47_88 bit_47_88 gnd C_bl
Cbb_47_88 bitb_47_88 gnd C_bl
Rb_47_89 bit_47_89 bit_47_90 R_bl
Rbb_47_89 bitb_47_89 bitb_47_90 R_bl
Cb_47_89 bit_47_89 gnd C_bl
Cbb_47_89 bitb_47_89 gnd C_bl
Rb_47_90 bit_47_90 bit_47_91 R_bl
Rbb_47_90 bitb_47_90 bitb_47_91 R_bl
Cb_47_90 bit_47_90 gnd C_bl
Cbb_47_90 bitb_47_90 gnd C_bl
Rb_47_91 bit_47_91 bit_47_92 R_bl
Rbb_47_91 bitb_47_91 bitb_47_92 R_bl
Cb_47_91 bit_47_91 gnd C_bl
Cbb_47_91 bitb_47_91 gnd C_bl
Rb_47_92 bit_47_92 bit_47_93 R_bl
Rbb_47_92 bitb_47_92 bitb_47_93 R_bl
Cb_47_92 bit_47_92 gnd C_bl
Cbb_47_92 bitb_47_92 gnd C_bl
Rb_47_93 bit_47_93 bit_47_94 R_bl
Rbb_47_93 bitb_47_93 bitb_47_94 R_bl
Cb_47_93 bit_47_93 gnd C_bl
Cbb_47_93 bitb_47_93 gnd C_bl
Rb_47_94 bit_47_94 bit_47_95 R_bl
Rbb_47_94 bitb_47_94 bitb_47_95 R_bl
Cb_47_94 bit_47_94 gnd C_bl
Cbb_47_94 bitb_47_94 gnd C_bl
Rb_47_95 bit_47_95 bit_47_96 R_bl
Rbb_47_95 bitb_47_95 bitb_47_96 R_bl
Cb_47_95 bit_47_95 gnd C_bl
Cbb_47_95 bitb_47_95 gnd C_bl
Rb_47_96 bit_47_96 bit_47_97 R_bl
Rbb_47_96 bitb_47_96 bitb_47_97 R_bl
Cb_47_96 bit_47_96 gnd C_bl
Cbb_47_96 bitb_47_96 gnd C_bl
Rb_47_97 bit_47_97 bit_47_98 R_bl
Rbb_47_97 bitb_47_97 bitb_47_98 R_bl
Cb_47_97 bit_47_97 gnd C_bl
Cbb_47_97 bitb_47_97 gnd C_bl
Rb_47_98 bit_47_98 bit_47_99 R_bl
Rbb_47_98 bitb_47_98 bitb_47_99 R_bl
Cb_47_98 bit_47_98 gnd C_bl
Cbb_47_98 bitb_47_98 gnd C_bl
Rb_47_99 bit_47_99 bit_47_100 R_bl
Rbb_47_99 bitb_47_99 bitb_47_100 R_bl
Cb_47_99 bit_47_99 gnd C_bl
Cbb_47_99 bitb_47_99 gnd C_bl
Rb_48_0 bit_48_0 bit_48_1 R_bl
Rbb_48_0 bitb_48_0 bitb_48_1 R_bl
Cb_48_0 bit_48_0 gnd C_bl
Cbb_48_0 bitb_48_0 gnd C_bl
Rb_48_1 bit_48_1 bit_48_2 R_bl
Rbb_48_1 bitb_48_1 bitb_48_2 R_bl
Cb_48_1 bit_48_1 gnd C_bl
Cbb_48_1 bitb_48_1 gnd C_bl
Rb_48_2 bit_48_2 bit_48_3 R_bl
Rbb_48_2 bitb_48_2 bitb_48_3 R_bl
Cb_48_2 bit_48_2 gnd C_bl
Cbb_48_2 bitb_48_2 gnd C_bl
Rb_48_3 bit_48_3 bit_48_4 R_bl
Rbb_48_3 bitb_48_3 bitb_48_4 R_bl
Cb_48_3 bit_48_3 gnd C_bl
Cbb_48_3 bitb_48_3 gnd C_bl
Rb_48_4 bit_48_4 bit_48_5 R_bl
Rbb_48_4 bitb_48_4 bitb_48_5 R_bl
Cb_48_4 bit_48_4 gnd C_bl
Cbb_48_4 bitb_48_4 gnd C_bl
Rb_48_5 bit_48_5 bit_48_6 R_bl
Rbb_48_5 bitb_48_5 bitb_48_6 R_bl
Cb_48_5 bit_48_5 gnd C_bl
Cbb_48_5 bitb_48_5 gnd C_bl
Rb_48_6 bit_48_6 bit_48_7 R_bl
Rbb_48_6 bitb_48_6 bitb_48_7 R_bl
Cb_48_6 bit_48_6 gnd C_bl
Cbb_48_6 bitb_48_6 gnd C_bl
Rb_48_7 bit_48_7 bit_48_8 R_bl
Rbb_48_7 bitb_48_7 bitb_48_8 R_bl
Cb_48_7 bit_48_7 gnd C_bl
Cbb_48_7 bitb_48_7 gnd C_bl
Rb_48_8 bit_48_8 bit_48_9 R_bl
Rbb_48_8 bitb_48_8 bitb_48_9 R_bl
Cb_48_8 bit_48_8 gnd C_bl
Cbb_48_8 bitb_48_8 gnd C_bl
Rb_48_9 bit_48_9 bit_48_10 R_bl
Rbb_48_9 bitb_48_9 bitb_48_10 R_bl
Cb_48_9 bit_48_9 gnd C_bl
Cbb_48_9 bitb_48_9 gnd C_bl
Rb_48_10 bit_48_10 bit_48_11 R_bl
Rbb_48_10 bitb_48_10 bitb_48_11 R_bl
Cb_48_10 bit_48_10 gnd C_bl
Cbb_48_10 bitb_48_10 gnd C_bl
Rb_48_11 bit_48_11 bit_48_12 R_bl
Rbb_48_11 bitb_48_11 bitb_48_12 R_bl
Cb_48_11 bit_48_11 gnd C_bl
Cbb_48_11 bitb_48_11 gnd C_bl
Rb_48_12 bit_48_12 bit_48_13 R_bl
Rbb_48_12 bitb_48_12 bitb_48_13 R_bl
Cb_48_12 bit_48_12 gnd C_bl
Cbb_48_12 bitb_48_12 gnd C_bl
Rb_48_13 bit_48_13 bit_48_14 R_bl
Rbb_48_13 bitb_48_13 bitb_48_14 R_bl
Cb_48_13 bit_48_13 gnd C_bl
Cbb_48_13 bitb_48_13 gnd C_bl
Rb_48_14 bit_48_14 bit_48_15 R_bl
Rbb_48_14 bitb_48_14 bitb_48_15 R_bl
Cb_48_14 bit_48_14 gnd C_bl
Cbb_48_14 bitb_48_14 gnd C_bl
Rb_48_15 bit_48_15 bit_48_16 R_bl
Rbb_48_15 bitb_48_15 bitb_48_16 R_bl
Cb_48_15 bit_48_15 gnd C_bl
Cbb_48_15 bitb_48_15 gnd C_bl
Rb_48_16 bit_48_16 bit_48_17 R_bl
Rbb_48_16 bitb_48_16 bitb_48_17 R_bl
Cb_48_16 bit_48_16 gnd C_bl
Cbb_48_16 bitb_48_16 gnd C_bl
Rb_48_17 bit_48_17 bit_48_18 R_bl
Rbb_48_17 bitb_48_17 bitb_48_18 R_bl
Cb_48_17 bit_48_17 gnd C_bl
Cbb_48_17 bitb_48_17 gnd C_bl
Rb_48_18 bit_48_18 bit_48_19 R_bl
Rbb_48_18 bitb_48_18 bitb_48_19 R_bl
Cb_48_18 bit_48_18 gnd C_bl
Cbb_48_18 bitb_48_18 gnd C_bl
Rb_48_19 bit_48_19 bit_48_20 R_bl
Rbb_48_19 bitb_48_19 bitb_48_20 R_bl
Cb_48_19 bit_48_19 gnd C_bl
Cbb_48_19 bitb_48_19 gnd C_bl
Rb_48_20 bit_48_20 bit_48_21 R_bl
Rbb_48_20 bitb_48_20 bitb_48_21 R_bl
Cb_48_20 bit_48_20 gnd C_bl
Cbb_48_20 bitb_48_20 gnd C_bl
Rb_48_21 bit_48_21 bit_48_22 R_bl
Rbb_48_21 bitb_48_21 bitb_48_22 R_bl
Cb_48_21 bit_48_21 gnd C_bl
Cbb_48_21 bitb_48_21 gnd C_bl
Rb_48_22 bit_48_22 bit_48_23 R_bl
Rbb_48_22 bitb_48_22 bitb_48_23 R_bl
Cb_48_22 bit_48_22 gnd C_bl
Cbb_48_22 bitb_48_22 gnd C_bl
Rb_48_23 bit_48_23 bit_48_24 R_bl
Rbb_48_23 bitb_48_23 bitb_48_24 R_bl
Cb_48_23 bit_48_23 gnd C_bl
Cbb_48_23 bitb_48_23 gnd C_bl
Rb_48_24 bit_48_24 bit_48_25 R_bl
Rbb_48_24 bitb_48_24 bitb_48_25 R_bl
Cb_48_24 bit_48_24 gnd C_bl
Cbb_48_24 bitb_48_24 gnd C_bl
Rb_48_25 bit_48_25 bit_48_26 R_bl
Rbb_48_25 bitb_48_25 bitb_48_26 R_bl
Cb_48_25 bit_48_25 gnd C_bl
Cbb_48_25 bitb_48_25 gnd C_bl
Rb_48_26 bit_48_26 bit_48_27 R_bl
Rbb_48_26 bitb_48_26 bitb_48_27 R_bl
Cb_48_26 bit_48_26 gnd C_bl
Cbb_48_26 bitb_48_26 gnd C_bl
Rb_48_27 bit_48_27 bit_48_28 R_bl
Rbb_48_27 bitb_48_27 bitb_48_28 R_bl
Cb_48_27 bit_48_27 gnd C_bl
Cbb_48_27 bitb_48_27 gnd C_bl
Rb_48_28 bit_48_28 bit_48_29 R_bl
Rbb_48_28 bitb_48_28 bitb_48_29 R_bl
Cb_48_28 bit_48_28 gnd C_bl
Cbb_48_28 bitb_48_28 gnd C_bl
Rb_48_29 bit_48_29 bit_48_30 R_bl
Rbb_48_29 bitb_48_29 bitb_48_30 R_bl
Cb_48_29 bit_48_29 gnd C_bl
Cbb_48_29 bitb_48_29 gnd C_bl
Rb_48_30 bit_48_30 bit_48_31 R_bl
Rbb_48_30 bitb_48_30 bitb_48_31 R_bl
Cb_48_30 bit_48_30 gnd C_bl
Cbb_48_30 bitb_48_30 gnd C_bl
Rb_48_31 bit_48_31 bit_48_32 R_bl
Rbb_48_31 bitb_48_31 bitb_48_32 R_bl
Cb_48_31 bit_48_31 gnd C_bl
Cbb_48_31 bitb_48_31 gnd C_bl
Rb_48_32 bit_48_32 bit_48_33 R_bl
Rbb_48_32 bitb_48_32 bitb_48_33 R_bl
Cb_48_32 bit_48_32 gnd C_bl
Cbb_48_32 bitb_48_32 gnd C_bl
Rb_48_33 bit_48_33 bit_48_34 R_bl
Rbb_48_33 bitb_48_33 bitb_48_34 R_bl
Cb_48_33 bit_48_33 gnd C_bl
Cbb_48_33 bitb_48_33 gnd C_bl
Rb_48_34 bit_48_34 bit_48_35 R_bl
Rbb_48_34 bitb_48_34 bitb_48_35 R_bl
Cb_48_34 bit_48_34 gnd C_bl
Cbb_48_34 bitb_48_34 gnd C_bl
Rb_48_35 bit_48_35 bit_48_36 R_bl
Rbb_48_35 bitb_48_35 bitb_48_36 R_bl
Cb_48_35 bit_48_35 gnd C_bl
Cbb_48_35 bitb_48_35 gnd C_bl
Rb_48_36 bit_48_36 bit_48_37 R_bl
Rbb_48_36 bitb_48_36 bitb_48_37 R_bl
Cb_48_36 bit_48_36 gnd C_bl
Cbb_48_36 bitb_48_36 gnd C_bl
Rb_48_37 bit_48_37 bit_48_38 R_bl
Rbb_48_37 bitb_48_37 bitb_48_38 R_bl
Cb_48_37 bit_48_37 gnd C_bl
Cbb_48_37 bitb_48_37 gnd C_bl
Rb_48_38 bit_48_38 bit_48_39 R_bl
Rbb_48_38 bitb_48_38 bitb_48_39 R_bl
Cb_48_38 bit_48_38 gnd C_bl
Cbb_48_38 bitb_48_38 gnd C_bl
Rb_48_39 bit_48_39 bit_48_40 R_bl
Rbb_48_39 bitb_48_39 bitb_48_40 R_bl
Cb_48_39 bit_48_39 gnd C_bl
Cbb_48_39 bitb_48_39 gnd C_bl
Rb_48_40 bit_48_40 bit_48_41 R_bl
Rbb_48_40 bitb_48_40 bitb_48_41 R_bl
Cb_48_40 bit_48_40 gnd C_bl
Cbb_48_40 bitb_48_40 gnd C_bl
Rb_48_41 bit_48_41 bit_48_42 R_bl
Rbb_48_41 bitb_48_41 bitb_48_42 R_bl
Cb_48_41 bit_48_41 gnd C_bl
Cbb_48_41 bitb_48_41 gnd C_bl
Rb_48_42 bit_48_42 bit_48_43 R_bl
Rbb_48_42 bitb_48_42 bitb_48_43 R_bl
Cb_48_42 bit_48_42 gnd C_bl
Cbb_48_42 bitb_48_42 gnd C_bl
Rb_48_43 bit_48_43 bit_48_44 R_bl
Rbb_48_43 bitb_48_43 bitb_48_44 R_bl
Cb_48_43 bit_48_43 gnd C_bl
Cbb_48_43 bitb_48_43 gnd C_bl
Rb_48_44 bit_48_44 bit_48_45 R_bl
Rbb_48_44 bitb_48_44 bitb_48_45 R_bl
Cb_48_44 bit_48_44 gnd C_bl
Cbb_48_44 bitb_48_44 gnd C_bl
Rb_48_45 bit_48_45 bit_48_46 R_bl
Rbb_48_45 bitb_48_45 bitb_48_46 R_bl
Cb_48_45 bit_48_45 gnd C_bl
Cbb_48_45 bitb_48_45 gnd C_bl
Rb_48_46 bit_48_46 bit_48_47 R_bl
Rbb_48_46 bitb_48_46 bitb_48_47 R_bl
Cb_48_46 bit_48_46 gnd C_bl
Cbb_48_46 bitb_48_46 gnd C_bl
Rb_48_47 bit_48_47 bit_48_48 R_bl
Rbb_48_47 bitb_48_47 bitb_48_48 R_bl
Cb_48_47 bit_48_47 gnd C_bl
Cbb_48_47 bitb_48_47 gnd C_bl
Rb_48_48 bit_48_48 bit_48_49 R_bl
Rbb_48_48 bitb_48_48 bitb_48_49 R_bl
Cb_48_48 bit_48_48 gnd C_bl
Cbb_48_48 bitb_48_48 gnd C_bl
Rb_48_49 bit_48_49 bit_48_50 R_bl
Rbb_48_49 bitb_48_49 bitb_48_50 R_bl
Cb_48_49 bit_48_49 gnd C_bl
Cbb_48_49 bitb_48_49 gnd C_bl
Rb_48_50 bit_48_50 bit_48_51 R_bl
Rbb_48_50 bitb_48_50 bitb_48_51 R_bl
Cb_48_50 bit_48_50 gnd C_bl
Cbb_48_50 bitb_48_50 gnd C_bl
Rb_48_51 bit_48_51 bit_48_52 R_bl
Rbb_48_51 bitb_48_51 bitb_48_52 R_bl
Cb_48_51 bit_48_51 gnd C_bl
Cbb_48_51 bitb_48_51 gnd C_bl
Rb_48_52 bit_48_52 bit_48_53 R_bl
Rbb_48_52 bitb_48_52 bitb_48_53 R_bl
Cb_48_52 bit_48_52 gnd C_bl
Cbb_48_52 bitb_48_52 gnd C_bl
Rb_48_53 bit_48_53 bit_48_54 R_bl
Rbb_48_53 bitb_48_53 bitb_48_54 R_bl
Cb_48_53 bit_48_53 gnd C_bl
Cbb_48_53 bitb_48_53 gnd C_bl
Rb_48_54 bit_48_54 bit_48_55 R_bl
Rbb_48_54 bitb_48_54 bitb_48_55 R_bl
Cb_48_54 bit_48_54 gnd C_bl
Cbb_48_54 bitb_48_54 gnd C_bl
Rb_48_55 bit_48_55 bit_48_56 R_bl
Rbb_48_55 bitb_48_55 bitb_48_56 R_bl
Cb_48_55 bit_48_55 gnd C_bl
Cbb_48_55 bitb_48_55 gnd C_bl
Rb_48_56 bit_48_56 bit_48_57 R_bl
Rbb_48_56 bitb_48_56 bitb_48_57 R_bl
Cb_48_56 bit_48_56 gnd C_bl
Cbb_48_56 bitb_48_56 gnd C_bl
Rb_48_57 bit_48_57 bit_48_58 R_bl
Rbb_48_57 bitb_48_57 bitb_48_58 R_bl
Cb_48_57 bit_48_57 gnd C_bl
Cbb_48_57 bitb_48_57 gnd C_bl
Rb_48_58 bit_48_58 bit_48_59 R_bl
Rbb_48_58 bitb_48_58 bitb_48_59 R_bl
Cb_48_58 bit_48_58 gnd C_bl
Cbb_48_58 bitb_48_58 gnd C_bl
Rb_48_59 bit_48_59 bit_48_60 R_bl
Rbb_48_59 bitb_48_59 bitb_48_60 R_bl
Cb_48_59 bit_48_59 gnd C_bl
Cbb_48_59 bitb_48_59 gnd C_bl
Rb_48_60 bit_48_60 bit_48_61 R_bl
Rbb_48_60 bitb_48_60 bitb_48_61 R_bl
Cb_48_60 bit_48_60 gnd C_bl
Cbb_48_60 bitb_48_60 gnd C_bl
Rb_48_61 bit_48_61 bit_48_62 R_bl
Rbb_48_61 bitb_48_61 bitb_48_62 R_bl
Cb_48_61 bit_48_61 gnd C_bl
Cbb_48_61 bitb_48_61 gnd C_bl
Rb_48_62 bit_48_62 bit_48_63 R_bl
Rbb_48_62 bitb_48_62 bitb_48_63 R_bl
Cb_48_62 bit_48_62 gnd C_bl
Cbb_48_62 bitb_48_62 gnd C_bl
Rb_48_63 bit_48_63 bit_48_64 R_bl
Rbb_48_63 bitb_48_63 bitb_48_64 R_bl
Cb_48_63 bit_48_63 gnd C_bl
Cbb_48_63 bitb_48_63 gnd C_bl
Rb_48_64 bit_48_64 bit_48_65 R_bl
Rbb_48_64 bitb_48_64 bitb_48_65 R_bl
Cb_48_64 bit_48_64 gnd C_bl
Cbb_48_64 bitb_48_64 gnd C_bl
Rb_48_65 bit_48_65 bit_48_66 R_bl
Rbb_48_65 bitb_48_65 bitb_48_66 R_bl
Cb_48_65 bit_48_65 gnd C_bl
Cbb_48_65 bitb_48_65 gnd C_bl
Rb_48_66 bit_48_66 bit_48_67 R_bl
Rbb_48_66 bitb_48_66 bitb_48_67 R_bl
Cb_48_66 bit_48_66 gnd C_bl
Cbb_48_66 bitb_48_66 gnd C_bl
Rb_48_67 bit_48_67 bit_48_68 R_bl
Rbb_48_67 bitb_48_67 bitb_48_68 R_bl
Cb_48_67 bit_48_67 gnd C_bl
Cbb_48_67 bitb_48_67 gnd C_bl
Rb_48_68 bit_48_68 bit_48_69 R_bl
Rbb_48_68 bitb_48_68 bitb_48_69 R_bl
Cb_48_68 bit_48_68 gnd C_bl
Cbb_48_68 bitb_48_68 gnd C_bl
Rb_48_69 bit_48_69 bit_48_70 R_bl
Rbb_48_69 bitb_48_69 bitb_48_70 R_bl
Cb_48_69 bit_48_69 gnd C_bl
Cbb_48_69 bitb_48_69 gnd C_bl
Rb_48_70 bit_48_70 bit_48_71 R_bl
Rbb_48_70 bitb_48_70 bitb_48_71 R_bl
Cb_48_70 bit_48_70 gnd C_bl
Cbb_48_70 bitb_48_70 gnd C_bl
Rb_48_71 bit_48_71 bit_48_72 R_bl
Rbb_48_71 bitb_48_71 bitb_48_72 R_bl
Cb_48_71 bit_48_71 gnd C_bl
Cbb_48_71 bitb_48_71 gnd C_bl
Rb_48_72 bit_48_72 bit_48_73 R_bl
Rbb_48_72 bitb_48_72 bitb_48_73 R_bl
Cb_48_72 bit_48_72 gnd C_bl
Cbb_48_72 bitb_48_72 gnd C_bl
Rb_48_73 bit_48_73 bit_48_74 R_bl
Rbb_48_73 bitb_48_73 bitb_48_74 R_bl
Cb_48_73 bit_48_73 gnd C_bl
Cbb_48_73 bitb_48_73 gnd C_bl
Rb_48_74 bit_48_74 bit_48_75 R_bl
Rbb_48_74 bitb_48_74 bitb_48_75 R_bl
Cb_48_74 bit_48_74 gnd C_bl
Cbb_48_74 bitb_48_74 gnd C_bl
Rb_48_75 bit_48_75 bit_48_76 R_bl
Rbb_48_75 bitb_48_75 bitb_48_76 R_bl
Cb_48_75 bit_48_75 gnd C_bl
Cbb_48_75 bitb_48_75 gnd C_bl
Rb_48_76 bit_48_76 bit_48_77 R_bl
Rbb_48_76 bitb_48_76 bitb_48_77 R_bl
Cb_48_76 bit_48_76 gnd C_bl
Cbb_48_76 bitb_48_76 gnd C_bl
Rb_48_77 bit_48_77 bit_48_78 R_bl
Rbb_48_77 bitb_48_77 bitb_48_78 R_bl
Cb_48_77 bit_48_77 gnd C_bl
Cbb_48_77 bitb_48_77 gnd C_bl
Rb_48_78 bit_48_78 bit_48_79 R_bl
Rbb_48_78 bitb_48_78 bitb_48_79 R_bl
Cb_48_78 bit_48_78 gnd C_bl
Cbb_48_78 bitb_48_78 gnd C_bl
Rb_48_79 bit_48_79 bit_48_80 R_bl
Rbb_48_79 bitb_48_79 bitb_48_80 R_bl
Cb_48_79 bit_48_79 gnd C_bl
Cbb_48_79 bitb_48_79 gnd C_bl
Rb_48_80 bit_48_80 bit_48_81 R_bl
Rbb_48_80 bitb_48_80 bitb_48_81 R_bl
Cb_48_80 bit_48_80 gnd C_bl
Cbb_48_80 bitb_48_80 gnd C_bl
Rb_48_81 bit_48_81 bit_48_82 R_bl
Rbb_48_81 bitb_48_81 bitb_48_82 R_bl
Cb_48_81 bit_48_81 gnd C_bl
Cbb_48_81 bitb_48_81 gnd C_bl
Rb_48_82 bit_48_82 bit_48_83 R_bl
Rbb_48_82 bitb_48_82 bitb_48_83 R_bl
Cb_48_82 bit_48_82 gnd C_bl
Cbb_48_82 bitb_48_82 gnd C_bl
Rb_48_83 bit_48_83 bit_48_84 R_bl
Rbb_48_83 bitb_48_83 bitb_48_84 R_bl
Cb_48_83 bit_48_83 gnd C_bl
Cbb_48_83 bitb_48_83 gnd C_bl
Rb_48_84 bit_48_84 bit_48_85 R_bl
Rbb_48_84 bitb_48_84 bitb_48_85 R_bl
Cb_48_84 bit_48_84 gnd C_bl
Cbb_48_84 bitb_48_84 gnd C_bl
Rb_48_85 bit_48_85 bit_48_86 R_bl
Rbb_48_85 bitb_48_85 bitb_48_86 R_bl
Cb_48_85 bit_48_85 gnd C_bl
Cbb_48_85 bitb_48_85 gnd C_bl
Rb_48_86 bit_48_86 bit_48_87 R_bl
Rbb_48_86 bitb_48_86 bitb_48_87 R_bl
Cb_48_86 bit_48_86 gnd C_bl
Cbb_48_86 bitb_48_86 gnd C_bl
Rb_48_87 bit_48_87 bit_48_88 R_bl
Rbb_48_87 bitb_48_87 bitb_48_88 R_bl
Cb_48_87 bit_48_87 gnd C_bl
Cbb_48_87 bitb_48_87 gnd C_bl
Rb_48_88 bit_48_88 bit_48_89 R_bl
Rbb_48_88 bitb_48_88 bitb_48_89 R_bl
Cb_48_88 bit_48_88 gnd C_bl
Cbb_48_88 bitb_48_88 gnd C_bl
Rb_48_89 bit_48_89 bit_48_90 R_bl
Rbb_48_89 bitb_48_89 bitb_48_90 R_bl
Cb_48_89 bit_48_89 gnd C_bl
Cbb_48_89 bitb_48_89 gnd C_bl
Rb_48_90 bit_48_90 bit_48_91 R_bl
Rbb_48_90 bitb_48_90 bitb_48_91 R_bl
Cb_48_90 bit_48_90 gnd C_bl
Cbb_48_90 bitb_48_90 gnd C_bl
Rb_48_91 bit_48_91 bit_48_92 R_bl
Rbb_48_91 bitb_48_91 bitb_48_92 R_bl
Cb_48_91 bit_48_91 gnd C_bl
Cbb_48_91 bitb_48_91 gnd C_bl
Rb_48_92 bit_48_92 bit_48_93 R_bl
Rbb_48_92 bitb_48_92 bitb_48_93 R_bl
Cb_48_92 bit_48_92 gnd C_bl
Cbb_48_92 bitb_48_92 gnd C_bl
Rb_48_93 bit_48_93 bit_48_94 R_bl
Rbb_48_93 bitb_48_93 bitb_48_94 R_bl
Cb_48_93 bit_48_93 gnd C_bl
Cbb_48_93 bitb_48_93 gnd C_bl
Rb_48_94 bit_48_94 bit_48_95 R_bl
Rbb_48_94 bitb_48_94 bitb_48_95 R_bl
Cb_48_94 bit_48_94 gnd C_bl
Cbb_48_94 bitb_48_94 gnd C_bl
Rb_48_95 bit_48_95 bit_48_96 R_bl
Rbb_48_95 bitb_48_95 bitb_48_96 R_bl
Cb_48_95 bit_48_95 gnd C_bl
Cbb_48_95 bitb_48_95 gnd C_bl
Rb_48_96 bit_48_96 bit_48_97 R_bl
Rbb_48_96 bitb_48_96 bitb_48_97 R_bl
Cb_48_96 bit_48_96 gnd C_bl
Cbb_48_96 bitb_48_96 gnd C_bl
Rb_48_97 bit_48_97 bit_48_98 R_bl
Rbb_48_97 bitb_48_97 bitb_48_98 R_bl
Cb_48_97 bit_48_97 gnd C_bl
Cbb_48_97 bitb_48_97 gnd C_bl
Rb_48_98 bit_48_98 bit_48_99 R_bl
Rbb_48_98 bitb_48_98 bitb_48_99 R_bl
Cb_48_98 bit_48_98 gnd C_bl
Cbb_48_98 bitb_48_98 gnd C_bl
Rb_48_99 bit_48_99 bit_48_100 R_bl
Rbb_48_99 bitb_48_99 bitb_48_100 R_bl
Cb_48_99 bit_48_99 gnd C_bl
Cbb_48_99 bitb_48_99 gnd C_bl
Rb_49_0 bit_49_0 bit_49_1 R_bl
Rbb_49_0 bitb_49_0 bitb_49_1 R_bl
Cb_49_0 bit_49_0 gnd C_bl
Cbb_49_0 bitb_49_0 gnd C_bl
Rb_49_1 bit_49_1 bit_49_2 R_bl
Rbb_49_1 bitb_49_1 bitb_49_2 R_bl
Cb_49_1 bit_49_1 gnd C_bl
Cbb_49_1 bitb_49_1 gnd C_bl
Rb_49_2 bit_49_2 bit_49_3 R_bl
Rbb_49_2 bitb_49_2 bitb_49_3 R_bl
Cb_49_2 bit_49_2 gnd C_bl
Cbb_49_2 bitb_49_2 gnd C_bl
Rb_49_3 bit_49_3 bit_49_4 R_bl
Rbb_49_3 bitb_49_3 bitb_49_4 R_bl
Cb_49_3 bit_49_3 gnd C_bl
Cbb_49_3 bitb_49_3 gnd C_bl
Rb_49_4 bit_49_4 bit_49_5 R_bl
Rbb_49_4 bitb_49_4 bitb_49_5 R_bl
Cb_49_4 bit_49_4 gnd C_bl
Cbb_49_4 bitb_49_4 gnd C_bl
Rb_49_5 bit_49_5 bit_49_6 R_bl
Rbb_49_5 bitb_49_5 bitb_49_6 R_bl
Cb_49_5 bit_49_5 gnd C_bl
Cbb_49_5 bitb_49_5 gnd C_bl
Rb_49_6 bit_49_6 bit_49_7 R_bl
Rbb_49_6 bitb_49_6 bitb_49_7 R_bl
Cb_49_6 bit_49_6 gnd C_bl
Cbb_49_6 bitb_49_6 gnd C_bl
Rb_49_7 bit_49_7 bit_49_8 R_bl
Rbb_49_7 bitb_49_7 bitb_49_8 R_bl
Cb_49_7 bit_49_7 gnd C_bl
Cbb_49_7 bitb_49_7 gnd C_bl
Rb_49_8 bit_49_8 bit_49_9 R_bl
Rbb_49_8 bitb_49_8 bitb_49_9 R_bl
Cb_49_8 bit_49_8 gnd C_bl
Cbb_49_8 bitb_49_8 gnd C_bl
Rb_49_9 bit_49_9 bit_49_10 R_bl
Rbb_49_9 bitb_49_9 bitb_49_10 R_bl
Cb_49_9 bit_49_9 gnd C_bl
Cbb_49_9 bitb_49_9 gnd C_bl
Rb_49_10 bit_49_10 bit_49_11 R_bl
Rbb_49_10 bitb_49_10 bitb_49_11 R_bl
Cb_49_10 bit_49_10 gnd C_bl
Cbb_49_10 bitb_49_10 gnd C_bl
Rb_49_11 bit_49_11 bit_49_12 R_bl
Rbb_49_11 bitb_49_11 bitb_49_12 R_bl
Cb_49_11 bit_49_11 gnd C_bl
Cbb_49_11 bitb_49_11 gnd C_bl
Rb_49_12 bit_49_12 bit_49_13 R_bl
Rbb_49_12 bitb_49_12 bitb_49_13 R_bl
Cb_49_12 bit_49_12 gnd C_bl
Cbb_49_12 bitb_49_12 gnd C_bl
Rb_49_13 bit_49_13 bit_49_14 R_bl
Rbb_49_13 bitb_49_13 bitb_49_14 R_bl
Cb_49_13 bit_49_13 gnd C_bl
Cbb_49_13 bitb_49_13 gnd C_bl
Rb_49_14 bit_49_14 bit_49_15 R_bl
Rbb_49_14 bitb_49_14 bitb_49_15 R_bl
Cb_49_14 bit_49_14 gnd C_bl
Cbb_49_14 bitb_49_14 gnd C_bl
Rb_49_15 bit_49_15 bit_49_16 R_bl
Rbb_49_15 bitb_49_15 bitb_49_16 R_bl
Cb_49_15 bit_49_15 gnd C_bl
Cbb_49_15 bitb_49_15 gnd C_bl
Rb_49_16 bit_49_16 bit_49_17 R_bl
Rbb_49_16 bitb_49_16 bitb_49_17 R_bl
Cb_49_16 bit_49_16 gnd C_bl
Cbb_49_16 bitb_49_16 gnd C_bl
Rb_49_17 bit_49_17 bit_49_18 R_bl
Rbb_49_17 bitb_49_17 bitb_49_18 R_bl
Cb_49_17 bit_49_17 gnd C_bl
Cbb_49_17 bitb_49_17 gnd C_bl
Rb_49_18 bit_49_18 bit_49_19 R_bl
Rbb_49_18 bitb_49_18 bitb_49_19 R_bl
Cb_49_18 bit_49_18 gnd C_bl
Cbb_49_18 bitb_49_18 gnd C_bl
Rb_49_19 bit_49_19 bit_49_20 R_bl
Rbb_49_19 bitb_49_19 bitb_49_20 R_bl
Cb_49_19 bit_49_19 gnd C_bl
Cbb_49_19 bitb_49_19 gnd C_bl
Rb_49_20 bit_49_20 bit_49_21 R_bl
Rbb_49_20 bitb_49_20 bitb_49_21 R_bl
Cb_49_20 bit_49_20 gnd C_bl
Cbb_49_20 bitb_49_20 gnd C_bl
Rb_49_21 bit_49_21 bit_49_22 R_bl
Rbb_49_21 bitb_49_21 bitb_49_22 R_bl
Cb_49_21 bit_49_21 gnd C_bl
Cbb_49_21 bitb_49_21 gnd C_bl
Rb_49_22 bit_49_22 bit_49_23 R_bl
Rbb_49_22 bitb_49_22 bitb_49_23 R_bl
Cb_49_22 bit_49_22 gnd C_bl
Cbb_49_22 bitb_49_22 gnd C_bl
Rb_49_23 bit_49_23 bit_49_24 R_bl
Rbb_49_23 bitb_49_23 bitb_49_24 R_bl
Cb_49_23 bit_49_23 gnd C_bl
Cbb_49_23 bitb_49_23 gnd C_bl
Rb_49_24 bit_49_24 bit_49_25 R_bl
Rbb_49_24 bitb_49_24 bitb_49_25 R_bl
Cb_49_24 bit_49_24 gnd C_bl
Cbb_49_24 bitb_49_24 gnd C_bl
Rb_49_25 bit_49_25 bit_49_26 R_bl
Rbb_49_25 bitb_49_25 bitb_49_26 R_bl
Cb_49_25 bit_49_25 gnd C_bl
Cbb_49_25 bitb_49_25 gnd C_bl
Rb_49_26 bit_49_26 bit_49_27 R_bl
Rbb_49_26 bitb_49_26 bitb_49_27 R_bl
Cb_49_26 bit_49_26 gnd C_bl
Cbb_49_26 bitb_49_26 gnd C_bl
Rb_49_27 bit_49_27 bit_49_28 R_bl
Rbb_49_27 bitb_49_27 bitb_49_28 R_bl
Cb_49_27 bit_49_27 gnd C_bl
Cbb_49_27 bitb_49_27 gnd C_bl
Rb_49_28 bit_49_28 bit_49_29 R_bl
Rbb_49_28 bitb_49_28 bitb_49_29 R_bl
Cb_49_28 bit_49_28 gnd C_bl
Cbb_49_28 bitb_49_28 gnd C_bl
Rb_49_29 bit_49_29 bit_49_30 R_bl
Rbb_49_29 bitb_49_29 bitb_49_30 R_bl
Cb_49_29 bit_49_29 gnd C_bl
Cbb_49_29 bitb_49_29 gnd C_bl
Rb_49_30 bit_49_30 bit_49_31 R_bl
Rbb_49_30 bitb_49_30 bitb_49_31 R_bl
Cb_49_30 bit_49_30 gnd C_bl
Cbb_49_30 bitb_49_30 gnd C_bl
Rb_49_31 bit_49_31 bit_49_32 R_bl
Rbb_49_31 bitb_49_31 bitb_49_32 R_bl
Cb_49_31 bit_49_31 gnd C_bl
Cbb_49_31 bitb_49_31 gnd C_bl
Rb_49_32 bit_49_32 bit_49_33 R_bl
Rbb_49_32 bitb_49_32 bitb_49_33 R_bl
Cb_49_32 bit_49_32 gnd C_bl
Cbb_49_32 bitb_49_32 gnd C_bl
Rb_49_33 bit_49_33 bit_49_34 R_bl
Rbb_49_33 bitb_49_33 bitb_49_34 R_bl
Cb_49_33 bit_49_33 gnd C_bl
Cbb_49_33 bitb_49_33 gnd C_bl
Rb_49_34 bit_49_34 bit_49_35 R_bl
Rbb_49_34 bitb_49_34 bitb_49_35 R_bl
Cb_49_34 bit_49_34 gnd C_bl
Cbb_49_34 bitb_49_34 gnd C_bl
Rb_49_35 bit_49_35 bit_49_36 R_bl
Rbb_49_35 bitb_49_35 bitb_49_36 R_bl
Cb_49_35 bit_49_35 gnd C_bl
Cbb_49_35 bitb_49_35 gnd C_bl
Rb_49_36 bit_49_36 bit_49_37 R_bl
Rbb_49_36 bitb_49_36 bitb_49_37 R_bl
Cb_49_36 bit_49_36 gnd C_bl
Cbb_49_36 bitb_49_36 gnd C_bl
Rb_49_37 bit_49_37 bit_49_38 R_bl
Rbb_49_37 bitb_49_37 bitb_49_38 R_bl
Cb_49_37 bit_49_37 gnd C_bl
Cbb_49_37 bitb_49_37 gnd C_bl
Rb_49_38 bit_49_38 bit_49_39 R_bl
Rbb_49_38 bitb_49_38 bitb_49_39 R_bl
Cb_49_38 bit_49_38 gnd C_bl
Cbb_49_38 bitb_49_38 gnd C_bl
Rb_49_39 bit_49_39 bit_49_40 R_bl
Rbb_49_39 bitb_49_39 bitb_49_40 R_bl
Cb_49_39 bit_49_39 gnd C_bl
Cbb_49_39 bitb_49_39 gnd C_bl
Rb_49_40 bit_49_40 bit_49_41 R_bl
Rbb_49_40 bitb_49_40 bitb_49_41 R_bl
Cb_49_40 bit_49_40 gnd C_bl
Cbb_49_40 bitb_49_40 gnd C_bl
Rb_49_41 bit_49_41 bit_49_42 R_bl
Rbb_49_41 bitb_49_41 bitb_49_42 R_bl
Cb_49_41 bit_49_41 gnd C_bl
Cbb_49_41 bitb_49_41 gnd C_bl
Rb_49_42 bit_49_42 bit_49_43 R_bl
Rbb_49_42 bitb_49_42 bitb_49_43 R_bl
Cb_49_42 bit_49_42 gnd C_bl
Cbb_49_42 bitb_49_42 gnd C_bl
Rb_49_43 bit_49_43 bit_49_44 R_bl
Rbb_49_43 bitb_49_43 bitb_49_44 R_bl
Cb_49_43 bit_49_43 gnd C_bl
Cbb_49_43 bitb_49_43 gnd C_bl
Rb_49_44 bit_49_44 bit_49_45 R_bl
Rbb_49_44 bitb_49_44 bitb_49_45 R_bl
Cb_49_44 bit_49_44 gnd C_bl
Cbb_49_44 bitb_49_44 gnd C_bl
Rb_49_45 bit_49_45 bit_49_46 R_bl
Rbb_49_45 bitb_49_45 bitb_49_46 R_bl
Cb_49_45 bit_49_45 gnd C_bl
Cbb_49_45 bitb_49_45 gnd C_bl
Rb_49_46 bit_49_46 bit_49_47 R_bl
Rbb_49_46 bitb_49_46 bitb_49_47 R_bl
Cb_49_46 bit_49_46 gnd C_bl
Cbb_49_46 bitb_49_46 gnd C_bl
Rb_49_47 bit_49_47 bit_49_48 R_bl
Rbb_49_47 bitb_49_47 bitb_49_48 R_bl
Cb_49_47 bit_49_47 gnd C_bl
Cbb_49_47 bitb_49_47 gnd C_bl
Rb_49_48 bit_49_48 bit_49_49 R_bl
Rbb_49_48 bitb_49_48 bitb_49_49 R_bl
Cb_49_48 bit_49_48 gnd C_bl
Cbb_49_48 bitb_49_48 gnd C_bl
Rb_49_49 bit_49_49 bit_49_50 R_bl
Rbb_49_49 bitb_49_49 bitb_49_50 R_bl
Cb_49_49 bit_49_49 gnd C_bl
Cbb_49_49 bitb_49_49 gnd C_bl
Rb_49_50 bit_49_50 bit_49_51 R_bl
Rbb_49_50 bitb_49_50 bitb_49_51 R_bl
Cb_49_50 bit_49_50 gnd C_bl
Cbb_49_50 bitb_49_50 gnd C_bl
Rb_49_51 bit_49_51 bit_49_52 R_bl
Rbb_49_51 bitb_49_51 bitb_49_52 R_bl
Cb_49_51 bit_49_51 gnd C_bl
Cbb_49_51 bitb_49_51 gnd C_bl
Rb_49_52 bit_49_52 bit_49_53 R_bl
Rbb_49_52 bitb_49_52 bitb_49_53 R_bl
Cb_49_52 bit_49_52 gnd C_bl
Cbb_49_52 bitb_49_52 gnd C_bl
Rb_49_53 bit_49_53 bit_49_54 R_bl
Rbb_49_53 bitb_49_53 bitb_49_54 R_bl
Cb_49_53 bit_49_53 gnd C_bl
Cbb_49_53 bitb_49_53 gnd C_bl
Rb_49_54 bit_49_54 bit_49_55 R_bl
Rbb_49_54 bitb_49_54 bitb_49_55 R_bl
Cb_49_54 bit_49_54 gnd C_bl
Cbb_49_54 bitb_49_54 gnd C_bl
Rb_49_55 bit_49_55 bit_49_56 R_bl
Rbb_49_55 bitb_49_55 bitb_49_56 R_bl
Cb_49_55 bit_49_55 gnd C_bl
Cbb_49_55 bitb_49_55 gnd C_bl
Rb_49_56 bit_49_56 bit_49_57 R_bl
Rbb_49_56 bitb_49_56 bitb_49_57 R_bl
Cb_49_56 bit_49_56 gnd C_bl
Cbb_49_56 bitb_49_56 gnd C_bl
Rb_49_57 bit_49_57 bit_49_58 R_bl
Rbb_49_57 bitb_49_57 bitb_49_58 R_bl
Cb_49_57 bit_49_57 gnd C_bl
Cbb_49_57 bitb_49_57 gnd C_bl
Rb_49_58 bit_49_58 bit_49_59 R_bl
Rbb_49_58 bitb_49_58 bitb_49_59 R_bl
Cb_49_58 bit_49_58 gnd C_bl
Cbb_49_58 bitb_49_58 gnd C_bl
Rb_49_59 bit_49_59 bit_49_60 R_bl
Rbb_49_59 bitb_49_59 bitb_49_60 R_bl
Cb_49_59 bit_49_59 gnd C_bl
Cbb_49_59 bitb_49_59 gnd C_bl
Rb_49_60 bit_49_60 bit_49_61 R_bl
Rbb_49_60 bitb_49_60 bitb_49_61 R_bl
Cb_49_60 bit_49_60 gnd C_bl
Cbb_49_60 bitb_49_60 gnd C_bl
Rb_49_61 bit_49_61 bit_49_62 R_bl
Rbb_49_61 bitb_49_61 bitb_49_62 R_bl
Cb_49_61 bit_49_61 gnd C_bl
Cbb_49_61 bitb_49_61 gnd C_bl
Rb_49_62 bit_49_62 bit_49_63 R_bl
Rbb_49_62 bitb_49_62 bitb_49_63 R_bl
Cb_49_62 bit_49_62 gnd C_bl
Cbb_49_62 bitb_49_62 gnd C_bl
Rb_49_63 bit_49_63 bit_49_64 R_bl
Rbb_49_63 bitb_49_63 bitb_49_64 R_bl
Cb_49_63 bit_49_63 gnd C_bl
Cbb_49_63 bitb_49_63 gnd C_bl
Rb_49_64 bit_49_64 bit_49_65 R_bl
Rbb_49_64 bitb_49_64 bitb_49_65 R_bl
Cb_49_64 bit_49_64 gnd C_bl
Cbb_49_64 bitb_49_64 gnd C_bl
Rb_49_65 bit_49_65 bit_49_66 R_bl
Rbb_49_65 bitb_49_65 bitb_49_66 R_bl
Cb_49_65 bit_49_65 gnd C_bl
Cbb_49_65 bitb_49_65 gnd C_bl
Rb_49_66 bit_49_66 bit_49_67 R_bl
Rbb_49_66 bitb_49_66 bitb_49_67 R_bl
Cb_49_66 bit_49_66 gnd C_bl
Cbb_49_66 bitb_49_66 gnd C_bl
Rb_49_67 bit_49_67 bit_49_68 R_bl
Rbb_49_67 bitb_49_67 bitb_49_68 R_bl
Cb_49_67 bit_49_67 gnd C_bl
Cbb_49_67 bitb_49_67 gnd C_bl
Rb_49_68 bit_49_68 bit_49_69 R_bl
Rbb_49_68 bitb_49_68 bitb_49_69 R_bl
Cb_49_68 bit_49_68 gnd C_bl
Cbb_49_68 bitb_49_68 gnd C_bl
Rb_49_69 bit_49_69 bit_49_70 R_bl
Rbb_49_69 bitb_49_69 bitb_49_70 R_bl
Cb_49_69 bit_49_69 gnd C_bl
Cbb_49_69 bitb_49_69 gnd C_bl
Rb_49_70 bit_49_70 bit_49_71 R_bl
Rbb_49_70 bitb_49_70 bitb_49_71 R_bl
Cb_49_70 bit_49_70 gnd C_bl
Cbb_49_70 bitb_49_70 gnd C_bl
Rb_49_71 bit_49_71 bit_49_72 R_bl
Rbb_49_71 bitb_49_71 bitb_49_72 R_bl
Cb_49_71 bit_49_71 gnd C_bl
Cbb_49_71 bitb_49_71 gnd C_bl
Rb_49_72 bit_49_72 bit_49_73 R_bl
Rbb_49_72 bitb_49_72 bitb_49_73 R_bl
Cb_49_72 bit_49_72 gnd C_bl
Cbb_49_72 bitb_49_72 gnd C_bl
Rb_49_73 bit_49_73 bit_49_74 R_bl
Rbb_49_73 bitb_49_73 bitb_49_74 R_bl
Cb_49_73 bit_49_73 gnd C_bl
Cbb_49_73 bitb_49_73 gnd C_bl
Rb_49_74 bit_49_74 bit_49_75 R_bl
Rbb_49_74 bitb_49_74 bitb_49_75 R_bl
Cb_49_74 bit_49_74 gnd C_bl
Cbb_49_74 bitb_49_74 gnd C_bl
Rb_49_75 bit_49_75 bit_49_76 R_bl
Rbb_49_75 bitb_49_75 bitb_49_76 R_bl
Cb_49_75 bit_49_75 gnd C_bl
Cbb_49_75 bitb_49_75 gnd C_bl
Rb_49_76 bit_49_76 bit_49_77 R_bl
Rbb_49_76 bitb_49_76 bitb_49_77 R_bl
Cb_49_76 bit_49_76 gnd C_bl
Cbb_49_76 bitb_49_76 gnd C_bl
Rb_49_77 bit_49_77 bit_49_78 R_bl
Rbb_49_77 bitb_49_77 bitb_49_78 R_bl
Cb_49_77 bit_49_77 gnd C_bl
Cbb_49_77 bitb_49_77 gnd C_bl
Rb_49_78 bit_49_78 bit_49_79 R_bl
Rbb_49_78 bitb_49_78 bitb_49_79 R_bl
Cb_49_78 bit_49_78 gnd C_bl
Cbb_49_78 bitb_49_78 gnd C_bl
Rb_49_79 bit_49_79 bit_49_80 R_bl
Rbb_49_79 bitb_49_79 bitb_49_80 R_bl
Cb_49_79 bit_49_79 gnd C_bl
Cbb_49_79 bitb_49_79 gnd C_bl
Rb_49_80 bit_49_80 bit_49_81 R_bl
Rbb_49_80 bitb_49_80 bitb_49_81 R_bl
Cb_49_80 bit_49_80 gnd C_bl
Cbb_49_80 bitb_49_80 gnd C_bl
Rb_49_81 bit_49_81 bit_49_82 R_bl
Rbb_49_81 bitb_49_81 bitb_49_82 R_bl
Cb_49_81 bit_49_81 gnd C_bl
Cbb_49_81 bitb_49_81 gnd C_bl
Rb_49_82 bit_49_82 bit_49_83 R_bl
Rbb_49_82 bitb_49_82 bitb_49_83 R_bl
Cb_49_82 bit_49_82 gnd C_bl
Cbb_49_82 bitb_49_82 gnd C_bl
Rb_49_83 bit_49_83 bit_49_84 R_bl
Rbb_49_83 bitb_49_83 bitb_49_84 R_bl
Cb_49_83 bit_49_83 gnd C_bl
Cbb_49_83 bitb_49_83 gnd C_bl
Rb_49_84 bit_49_84 bit_49_85 R_bl
Rbb_49_84 bitb_49_84 bitb_49_85 R_bl
Cb_49_84 bit_49_84 gnd C_bl
Cbb_49_84 bitb_49_84 gnd C_bl
Rb_49_85 bit_49_85 bit_49_86 R_bl
Rbb_49_85 bitb_49_85 bitb_49_86 R_bl
Cb_49_85 bit_49_85 gnd C_bl
Cbb_49_85 bitb_49_85 gnd C_bl
Rb_49_86 bit_49_86 bit_49_87 R_bl
Rbb_49_86 bitb_49_86 bitb_49_87 R_bl
Cb_49_86 bit_49_86 gnd C_bl
Cbb_49_86 bitb_49_86 gnd C_bl
Rb_49_87 bit_49_87 bit_49_88 R_bl
Rbb_49_87 bitb_49_87 bitb_49_88 R_bl
Cb_49_87 bit_49_87 gnd C_bl
Cbb_49_87 bitb_49_87 gnd C_bl
Rb_49_88 bit_49_88 bit_49_89 R_bl
Rbb_49_88 bitb_49_88 bitb_49_89 R_bl
Cb_49_88 bit_49_88 gnd C_bl
Cbb_49_88 bitb_49_88 gnd C_bl
Rb_49_89 bit_49_89 bit_49_90 R_bl
Rbb_49_89 bitb_49_89 bitb_49_90 R_bl
Cb_49_89 bit_49_89 gnd C_bl
Cbb_49_89 bitb_49_89 gnd C_bl
Rb_49_90 bit_49_90 bit_49_91 R_bl
Rbb_49_90 bitb_49_90 bitb_49_91 R_bl
Cb_49_90 bit_49_90 gnd C_bl
Cbb_49_90 bitb_49_90 gnd C_bl
Rb_49_91 bit_49_91 bit_49_92 R_bl
Rbb_49_91 bitb_49_91 bitb_49_92 R_bl
Cb_49_91 bit_49_91 gnd C_bl
Cbb_49_91 bitb_49_91 gnd C_bl
Rb_49_92 bit_49_92 bit_49_93 R_bl
Rbb_49_92 bitb_49_92 bitb_49_93 R_bl
Cb_49_92 bit_49_92 gnd C_bl
Cbb_49_92 bitb_49_92 gnd C_bl
Rb_49_93 bit_49_93 bit_49_94 R_bl
Rbb_49_93 bitb_49_93 bitb_49_94 R_bl
Cb_49_93 bit_49_93 gnd C_bl
Cbb_49_93 bitb_49_93 gnd C_bl
Rb_49_94 bit_49_94 bit_49_95 R_bl
Rbb_49_94 bitb_49_94 bitb_49_95 R_bl
Cb_49_94 bit_49_94 gnd C_bl
Cbb_49_94 bitb_49_94 gnd C_bl
Rb_49_95 bit_49_95 bit_49_96 R_bl
Rbb_49_95 bitb_49_95 bitb_49_96 R_bl
Cb_49_95 bit_49_95 gnd C_bl
Cbb_49_95 bitb_49_95 gnd C_bl
Rb_49_96 bit_49_96 bit_49_97 R_bl
Rbb_49_96 bitb_49_96 bitb_49_97 R_bl
Cb_49_96 bit_49_96 gnd C_bl
Cbb_49_96 bitb_49_96 gnd C_bl
Rb_49_97 bit_49_97 bit_49_98 R_bl
Rbb_49_97 bitb_49_97 bitb_49_98 R_bl
Cb_49_97 bit_49_97 gnd C_bl
Cbb_49_97 bitb_49_97 gnd C_bl
Rb_49_98 bit_49_98 bit_49_99 R_bl
Rbb_49_98 bitb_49_98 bitb_49_99 R_bl
Cb_49_98 bit_49_98 gnd C_bl
Cbb_49_98 bitb_49_98 gnd C_bl
Rb_49_99 bit_49_99 bit_49_100 R_bl
Rbb_49_99 bitb_49_99 bitb_49_100 R_bl
Cb_49_99 bit_49_99 gnd C_bl
Cbb_49_99 bitb_49_99 gnd C_bl
Rb_50_0 bit_50_0 bit_50_1 R_bl
Rbb_50_0 bitb_50_0 bitb_50_1 R_bl
Cb_50_0 bit_50_0 gnd C_bl
Cbb_50_0 bitb_50_0 gnd C_bl
Rb_50_1 bit_50_1 bit_50_2 R_bl
Rbb_50_1 bitb_50_1 bitb_50_2 R_bl
Cb_50_1 bit_50_1 gnd C_bl
Cbb_50_1 bitb_50_1 gnd C_bl
Rb_50_2 bit_50_2 bit_50_3 R_bl
Rbb_50_2 bitb_50_2 bitb_50_3 R_bl
Cb_50_2 bit_50_2 gnd C_bl
Cbb_50_2 bitb_50_2 gnd C_bl
Rb_50_3 bit_50_3 bit_50_4 R_bl
Rbb_50_3 bitb_50_3 bitb_50_4 R_bl
Cb_50_3 bit_50_3 gnd C_bl
Cbb_50_3 bitb_50_3 gnd C_bl
Rb_50_4 bit_50_4 bit_50_5 R_bl
Rbb_50_4 bitb_50_4 bitb_50_5 R_bl
Cb_50_4 bit_50_4 gnd C_bl
Cbb_50_4 bitb_50_4 gnd C_bl
Rb_50_5 bit_50_5 bit_50_6 R_bl
Rbb_50_5 bitb_50_5 bitb_50_6 R_bl
Cb_50_5 bit_50_5 gnd C_bl
Cbb_50_5 bitb_50_5 gnd C_bl
Rb_50_6 bit_50_6 bit_50_7 R_bl
Rbb_50_6 bitb_50_6 bitb_50_7 R_bl
Cb_50_6 bit_50_6 gnd C_bl
Cbb_50_6 bitb_50_6 gnd C_bl
Rb_50_7 bit_50_7 bit_50_8 R_bl
Rbb_50_7 bitb_50_7 bitb_50_8 R_bl
Cb_50_7 bit_50_7 gnd C_bl
Cbb_50_7 bitb_50_7 gnd C_bl
Rb_50_8 bit_50_8 bit_50_9 R_bl
Rbb_50_8 bitb_50_8 bitb_50_9 R_bl
Cb_50_8 bit_50_8 gnd C_bl
Cbb_50_8 bitb_50_8 gnd C_bl
Rb_50_9 bit_50_9 bit_50_10 R_bl
Rbb_50_9 bitb_50_9 bitb_50_10 R_bl
Cb_50_9 bit_50_9 gnd C_bl
Cbb_50_9 bitb_50_9 gnd C_bl
Rb_50_10 bit_50_10 bit_50_11 R_bl
Rbb_50_10 bitb_50_10 bitb_50_11 R_bl
Cb_50_10 bit_50_10 gnd C_bl
Cbb_50_10 bitb_50_10 gnd C_bl
Rb_50_11 bit_50_11 bit_50_12 R_bl
Rbb_50_11 bitb_50_11 bitb_50_12 R_bl
Cb_50_11 bit_50_11 gnd C_bl
Cbb_50_11 bitb_50_11 gnd C_bl
Rb_50_12 bit_50_12 bit_50_13 R_bl
Rbb_50_12 bitb_50_12 bitb_50_13 R_bl
Cb_50_12 bit_50_12 gnd C_bl
Cbb_50_12 bitb_50_12 gnd C_bl
Rb_50_13 bit_50_13 bit_50_14 R_bl
Rbb_50_13 bitb_50_13 bitb_50_14 R_bl
Cb_50_13 bit_50_13 gnd C_bl
Cbb_50_13 bitb_50_13 gnd C_bl
Rb_50_14 bit_50_14 bit_50_15 R_bl
Rbb_50_14 bitb_50_14 bitb_50_15 R_bl
Cb_50_14 bit_50_14 gnd C_bl
Cbb_50_14 bitb_50_14 gnd C_bl
Rb_50_15 bit_50_15 bit_50_16 R_bl
Rbb_50_15 bitb_50_15 bitb_50_16 R_bl
Cb_50_15 bit_50_15 gnd C_bl
Cbb_50_15 bitb_50_15 gnd C_bl
Rb_50_16 bit_50_16 bit_50_17 R_bl
Rbb_50_16 bitb_50_16 bitb_50_17 R_bl
Cb_50_16 bit_50_16 gnd C_bl
Cbb_50_16 bitb_50_16 gnd C_bl
Rb_50_17 bit_50_17 bit_50_18 R_bl
Rbb_50_17 bitb_50_17 bitb_50_18 R_bl
Cb_50_17 bit_50_17 gnd C_bl
Cbb_50_17 bitb_50_17 gnd C_bl
Rb_50_18 bit_50_18 bit_50_19 R_bl
Rbb_50_18 bitb_50_18 bitb_50_19 R_bl
Cb_50_18 bit_50_18 gnd C_bl
Cbb_50_18 bitb_50_18 gnd C_bl
Rb_50_19 bit_50_19 bit_50_20 R_bl
Rbb_50_19 bitb_50_19 bitb_50_20 R_bl
Cb_50_19 bit_50_19 gnd C_bl
Cbb_50_19 bitb_50_19 gnd C_bl
Rb_50_20 bit_50_20 bit_50_21 R_bl
Rbb_50_20 bitb_50_20 bitb_50_21 R_bl
Cb_50_20 bit_50_20 gnd C_bl
Cbb_50_20 bitb_50_20 gnd C_bl
Rb_50_21 bit_50_21 bit_50_22 R_bl
Rbb_50_21 bitb_50_21 bitb_50_22 R_bl
Cb_50_21 bit_50_21 gnd C_bl
Cbb_50_21 bitb_50_21 gnd C_bl
Rb_50_22 bit_50_22 bit_50_23 R_bl
Rbb_50_22 bitb_50_22 bitb_50_23 R_bl
Cb_50_22 bit_50_22 gnd C_bl
Cbb_50_22 bitb_50_22 gnd C_bl
Rb_50_23 bit_50_23 bit_50_24 R_bl
Rbb_50_23 bitb_50_23 bitb_50_24 R_bl
Cb_50_23 bit_50_23 gnd C_bl
Cbb_50_23 bitb_50_23 gnd C_bl
Rb_50_24 bit_50_24 bit_50_25 R_bl
Rbb_50_24 bitb_50_24 bitb_50_25 R_bl
Cb_50_24 bit_50_24 gnd C_bl
Cbb_50_24 bitb_50_24 gnd C_bl
Rb_50_25 bit_50_25 bit_50_26 R_bl
Rbb_50_25 bitb_50_25 bitb_50_26 R_bl
Cb_50_25 bit_50_25 gnd C_bl
Cbb_50_25 bitb_50_25 gnd C_bl
Rb_50_26 bit_50_26 bit_50_27 R_bl
Rbb_50_26 bitb_50_26 bitb_50_27 R_bl
Cb_50_26 bit_50_26 gnd C_bl
Cbb_50_26 bitb_50_26 gnd C_bl
Rb_50_27 bit_50_27 bit_50_28 R_bl
Rbb_50_27 bitb_50_27 bitb_50_28 R_bl
Cb_50_27 bit_50_27 gnd C_bl
Cbb_50_27 bitb_50_27 gnd C_bl
Rb_50_28 bit_50_28 bit_50_29 R_bl
Rbb_50_28 bitb_50_28 bitb_50_29 R_bl
Cb_50_28 bit_50_28 gnd C_bl
Cbb_50_28 bitb_50_28 gnd C_bl
Rb_50_29 bit_50_29 bit_50_30 R_bl
Rbb_50_29 bitb_50_29 bitb_50_30 R_bl
Cb_50_29 bit_50_29 gnd C_bl
Cbb_50_29 bitb_50_29 gnd C_bl
Rb_50_30 bit_50_30 bit_50_31 R_bl
Rbb_50_30 bitb_50_30 bitb_50_31 R_bl
Cb_50_30 bit_50_30 gnd C_bl
Cbb_50_30 bitb_50_30 gnd C_bl
Rb_50_31 bit_50_31 bit_50_32 R_bl
Rbb_50_31 bitb_50_31 bitb_50_32 R_bl
Cb_50_31 bit_50_31 gnd C_bl
Cbb_50_31 bitb_50_31 gnd C_bl
Rb_50_32 bit_50_32 bit_50_33 R_bl
Rbb_50_32 bitb_50_32 bitb_50_33 R_bl
Cb_50_32 bit_50_32 gnd C_bl
Cbb_50_32 bitb_50_32 gnd C_bl
Rb_50_33 bit_50_33 bit_50_34 R_bl
Rbb_50_33 bitb_50_33 bitb_50_34 R_bl
Cb_50_33 bit_50_33 gnd C_bl
Cbb_50_33 bitb_50_33 gnd C_bl
Rb_50_34 bit_50_34 bit_50_35 R_bl
Rbb_50_34 bitb_50_34 bitb_50_35 R_bl
Cb_50_34 bit_50_34 gnd C_bl
Cbb_50_34 bitb_50_34 gnd C_bl
Rb_50_35 bit_50_35 bit_50_36 R_bl
Rbb_50_35 bitb_50_35 bitb_50_36 R_bl
Cb_50_35 bit_50_35 gnd C_bl
Cbb_50_35 bitb_50_35 gnd C_bl
Rb_50_36 bit_50_36 bit_50_37 R_bl
Rbb_50_36 bitb_50_36 bitb_50_37 R_bl
Cb_50_36 bit_50_36 gnd C_bl
Cbb_50_36 bitb_50_36 gnd C_bl
Rb_50_37 bit_50_37 bit_50_38 R_bl
Rbb_50_37 bitb_50_37 bitb_50_38 R_bl
Cb_50_37 bit_50_37 gnd C_bl
Cbb_50_37 bitb_50_37 gnd C_bl
Rb_50_38 bit_50_38 bit_50_39 R_bl
Rbb_50_38 bitb_50_38 bitb_50_39 R_bl
Cb_50_38 bit_50_38 gnd C_bl
Cbb_50_38 bitb_50_38 gnd C_bl
Rb_50_39 bit_50_39 bit_50_40 R_bl
Rbb_50_39 bitb_50_39 bitb_50_40 R_bl
Cb_50_39 bit_50_39 gnd C_bl
Cbb_50_39 bitb_50_39 gnd C_bl
Rb_50_40 bit_50_40 bit_50_41 R_bl
Rbb_50_40 bitb_50_40 bitb_50_41 R_bl
Cb_50_40 bit_50_40 gnd C_bl
Cbb_50_40 bitb_50_40 gnd C_bl
Rb_50_41 bit_50_41 bit_50_42 R_bl
Rbb_50_41 bitb_50_41 bitb_50_42 R_bl
Cb_50_41 bit_50_41 gnd C_bl
Cbb_50_41 bitb_50_41 gnd C_bl
Rb_50_42 bit_50_42 bit_50_43 R_bl
Rbb_50_42 bitb_50_42 bitb_50_43 R_bl
Cb_50_42 bit_50_42 gnd C_bl
Cbb_50_42 bitb_50_42 gnd C_bl
Rb_50_43 bit_50_43 bit_50_44 R_bl
Rbb_50_43 bitb_50_43 bitb_50_44 R_bl
Cb_50_43 bit_50_43 gnd C_bl
Cbb_50_43 bitb_50_43 gnd C_bl
Rb_50_44 bit_50_44 bit_50_45 R_bl
Rbb_50_44 bitb_50_44 bitb_50_45 R_bl
Cb_50_44 bit_50_44 gnd C_bl
Cbb_50_44 bitb_50_44 gnd C_bl
Rb_50_45 bit_50_45 bit_50_46 R_bl
Rbb_50_45 bitb_50_45 bitb_50_46 R_bl
Cb_50_45 bit_50_45 gnd C_bl
Cbb_50_45 bitb_50_45 gnd C_bl
Rb_50_46 bit_50_46 bit_50_47 R_bl
Rbb_50_46 bitb_50_46 bitb_50_47 R_bl
Cb_50_46 bit_50_46 gnd C_bl
Cbb_50_46 bitb_50_46 gnd C_bl
Rb_50_47 bit_50_47 bit_50_48 R_bl
Rbb_50_47 bitb_50_47 bitb_50_48 R_bl
Cb_50_47 bit_50_47 gnd C_bl
Cbb_50_47 bitb_50_47 gnd C_bl
Rb_50_48 bit_50_48 bit_50_49 R_bl
Rbb_50_48 bitb_50_48 bitb_50_49 R_bl
Cb_50_48 bit_50_48 gnd C_bl
Cbb_50_48 bitb_50_48 gnd C_bl
Rb_50_49 bit_50_49 bit_50_50 R_bl
Rbb_50_49 bitb_50_49 bitb_50_50 R_bl
Cb_50_49 bit_50_49 gnd C_bl
Cbb_50_49 bitb_50_49 gnd C_bl
Rb_50_50 bit_50_50 bit_50_51 R_bl
Rbb_50_50 bitb_50_50 bitb_50_51 R_bl
Cb_50_50 bit_50_50 gnd C_bl
Cbb_50_50 bitb_50_50 gnd C_bl
Rb_50_51 bit_50_51 bit_50_52 R_bl
Rbb_50_51 bitb_50_51 bitb_50_52 R_bl
Cb_50_51 bit_50_51 gnd C_bl
Cbb_50_51 bitb_50_51 gnd C_bl
Rb_50_52 bit_50_52 bit_50_53 R_bl
Rbb_50_52 bitb_50_52 bitb_50_53 R_bl
Cb_50_52 bit_50_52 gnd C_bl
Cbb_50_52 bitb_50_52 gnd C_bl
Rb_50_53 bit_50_53 bit_50_54 R_bl
Rbb_50_53 bitb_50_53 bitb_50_54 R_bl
Cb_50_53 bit_50_53 gnd C_bl
Cbb_50_53 bitb_50_53 gnd C_bl
Rb_50_54 bit_50_54 bit_50_55 R_bl
Rbb_50_54 bitb_50_54 bitb_50_55 R_bl
Cb_50_54 bit_50_54 gnd C_bl
Cbb_50_54 bitb_50_54 gnd C_bl
Rb_50_55 bit_50_55 bit_50_56 R_bl
Rbb_50_55 bitb_50_55 bitb_50_56 R_bl
Cb_50_55 bit_50_55 gnd C_bl
Cbb_50_55 bitb_50_55 gnd C_bl
Rb_50_56 bit_50_56 bit_50_57 R_bl
Rbb_50_56 bitb_50_56 bitb_50_57 R_bl
Cb_50_56 bit_50_56 gnd C_bl
Cbb_50_56 bitb_50_56 gnd C_bl
Rb_50_57 bit_50_57 bit_50_58 R_bl
Rbb_50_57 bitb_50_57 bitb_50_58 R_bl
Cb_50_57 bit_50_57 gnd C_bl
Cbb_50_57 bitb_50_57 gnd C_bl
Rb_50_58 bit_50_58 bit_50_59 R_bl
Rbb_50_58 bitb_50_58 bitb_50_59 R_bl
Cb_50_58 bit_50_58 gnd C_bl
Cbb_50_58 bitb_50_58 gnd C_bl
Rb_50_59 bit_50_59 bit_50_60 R_bl
Rbb_50_59 bitb_50_59 bitb_50_60 R_bl
Cb_50_59 bit_50_59 gnd C_bl
Cbb_50_59 bitb_50_59 gnd C_bl
Rb_50_60 bit_50_60 bit_50_61 R_bl
Rbb_50_60 bitb_50_60 bitb_50_61 R_bl
Cb_50_60 bit_50_60 gnd C_bl
Cbb_50_60 bitb_50_60 gnd C_bl
Rb_50_61 bit_50_61 bit_50_62 R_bl
Rbb_50_61 bitb_50_61 bitb_50_62 R_bl
Cb_50_61 bit_50_61 gnd C_bl
Cbb_50_61 bitb_50_61 gnd C_bl
Rb_50_62 bit_50_62 bit_50_63 R_bl
Rbb_50_62 bitb_50_62 bitb_50_63 R_bl
Cb_50_62 bit_50_62 gnd C_bl
Cbb_50_62 bitb_50_62 gnd C_bl
Rb_50_63 bit_50_63 bit_50_64 R_bl
Rbb_50_63 bitb_50_63 bitb_50_64 R_bl
Cb_50_63 bit_50_63 gnd C_bl
Cbb_50_63 bitb_50_63 gnd C_bl
Rb_50_64 bit_50_64 bit_50_65 R_bl
Rbb_50_64 bitb_50_64 bitb_50_65 R_bl
Cb_50_64 bit_50_64 gnd C_bl
Cbb_50_64 bitb_50_64 gnd C_bl
Rb_50_65 bit_50_65 bit_50_66 R_bl
Rbb_50_65 bitb_50_65 bitb_50_66 R_bl
Cb_50_65 bit_50_65 gnd C_bl
Cbb_50_65 bitb_50_65 gnd C_bl
Rb_50_66 bit_50_66 bit_50_67 R_bl
Rbb_50_66 bitb_50_66 bitb_50_67 R_bl
Cb_50_66 bit_50_66 gnd C_bl
Cbb_50_66 bitb_50_66 gnd C_bl
Rb_50_67 bit_50_67 bit_50_68 R_bl
Rbb_50_67 bitb_50_67 bitb_50_68 R_bl
Cb_50_67 bit_50_67 gnd C_bl
Cbb_50_67 bitb_50_67 gnd C_bl
Rb_50_68 bit_50_68 bit_50_69 R_bl
Rbb_50_68 bitb_50_68 bitb_50_69 R_bl
Cb_50_68 bit_50_68 gnd C_bl
Cbb_50_68 bitb_50_68 gnd C_bl
Rb_50_69 bit_50_69 bit_50_70 R_bl
Rbb_50_69 bitb_50_69 bitb_50_70 R_bl
Cb_50_69 bit_50_69 gnd C_bl
Cbb_50_69 bitb_50_69 gnd C_bl
Rb_50_70 bit_50_70 bit_50_71 R_bl
Rbb_50_70 bitb_50_70 bitb_50_71 R_bl
Cb_50_70 bit_50_70 gnd C_bl
Cbb_50_70 bitb_50_70 gnd C_bl
Rb_50_71 bit_50_71 bit_50_72 R_bl
Rbb_50_71 bitb_50_71 bitb_50_72 R_bl
Cb_50_71 bit_50_71 gnd C_bl
Cbb_50_71 bitb_50_71 gnd C_bl
Rb_50_72 bit_50_72 bit_50_73 R_bl
Rbb_50_72 bitb_50_72 bitb_50_73 R_bl
Cb_50_72 bit_50_72 gnd C_bl
Cbb_50_72 bitb_50_72 gnd C_bl
Rb_50_73 bit_50_73 bit_50_74 R_bl
Rbb_50_73 bitb_50_73 bitb_50_74 R_bl
Cb_50_73 bit_50_73 gnd C_bl
Cbb_50_73 bitb_50_73 gnd C_bl
Rb_50_74 bit_50_74 bit_50_75 R_bl
Rbb_50_74 bitb_50_74 bitb_50_75 R_bl
Cb_50_74 bit_50_74 gnd C_bl
Cbb_50_74 bitb_50_74 gnd C_bl
Rb_50_75 bit_50_75 bit_50_76 R_bl
Rbb_50_75 bitb_50_75 bitb_50_76 R_bl
Cb_50_75 bit_50_75 gnd C_bl
Cbb_50_75 bitb_50_75 gnd C_bl
Rb_50_76 bit_50_76 bit_50_77 R_bl
Rbb_50_76 bitb_50_76 bitb_50_77 R_bl
Cb_50_76 bit_50_76 gnd C_bl
Cbb_50_76 bitb_50_76 gnd C_bl
Rb_50_77 bit_50_77 bit_50_78 R_bl
Rbb_50_77 bitb_50_77 bitb_50_78 R_bl
Cb_50_77 bit_50_77 gnd C_bl
Cbb_50_77 bitb_50_77 gnd C_bl
Rb_50_78 bit_50_78 bit_50_79 R_bl
Rbb_50_78 bitb_50_78 bitb_50_79 R_bl
Cb_50_78 bit_50_78 gnd C_bl
Cbb_50_78 bitb_50_78 gnd C_bl
Rb_50_79 bit_50_79 bit_50_80 R_bl
Rbb_50_79 bitb_50_79 bitb_50_80 R_bl
Cb_50_79 bit_50_79 gnd C_bl
Cbb_50_79 bitb_50_79 gnd C_bl
Rb_50_80 bit_50_80 bit_50_81 R_bl
Rbb_50_80 bitb_50_80 bitb_50_81 R_bl
Cb_50_80 bit_50_80 gnd C_bl
Cbb_50_80 bitb_50_80 gnd C_bl
Rb_50_81 bit_50_81 bit_50_82 R_bl
Rbb_50_81 bitb_50_81 bitb_50_82 R_bl
Cb_50_81 bit_50_81 gnd C_bl
Cbb_50_81 bitb_50_81 gnd C_bl
Rb_50_82 bit_50_82 bit_50_83 R_bl
Rbb_50_82 bitb_50_82 bitb_50_83 R_bl
Cb_50_82 bit_50_82 gnd C_bl
Cbb_50_82 bitb_50_82 gnd C_bl
Rb_50_83 bit_50_83 bit_50_84 R_bl
Rbb_50_83 bitb_50_83 bitb_50_84 R_bl
Cb_50_83 bit_50_83 gnd C_bl
Cbb_50_83 bitb_50_83 gnd C_bl
Rb_50_84 bit_50_84 bit_50_85 R_bl
Rbb_50_84 bitb_50_84 bitb_50_85 R_bl
Cb_50_84 bit_50_84 gnd C_bl
Cbb_50_84 bitb_50_84 gnd C_bl
Rb_50_85 bit_50_85 bit_50_86 R_bl
Rbb_50_85 bitb_50_85 bitb_50_86 R_bl
Cb_50_85 bit_50_85 gnd C_bl
Cbb_50_85 bitb_50_85 gnd C_bl
Rb_50_86 bit_50_86 bit_50_87 R_bl
Rbb_50_86 bitb_50_86 bitb_50_87 R_bl
Cb_50_86 bit_50_86 gnd C_bl
Cbb_50_86 bitb_50_86 gnd C_bl
Rb_50_87 bit_50_87 bit_50_88 R_bl
Rbb_50_87 bitb_50_87 bitb_50_88 R_bl
Cb_50_87 bit_50_87 gnd C_bl
Cbb_50_87 bitb_50_87 gnd C_bl
Rb_50_88 bit_50_88 bit_50_89 R_bl
Rbb_50_88 bitb_50_88 bitb_50_89 R_bl
Cb_50_88 bit_50_88 gnd C_bl
Cbb_50_88 bitb_50_88 gnd C_bl
Rb_50_89 bit_50_89 bit_50_90 R_bl
Rbb_50_89 bitb_50_89 bitb_50_90 R_bl
Cb_50_89 bit_50_89 gnd C_bl
Cbb_50_89 bitb_50_89 gnd C_bl
Rb_50_90 bit_50_90 bit_50_91 R_bl
Rbb_50_90 bitb_50_90 bitb_50_91 R_bl
Cb_50_90 bit_50_90 gnd C_bl
Cbb_50_90 bitb_50_90 gnd C_bl
Rb_50_91 bit_50_91 bit_50_92 R_bl
Rbb_50_91 bitb_50_91 bitb_50_92 R_bl
Cb_50_91 bit_50_91 gnd C_bl
Cbb_50_91 bitb_50_91 gnd C_bl
Rb_50_92 bit_50_92 bit_50_93 R_bl
Rbb_50_92 bitb_50_92 bitb_50_93 R_bl
Cb_50_92 bit_50_92 gnd C_bl
Cbb_50_92 bitb_50_92 gnd C_bl
Rb_50_93 bit_50_93 bit_50_94 R_bl
Rbb_50_93 bitb_50_93 bitb_50_94 R_bl
Cb_50_93 bit_50_93 gnd C_bl
Cbb_50_93 bitb_50_93 gnd C_bl
Rb_50_94 bit_50_94 bit_50_95 R_bl
Rbb_50_94 bitb_50_94 bitb_50_95 R_bl
Cb_50_94 bit_50_94 gnd C_bl
Cbb_50_94 bitb_50_94 gnd C_bl
Rb_50_95 bit_50_95 bit_50_96 R_bl
Rbb_50_95 bitb_50_95 bitb_50_96 R_bl
Cb_50_95 bit_50_95 gnd C_bl
Cbb_50_95 bitb_50_95 gnd C_bl
Rb_50_96 bit_50_96 bit_50_97 R_bl
Rbb_50_96 bitb_50_96 bitb_50_97 R_bl
Cb_50_96 bit_50_96 gnd C_bl
Cbb_50_96 bitb_50_96 gnd C_bl
Rb_50_97 bit_50_97 bit_50_98 R_bl
Rbb_50_97 bitb_50_97 bitb_50_98 R_bl
Cb_50_97 bit_50_97 gnd C_bl
Cbb_50_97 bitb_50_97 gnd C_bl
Rb_50_98 bit_50_98 bit_50_99 R_bl
Rbb_50_98 bitb_50_98 bitb_50_99 R_bl
Cb_50_98 bit_50_98 gnd C_bl
Cbb_50_98 bitb_50_98 gnd C_bl
Rb_50_99 bit_50_99 bit_50_100 R_bl
Rbb_50_99 bitb_50_99 bitb_50_100 R_bl
Cb_50_99 bit_50_99 gnd C_bl
Cbb_50_99 bitb_50_99 gnd C_bl
Rb_51_0 bit_51_0 bit_51_1 R_bl
Rbb_51_0 bitb_51_0 bitb_51_1 R_bl
Cb_51_0 bit_51_0 gnd C_bl
Cbb_51_0 bitb_51_0 gnd C_bl
Rb_51_1 bit_51_1 bit_51_2 R_bl
Rbb_51_1 bitb_51_1 bitb_51_2 R_bl
Cb_51_1 bit_51_1 gnd C_bl
Cbb_51_1 bitb_51_1 gnd C_bl
Rb_51_2 bit_51_2 bit_51_3 R_bl
Rbb_51_2 bitb_51_2 bitb_51_3 R_bl
Cb_51_2 bit_51_2 gnd C_bl
Cbb_51_2 bitb_51_2 gnd C_bl
Rb_51_3 bit_51_3 bit_51_4 R_bl
Rbb_51_3 bitb_51_3 bitb_51_4 R_bl
Cb_51_3 bit_51_3 gnd C_bl
Cbb_51_3 bitb_51_3 gnd C_bl
Rb_51_4 bit_51_4 bit_51_5 R_bl
Rbb_51_4 bitb_51_4 bitb_51_5 R_bl
Cb_51_4 bit_51_4 gnd C_bl
Cbb_51_4 bitb_51_4 gnd C_bl
Rb_51_5 bit_51_5 bit_51_6 R_bl
Rbb_51_5 bitb_51_5 bitb_51_6 R_bl
Cb_51_5 bit_51_5 gnd C_bl
Cbb_51_5 bitb_51_5 gnd C_bl
Rb_51_6 bit_51_6 bit_51_7 R_bl
Rbb_51_6 bitb_51_6 bitb_51_7 R_bl
Cb_51_6 bit_51_6 gnd C_bl
Cbb_51_6 bitb_51_6 gnd C_bl
Rb_51_7 bit_51_7 bit_51_8 R_bl
Rbb_51_7 bitb_51_7 bitb_51_8 R_bl
Cb_51_7 bit_51_7 gnd C_bl
Cbb_51_7 bitb_51_7 gnd C_bl
Rb_51_8 bit_51_8 bit_51_9 R_bl
Rbb_51_8 bitb_51_8 bitb_51_9 R_bl
Cb_51_8 bit_51_8 gnd C_bl
Cbb_51_8 bitb_51_8 gnd C_bl
Rb_51_9 bit_51_9 bit_51_10 R_bl
Rbb_51_9 bitb_51_9 bitb_51_10 R_bl
Cb_51_9 bit_51_9 gnd C_bl
Cbb_51_9 bitb_51_9 gnd C_bl
Rb_51_10 bit_51_10 bit_51_11 R_bl
Rbb_51_10 bitb_51_10 bitb_51_11 R_bl
Cb_51_10 bit_51_10 gnd C_bl
Cbb_51_10 bitb_51_10 gnd C_bl
Rb_51_11 bit_51_11 bit_51_12 R_bl
Rbb_51_11 bitb_51_11 bitb_51_12 R_bl
Cb_51_11 bit_51_11 gnd C_bl
Cbb_51_11 bitb_51_11 gnd C_bl
Rb_51_12 bit_51_12 bit_51_13 R_bl
Rbb_51_12 bitb_51_12 bitb_51_13 R_bl
Cb_51_12 bit_51_12 gnd C_bl
Cbb_51_12 bitb_51_12 gnd C_bl
Rb_51_13 bit_51_13 bit_51_14 R_bl
Rbb_51_13 bitb_51_13 bitb_51_14 R_bl
Cb_51_13 bit_51_13 gnd C_bl
Cbb_51_13 bitb_51_13 gnd C_bl
Rb_51_14 bit_51_14 bit_51_15 R_bl
Rbb_51_14 bitb_51_14 bitb_51_15 R_bl
Cb_51_14 bit_51_14 gnd C_bl
Cbb_51_14 bitb_51_14 gnd C_bl
Rb_51_15 bit_51_15 bit_51_16 R_bl
Rbb_51_15 bitb_51_15 bitb_51_16 R_bl
Cb_51_15 bit_51_15 gnd C_bl
Cbb_51_15 bitb_51_15 gnd C_bl
Rb_51_16 bit_51_16 bit_51_17 R_bl
Rbb_51_16 bitb_51_16 bitb_51_17 R_bl
Cb_51_16 bit_51_16 gnd C_bl
Cbb_51_16 bitb_51_16 gnd C_bl
Rb_51_17 bit_51_17 bit_51_18 R_bl
Rbb_51_17 bitb_51_17 bitb_51_18 R_bl
Cb_51_17 bit_51_17 gnd C_bl
Cbb_51_17 bitb_51_17 gnd C_bl
Rb_51_18 bit_51_18 bit_51_19 R_bl
Rbb_51_18 bitb_51_18 bitb_51_19 R_bl
Cb_51_18 bit_51_18 gnd C_bl
Cbb_51_18 bitb_51_18 gnd C_bl
Rb_51_19 bit_51_19 bit_51_20 R_bl
Rbb_51_19 bitb_51_19 bitb_51_20 R_bl
Cb_51_19 bit_51_19 gnd C_bl
Cbb_51_19 bitb_51_19 gnd C_bl
Rb_51_20 bit_51_20 bit_51_21 R_bl
Rbb_51_20 bitb_51_20 bitb_51_21 R_bl
Cb_51_20 bit_51_20 gnd C_bl
Cbb_51_20 bitb_51_20 gnd C_bl
Rb_51_21 bit_51_21 bit_51_22 R_bl
Rbb_51_21 bitb_51_21 bitb_51_22 R_bl
Cb_51_21 bit_51_21 gnd C_bl
Cbb_51_21 bitb_51_21 gnd C_bl
Rb_51_22 bit_51_22 bit_51_23 R_bl
Rbb_51_22 bitb_51_22 bitb_51_23 R_bl
Cb_51_22 bit_51_22 gnd C_bl
Cbb_51_22 bitb_51_22 gnd C_bl
Rb_51_23 bit_51_23 bit_51_24 R_bl
Rbb_51_23 bitb_51_23 bitb_51_24 R_bl
Cb_51_23 bit_51_23 gnd C_bl
Cbb_51_23 bitb_51_23 gnd C_bl
Rb_51_24 bit_51_24 bit_51_25 R_bl
Rbb_51_24 bitb_51_24 bitb_51_25 R_bl
Cb_51_24 bit_51_24 gnd C_bl
Cbb_51_24 bitb_51_24 gnd C_bl
Rb_51_25 bit_51_25 bit_51_26 R_bl
Rbb_51_25 bitb_51_25 bitb_51_26 R_bl
Cb_51_25 bit_51_25 gnd C_bl
Cbb_51_25 bitb_51_25 gnd C_bl
Rb_51_26 bit_51_26 bit_51_27 R_bl
Rbb_51_26 bitb_51_26 bitb_51_27 R_bl
Cb_51_26 bit_51_26 gnd C_bl
Cbb_51_26 bitb_51_26 gnd C_bl
Rb_51_27 bit_51_27 bit_51_28 R_bl
Rbb_51_27 bitb_51_27 bitb_51_28 R_bl
Cb_51_27 bit_51_27 gnd C_bl
Cbb_51_27 bitb_51_27 gnd C_bl
Rb_51_28 bit_51_28 bit_51_29 R_bl
Rbb_51_28 bitb_51_28 bitb_51_29 R_bl
Cb_51_28 bit_51_28 gnd C_bl
Cbb_51_28 bitb_51_28 gnd C_bl
Rb_51_29 bit_51_29 bit_51_30 R_bl
Rbb_51_29 bitb_51_29 bitb_51_30 R_bl
Cb_51_29 bit_51_29 gnd C_bl
Cbb_51_29 bitb_51_29 gnd C_bl
Rb_51_30 bit_51_30 bit_51_31 R_bl
Rbb_51_30 bitb_51_30 bitb_51_31 R_bl
Cb_51_30 bit_51_30 gnd C_bl
Cbb_51_30 bitb_51_30 gnd C_bl
Rb_51_31 bit_51_31 bit_51_32 R_bl
Rbb_51_31 bitb_51_31 bitb_51_32 R_bl
Cb_51_31 bit_51_31 gnd C_bl
Cbb_51_31 bitb_51_31 gnd C_bl
Rb_51_32 bit_51_32 bit_51_33 R_bl
Rbb_51_32 bitb_51_32 bitb_51_33 R_bl
Cb_51_32 bit_51_32 gnd C_bl
Cbb_51_32 bitb_51_32 gnd C_bl
Rb_51_33 bit_51_33 bit_51_34 R_bl
Rbb_51_33 bitb_51_33 bitb_51_34 R_bl
Cb_51_33 bit_51_33 gnd C_bl
Cbb_51_33 bitb_51_33 gnd C_bl
Rb_51_34 bit_51_34 bit_51_35 R_bl
Rbb_51_34 bitb_51_34 bitb_51_35 R_bl
Cb_51_34 bit_51_34 gnd C_bl
Cbb_51_34 bitb_51_34 gnd C_bl
Rb_51_35 bit_51_35 bit_51_36 R_bl
Rbb_51_35 bitb_51_35 bitb_51_36 R_bl
Cb_51_35 bit_51_35 gnd C_bl
Cbb_51_35 bitb_51_35 gnd C_bl
Rb_51_36 bit_51_36 bit_51_37 R_bl
Rbb_51_36 bitb_51_36 bitb_51_37 R_bl
Cb_51_36 bit_51_36 gnd C_bl
Cbb_51_36 bitb_51_36 gnd C_bl
Rb_51_37 bit_51_37 bit_51_38 R_bl
Rbb_51_37 bitb_51_37 bitb_51_38 R_bl
Cb_51_37 bit_51_37 gnd C_bl
Cbb_51_37 bitb_51_37 gnd C_bl
Rb_51_38 bit_51_38 bit_51_39 R_bl
Rbb_51_38 bitb_51_38 bitb_51_39 R_bl
Cb_51_38 bit_51_38 gnd C_bl
Cbb_51_38 bitb_51_38 gnd C_bl
Rb_51_39 bit_51_39 bit_51_40 R_bl
Rbb_51_39 bitb_51_39 bitb_51_40 R_bl
Cb_51_39 bit_51_39 gnd C_bl
Cbb_51_39 bitb_51_39 gnd C_bl
Rb_51_40 bit_51_40 bit_51_41 R_bl
Rbb_51_40 bitb_51_40 bitb_51_41 R_bl
Cb_51_40 bit_51_40 gnd C_bl
Cbb_51_40 bitb_51_40 gnd C_bl
Rb_51_41 bit_51_41 bit_51_42 R_bl
Rbb_51_41 bitb_51_41 bitb_51_42 R_bl
Cb_51_41 bit_51_41 gnd C_bl
Cbb_51_41 bitb_51_41 gnd C_bl
Rb_51_42 bit_51_42 bit_51_43 R_bl
Rbb_51_42 bitb_51_42 bitb_51_43 R_bl
Cb_51_42 bit_51_42 gnd C_bl
Cbb_51_42 bitb_51_42 gnd C_bl
Rb_51_43 bit_51_43 bit_51_44 R_bl
Rbb_51_43 bitb_51_43 bitb_51_44 R_bl
Cb_51_43 bit_51_43 gnd C_bl
Cbb_51_43 bitb_51_43 gnd C_bl
Rb_51_44 bit_51_44 bit_51_45 R_bl
Rbb_51_44 bitb_51_44 bitb_51_45 R_bl
Cb_51_44 bit_51_44 gnd C_bl
Cbb_51_44 bitb_51_44 gnd C_bl
Rb_51_45 bit_51_45 bit_51_46 R_bl
Rbb_51_45 bitb_51_45 bitb_51_46 R_bl
Cb_51_45 bit_51_45 gnd C_bl
Cbb_51_45 bitb_51_45 gnd C_bl
Rb_51_46 bit_51_46 bit_51_47 R_bl
Rbb_51_46 bitb_51_46 bitb_51_47 R_bl
Cb_51_46 bit_51_46 gnd C_bl
Cbb_51_46 bitb_51_46 gnd C_bl
Rb_51_47 bit_51_47 bit_51_48 R_bl
Rbb_51_47 bitb_51_47 bitb_51_48 R_bl
Cb_51_47 bit_51_47 gnd C_bl
Cbb_51_47 bitb_51_47 gnd C_bl
Rb_51_48 bit_51_48 bit_51_49 R_bl
Rbb_51_48 bitb_51_48 bitb_51_49 R_bl
Cb_51_48 bit_51_48 gnd C_bl
Cbb_51_48 bitb_51_48 gnd C_bl
Rb_51_49 bit_51_49 bit_51_50 R_bl
Rbb_51_49 bitb_51_49 bitb_51_50 R_bl
Cb_51_49 bit_51_49 gnd C_bl
Cbb_51_49 bitb_51_49 gnd C_bl
Rb_51_50 bit_51_50 bit_51_51 R_bl
Rbb_51_50 bitb_51_50 bitb_51_51 R_bl
Cb_51_50 bit_51_50 gnd C_bl
Cbb_51_50 bitb_51_50 gnd C_bl
Rb_51_51 bit_51_51 bit_51_52 R_bl
Rbb_51_51 bitb_51_51 bitb_51_52 R_bl
Cb_51_51 bit_51_51 gnd C_bl
Cbb_51_51 bitb_51_51 gnd C_bl
Rb_51_52 bit_51_52 bit_51_53 R_bl
Rbb_51_52 bitb_51_52 bitb_51_53 R_bl
Cb_51_52 bit_51_52 gnd C_bl
Cbb_51_52 bitb_51_52 gnd C_bl
Rb_51_53 bit_51_53 bit_51_54 R_bl
Rbb_51_53 bitb_51_53 bitb_51_54 R_bl
Cb_51_53 bit_51_53 gnd C_bl
Cbb_51_53 bitb_51_53 gnd C_bl
Rb_51_54 bit_51_54 bit_51_55 R_bl
Rbb_51_54 bitb_51_54 bitb_51_55 R_bl
Cb_51_54 bit_51_54 gnd C_bl
Cbb_51_54 bitb_51_54 gnd C_bl
Rb_51_55 bit_51_55 bit_51_56 R_bl
Rbb_51_55 bitb_51_55 bitb_51_56 R_bl
Cb_51_55 bit_51_55 gnd C_bl
Cbb_51_55 bitb_51_55 gnd C_bl
Rb_51_56 bit_51_56 bit_51_57 R_bl
Rbb_51_56 bitb_51_56 bitb_51_57 R_bl
Cb_51_56 bit_51_56 gnd C_bl
Cbb_51_56 bitb_51_56 gnd C_bl
Rb_51_57 bit_51_57 bit_51_58 R_bl
Rbb_51_57 bitb_51_57 bitb_51_58 R_bl
Cb_51_57 bit_51_57 gnd C_bl
Cbb_51_57 bitb_51_57 gnd C_bl
Rb_51_58 bit_51_58 bit_51_59 R_bl
Rbb_51_58 bitb_51_58 bitb_51_59 R_bl
Cb_51_58 bit_51_58 gnd C_bl
Cbb_51_58 bitb_51_58 gnd C_bl
Rb_51_59 bit_51_59 bit_51_60 R_bl
Rbb_51_59 bitb_51_59 bitb_51_60 R_bl
Cb_51_59 bit_51_59 gnd C_bl
Cbb_51_59 bitb_51_59 gnd C_bl
Rb_51_60 bit_51_60 bit_51_61 R_bl
Rbb_51_60 bitb_51_60 bitb_51_61 R_bl
Cb_51_60 bit_51_60 gnd C_bl
Cbb_51_60 bitb_51_60 gnd C_bl
Rb_51_61 bit_51_61 bit_51_62 R_bl
Rbb_51_61 bitb_51_61 bitb_51_62 R_bl
Cb_51_61 bit_51_61 gnd C_bl
Cbb_51_61 bitb_51_61 gnd C_bl
Rb_51_62 bit_51_62 bit_51_63 R_bl
Rbb_51_62 bitb_51_62 bitb_51_63 R_bl
Cb_51_62 bit_51_62 gnd C_bl
Cbb_51_62 bitb_51_62 gnd C_bl
Rb_51_63 bit_51_63 bit_51_64 R_bl
Rbb_51_63 bitb_51_63 bitb_51_64 R_bl
Cb_51_63 bit_51_63 gnd C_bl
Cbb_51_63 bitb_51_63 gnd C_bl
Rb_51_64 bit_51_64 bit_51_65 R_bl
Rbb_51_64 bitb_51_64 bitb_51_65 R_bl
Cb_51_64 bit_51_64 gnd C_bl
Cbb_51_64 bitb_51_64 gnd C_bl
Rb_51_65 bit_51_65 bit_51_66 R_bl
Rbb_51_65 bitb_51_65 bitb_51_66 R_bl
Cb_51_65 bit_51_65 gnd C_bl
Cbb_51_65 bitb_51_65 gnd C_bl
Rb_51_66 bit_51_66 bit_51_67 R_bl
Rbb_51_66 bitb_51_66 bitb_51_67 R_bl
Cb_51_66 bit_51_66 gnd C_bl
Cbb_51_66 bitb_51_66 gnd C_bl
Rb_51_67 bit_51_67 bit_51_68 R_bl
Rbb_51_67 bitb_51_67 bitb_51_68 R_bl
Cb_51_67 bit_51_67 gnd C_bl
Cbb_51_67 bitb_51_67 gnd C_bl
Rb_51_68 bit_51_68 bit_51_69 R_bl
Rbb_51_68 bitb_51_68 bitb_51_69 R_bl
Cb_51_68 bit_51_68 gnd C_bl
Cbb_51_68 bitb_51_68 gnd C_bl
Rb_51_69 bit_51_69 bit_51_70 R_bl
Rbb_51_69 bitb_51_69 bitb_51_70 R_bl
Cb_51_69 bit_51_69 gnd C_bl
Cbb_51_69 bitb_51_69 gnd C_bl
Rb_51_70 bit_51_70 bit_51_71 R_bl
Rbb_51_70 bitb_51_70 bitb_51_71 R_bl
Cb_51_70 bit_51_70 gnd C_bl
Cbb_51_70 bitb_51_70 gnd C_bl
Rb_51_71 bit_51_71 bit_51_72 R_bl
Rbb_51_71 bitb_51_71 bitb_51_72 R_bl
Cb_51_71 bit_51_71 gnd C_bl
Cbb_51_71 bitb_51_71 gnd C_bl
Rb_51_72 bit_51_72 bit_51_73 R_bl
Rbb_51_72 bitb_51_72 bitb_51_73 R_bl
Cb_51_72 bit_51_72 gnd C_bl
Cbb_51_72 bitb_51_72 gnd C_bl
Rb_51_73 bit_51_73 bit_51_74 R_bl
Rbb_51_73 bitb_51_73 bitb_51_74 R_bl
Cb_51_73 bit_51_73 gnd C_bl
Cbb_51_73 bitb_51_73 gnd C_bl
Rb_51_74 bit_51_74 bit_51_75 R_bl
Rbb_51_74 bitb_51_74 bitb_51_75 R_bl
Cb_51_74 bit_51_74 gnd C_bl
Cbb_51_74 bitb_51_74 gnd C_bl
Rb_51_75 bit_51_75 bit_51_76 R_bl
Rbb_51_75 bitb_51_75 bitb_51_76 R_bl
Cb_51_75 bit_51_75 gnd C_bl
Cbb_51_75 bitb_51_75 gnd C_bl
Rb_51_76 bit_51_76 bit_51_77 R_bl
Rbb_51_76 bitb_51_76 bitb_51_77 R_bl
Cb_51_76 bit_51_76 gnd C_bl
Cbb_51_76 bitb_51_76 gnd C_bl
Rb_51_77 bit_51_77 bit_51_78 R_bl
Rbb_51_77 bitb_51_77 bitb_51_78 R_bl
Cb_51_77 bit_51_77 gnd C_bl
Cbb_51_77 bitb_51_77 gnd C_bl
Rb_51_78 bit_51_78 bit_51_79 R_bl
Rbb_51_78 bitb_51_78 bitb_51_79 R_bl
Cb_51_78 bit_51_78 gnd C_bl
Cbb_51_78 bitb_51_78 gnd C_bl
Rb_51_79 bit_51_79 bit_51_80 R_bl
Rbb_51_79 bitb_51_79 bitb_51_80 R_bl
Cb_51_79 bit_51_79 gnd C_bl
Cbb_51_79 bitb_51_79 gnd C_bl
Rb_51_80 bit_51_80 bit_51_81 R_bl
Rbb_51_80 bitb_51_80 bitb_51_81 R_bl
Cb_51_80 bit_51_80 gnd C_bl
Cbb_51_80 bitb_51_80 gnd C_bl
Rb_51_81 bit_51_81 bit_51_82 R_bl
Rbb_51_81 bitb_51_81 bitb_51_82 R_bl
Cb_51_81 bit_51_81 gnd C_bl
Cbb_51_81 bitb_51_81 gnd C_bl
Rb_51_82 bit_51_82 bit_51_83 R_bl
Rbb_51_82 bitb_51_82 bitb_51_83 R_bl
Cb_51_82 bit_51_82 gnd C_bl
Cbb_51_82 bitb_51_82 gnd C_bl
Rb_51_83 bit_51_83 bit_51_84 R_bl
Rbb_51_83 bitb_51_83 bitb_51_84 R_bl
Cb_51_83 bit_51_83 gnd C_bl
Cbb_51_83 bitb_51_83 gnd C_bl
Rb_51_84 bit_51_84 bit_51_85 R_bl
Rbb_51_84 bitb_51_84 bitb_51_85 R_bl
Cb_51_84 bit_51_84 gnd C_bl
Cbb_51_84 bitb_51_84 gnd C_bl
Rb_51_85 bit_51_85 bit_51_86 R_bl
Rbb_51_85 bitb_51_85 bitb_51_86 R_bl
Cb_51_85 bit_51_85 gnd C_bl
Cbb_51_85 bitb_51_85 gnd C_bl
Rb_51_86 bit_51_86 bit_51_87 R_bl
Rbb_51_86 bitb_51_86 bitb_51_87 R_bl
Cb_51_86 bit_51_86 gnd C_bl
Cbb_51_86 bitb_51_86 gnd C_bl
Rb_51_87 bit_51_87 bit_51_88 R_bl
Rbb_51_87 bitb_51_87 bitb_51_88 R_bl
Cb_51_87 bit_51_87 gnd C_bl
Cbb_51_87 bitb_51_87 gnd C_bl
Rb_51_88 bit_51_88 bit_51_89 R_bl
Rbb_51_88 bitb_51_88 bitb_51_89 R_bl
Cb_51_88 bit_51_88 gnd C_bl
Cbb_51_88 bitb_51_88 gnd C_bl
Rb_51_89 bit_51_89 bit_51_90 R_bl
Rbb_51_89 bitb_51_89 bitb_51_90 R_bl
Cb_51_89 bit_51_89 gnd C_bl
Cbb_51_89 bitb_51_89 gnd C_bl
Rb_51_90 bit_51_90 bit_51_91 R_bl
Rbb_51_90 bitb_51_90 bitb_51_91 R_bl
Cb_51_90 bit_51_90 gnd C_bl
Cbb_51_90 bitb_51_90 gnd C_bl
Rb_51_91 bit_51_91 bit_51_92 R_bl
Rbb_51_91 bitb_51_91 bitb_51_92 R_bl
Cb_51_91 bit_51_91 gnd C_bl
Cbb_51_91 bitb_51_91 gnd C_bl
Rb_51_92 bit_51_92 bit_51_93 R_bl
Rbb_51_92 bitb_51_92 bitb_51_93 R_bl
Cb_51_92 bit_51_92 gnd C_bl
Cbb_51_92 bitb_51_92 gnd C_bl
Rb_51_93 bit_51_93 bit_51_94 R_bl
Rbb_51_93 bitb_51_93 bitb_51_94 R_bl
Cb_51_93 bit_51_93 gnd C_bl
Cbb_51_93 bitb_51_93 gnd C_bl
Rb_51_94 bit_51_94 bit_51_95 R_bl
Rbb_51_94 bitb_51_94 bitb_51_95 R_bl
Cb_51_94 bit_51_94 gnd C_bl
Cbb_51_94 bitb_51_94 gnd C_bl
Rb_51_95 bit_51_95 bit_51_96 R_bl
Rbb_51_95 bitb_51_95 bitb_51_96 R_bl
Cb_51_95 bit_51_95 gnd C_bl
Cbb_51_95 bitb_51_95 gnd C_bl
Rb_51_96 bit_51_96 bit_51_97 R_bl
Rbb_51_96 bitb_51_96 bitb_51_97 R_bl
Cb_51_96 bit_51_96 gnd C_bl
Cbb_51_96 bitb_51_96 gnd C_bl
Rb_51_97 bit_51_97 bit_51_98 R_bl
Rbb_51_97 bitb_51_97 bitb_51_98 R_bl
Cb_51_97 bit_51_97 gnd C_bl
Cbb_51_97 bitb_51_97 gnd C_bl
Rb_51_98 bit_51_98 bit_51_99 R_bl
Rbb_51_98 bitb_51_98 bitb_51_99 R_bl
Cb_51_98 bit_51_98 gnd C_bl
Cbb_51_98 bitb_51_98 gnd C_bl
Rb_51_99 bit_51_99 bit_51_100 R_bl
Rbb_51_99 bitb_51_99 bitb_51_100 R_bl
Cb_51_99 bit_51_99 gnd C_bl
Cbb_51_99 bitb_51_99 gnd C_bl
Rb_52_0 bit_52_0 bit_52_1 R_bl
Rbb_52_0 bitb_52_0 bitb_52_1 R_bl
Cb_52_0 bit_52_0 gnd C_bl
Cbb_52_0 bitb_52_0 gnd C_bl
Rb_52_1 bit_52_1 bit_52_2 R_bl
Rbb_52_1 bitb_52_1 bitb_52_2 R_bl
Cb_52_1 bit_52_1 gnd C_bl
Cbb_52_1 bitb_52_1 gnd C_bl
Rb_52_2 bit_52_2 bit_52_3 R_bl
Rbb_52_2 bitb_52_2 bitb_52_3 R_bl
Cb_52_2 bit_52_2 gnd C_bl
Cbb_52_2 bitb_52_2 gnd C_bl
Rb_52_3 bit_52_3 bit_52_4 R_bl
Rbb_52_3 bitb_52_3 bitb_52_4 R_bl
Cb_52_3 bit_52_3 gnd C_bl
Cbb_52_3 bitb_52_3 gnd C_bl
Rb_52_4 bit_52_4 bit_52_5 R_bl
Rbb_52_4 bitb_52_4 bitb_52_5 R_bl
Cb_52_4 bit_52_4 gnd C_bl
Cbb_52_4 bitb_52_4 gnd C_bl
Rb_52_5 bit_52_5 bit_52_6 R_bl
Rbb_52_5 bitb_52_5 bitb_52_6 R_bl
Cb_52_5 bit_52_5 gnd C_bl
Cbb_52_5 bitb_52_5 gnd C_bl
Rb_52_6 bit_52_6 bit_52_7 R_bl
Rbb_52_6 bitb_52_6 bitb_52_7 R_bl
Cb_52_6 bit_52_6 gnd C_bl
Cbb_52_6 bitb_52_6 gnd C_bl
Rb_52_7 bit_52_7 bit_52_8 R_bl
Rbb_52_7 bitb_52_7 bitb_52_8 R_bl
Cb_52_7 bit_52_7 gnd C_bl
Cbb_52_7 bitb_52_7 gnd C_bl
Rb_52_8 bit_52_8 bit_52_9 R_bl
Rbb_52_8 bitb_52_8 bitb_52_9 R_bl
Cb_52_8 bit_52_8 gnd C_bl
Cbb_52_8 bitb_52_8 gnd C_bl
Rb_52_9 bit_52_9 bit_52_10 R_bl
Rbb_52_9 bitb_52_9 bitb_52_10 R_bl
Cb_52_9 bit_52_9 gnd C_bl
Cbb_52_9 bitb_52_9 gnd C_bl
Rb_52_10 bit_52_10 bit_52_11 R_bl
Rbb_52_10 bitb_52_10 bitb_52_11 R_bl
Cb_52_10 bit_52_10 gnd C_bl
Cbb_52_10 bitb_52_10 gnd C_bl
Rb_52_11 bit_52_11 bit_52_12 R_bl
Rbb_52_11 bitb_52_11 bitb_52_12 R_bl
Cb_52_11 bit_52_11 gnd C_bl
Cbb_52_11 bitb_52_11 gnd C_bl
Rb_52_12 bit_52_12 bit_52_13 R_bl
Rbb_52_12 bitb_52_12 bitb_52_13 R_bl
Cb_52_12 bit_52_12 gnd C_bl
Cbb_52_12 bitb_52_12 gnd C_bl
Rb_52_13 bit_52_13 bit_52_14 R_bl
Rbb_52_13 bitb_52_13 bitb_52_14 R_bl
Cb_52_13 bit_52_13 gnd C_bl
Cbb_52_13 bitb_52_13 gnd C_bl
Rb_52_14 bit_52_14 bit_52_15 R_bl
Rbb_52_14 bitb_52_14 bitb_52_15 R_bl
Cb_52_14 bit_52_14 gnd C_bl
Cbb_52_14 bitb_52_14 gnd C_bl
Rb_52_15 bit_52_15 bit_52_16 R_bl
Rbb_52_15 bitb_52_15 bitb_52_16 R_bl
Cb_52_15 bit_52_15 gnd C_bl
Cbb_52_15 bitb_52_15 gnd C_bl
Rb_52_16 bit_52_16 bit_52_17 R_bl
Rbb_52_16 bitb_52_16 bitb_52_17 R_bl
Cb_52_16 bit_52_16 gnd C_bl
Cbb_52_16 bitb_52_16 gnd C_bl
Rb_52_17 bit_52_17 bit_52_18 R_bl
Rbb_52_17 bitb_52_17 bitb_52_18 R_bl
Cb_52_17 bit_52_17 gnd C_bl
Cbb_52_17 bitb_52_17 gnd C_bl
Rb_52_18 bit_52_18 bit_52_19 R_bl
Rbb_52_18 bitb_52_18 bitb_52_19 R_bl
Cb_52_18 bit_52_18 gnd C_bl
Cbb_52_18 bitb_52_18 gnd C_bl
Rb_52_19 bit_52_19 bit_52_20 R_bl
Rbb_52_19 bitb_52_19 bitb_52_20 R_bl
Cb_52_19 bit_52_19 gnd C_bl
Cbb_52_19 bitb_52_19 gnd C_bl
Rb_52_20 bit_52_20 bit_52_21 R_bl
Rbb_52_20 bitb_52_20 bitb_52_21 R_bl
Cb_52_20 bit_52_20 gnd C_bl
Cbb_52_20 bitb_52_20 gnd C_bl
Rb_52_21 bit_52_21 bit_52_22 R_bl
Rbb_52_21 bitb_52_21 bitb_52_22 R_bl
Cb_52_21 bit_52_21 gnd C_bl
Cbb_52_21 bitb_52_21 gnd C_bl
Rb_52_22 bit_52_22 bit_52_23 R_bl
Rbb_52_22 bitb_52_22 bitb_52_23 R_bl
Cb_52_22 bit_52_22 gnd C_bl
Cbb_52_22 bitb_52_22 gnd C_bl
Rb_52_23 bit_52_23 bit_52_24 R_bl
Rbb_52_23 bitb_52_23 bitb_52_24 R_bl
Cb_52_23 bit_52_23 gnd C_bl
Cbb_52_23 bitb_52_23 gnd C_bl
Rb_52_24 bit_52_24 bit_52_25 R_bl
Rbb_52_24 bitb_52_24 bitb_52_25 R_bl
Cb_52_24 bit_52_24 gnd C_bl
Cbb_52_24 bitb_52_24 gnd C_bl
Rb_52_25 bit_52_25 bit_52_26 R_bl
Rbb_52_25 bitb_52_25 bitb_52_26 R_bl
Cb_52_25 bit_52_25 gnd C_bl
Cbb_52_25 bitb_52_25 gnd C_bl
Rb_52_26 bit_52_26 bit_52_27 R_bl
Rbb_52_26 bitb_52_26 bitb_52_27 R_bl
Cb_52_26 bit_52_26 gnd C_bl
Cbb_52_26 bitb_52_26 gnd C_bl
Rb_52_27 bit_52_27 bit_52_28 R_bl
Rbb_52_27 bitb_52_27 bitb_52_28 R_bl
Cb_52_27 bit_52_27 gnd C_bl
Cbb_52_27 bitb_52_27 gnd C_bl
Rb_52_28 bit_52_28 bit_52_29 R_bl
Rbb_52_28 bitb_52_28 bitb_52_29 R_bl
Cb_52_28 bit_52_28 gnd C_bl
Cbb_52_28 bitb_52_28 gnd C_bl
Rb_52_29 bit_52_29 bit_52_30 R_bl
Rbb_52_29 bitb_52_29 bitb_52_30 R_bl
Cb_52_29 bit_52_29 gnd C_bl
Cbb_52_29 bitb_52_29 gnd C_bl
Rb_52_30 bit_52_30 bit_52_31 R_bl
Rbb_52_30 bitb_52_30 bitb_52_31 R_bl
Cb_52_30 bit_52_30 gnd C_bl
Cbb_52_30 bitb_52_30 gnd C_bl
Rb_52_31 bit_52_31 bit_52_32 R_bl
Rbb_52_31 bitb_52_31 bitb_52_32 R_bl
Cb_52_31 bit_52_31 gnd C_bl
Cbb_52_31 bitb_52_31 gnd C_bl
Rb_52_32 bit_52_32 bit_52_33 R_bl
Rbb_52_32 bitb_52_32 bitb_52_33 R_bl
Cb_52_32 bit_52_32 gnd C_bl
Cbb_52_32 bitb_52_32 gnd C_bl
Rb_52_33 bit_52_33 bit_52_34 R_bl
Rbb_52_33 bitb_52_33 bitb_52_34 R_bl
Cb_52_33 bit_52_33 gnd C_bl
Cbb_52_33 bitb_52_33 gnd C_bl
Rb_52_34 bit_52_34 bit_52_35 R_bl
Rbb_52_34 bitb_52_34 bitb_52_35 R_bl
Cb_52_34 bit_52_34 gnd C_bl
Cbb_52_34 bitb_52_34 gnd C_bl
Rb_52_35 bit_52_35 bit_52_36 R_bl
Rbb_52_35 bitb_52_35 bitb_52_36 R_bl
Cb_52_35 bit_52_35 gnd C_bl
Cbb_52_35 bitb_52_35 gnd C_bl
Rb_52_36 bit_52_36 bit_52_37 R_bl
Rbb_52_36 bitb_52_36 bitb_52_37 R_bl
Cb_52_36 bit_52_36 gnd C_bl
Cbb_52_36 bitb_52_36 gnd C_bl
Rb_52_37 bit_52_37 bit_52_38 R_bl
Rbb_52_37 bitb_52_37 bitb_52_38 R_bl
Cb_52_37 bit_52_37 gnd C_bl
Cbb_52_37 bitb_52_37 gnd C_bl
Rb_52_38 bit_52_38 bit_52_39 R_bl
Rbb_52_38 bitb_52_38 bitb_52_39 R_bl
Cb_52_38 bit_52_38 gnd C_bl
Cbb_52_38 bitb_52_38 gnd C_bl
Rb_52_39 bit_52_39 bit_52_40 R_bl
Rbb_52_39 bitb_52_39 bitb_52_40 R_bl
Cb_52_39 bit_52_39 gnd C_bl
Cbb_52_39 bitb_52_39 gnd C_bl
Rb_52_40 bit_52_40 bit_52_41 R_bl
Rbb_52_40 bitb_52_40 bitb_52_41 R_bl
Cb_52_40 bit_52_40 gnd C_bl
Cbb_52_40 bitb_52_40 gnd C_bl
Rb_52_41 bit_52_41 bit_52_42 R_bl
Rbb_52_41 bitb_52_41 bitb_52_42 R_bl
Cb_52_41 bit_52_41 gnd C_bl
Cbb_52_41 bitb_52_41 gnd C_bl
Rb_52_42 bit_52_42 bit_52_43 R_bl
Rbb_52_42 bitb_52_42 bitb_52_43 R_bl
Cb_52_42 bit_52_42 gnd C_bl
Cbb_52_42 bitb_52_42 gnd C_bl
Rb_52_43 bit_52_43 bit_52_44 R_bl
Rbb_52_43 bitb_52_43 bitb_52_44 R_bl
Cb_52_43 bit_52_43 gnd C_bl
Cbb_52_43 bitb_52_43 gnd C_bl
Rb_52_44 bit_52_44 bit_52_45 R_bl
Rbb_52_44 bitb_52_44 bitb_52_45 R_bl
Cb_52_44 bit_52_44 gnd C_bl
Cbb_52_44 bitb_52_44 gnd C_bl
Rb_52_45 bit_52_45 bit_52_46 R_bl
Rbb_52_45 bitb_52_45 bitb_52_46 R_bl
Cb_52_45 bit_52_45 gnd C_bl
Cbb_52_45 bitb_52_45 gnd C_bl
Rb_52_46 bit_52_46 bit_52_47 R_bl
Rbb_52_46 bitb_52_46 bitb_52_47 R_bl
Cb_52_46 bit_52_46 gnd C_bl
Cbb_52_46 bitb_52_46 gnd C_bl
Rb_52_47 bit_52_47 bit_52_48 R_bl
Rbb_52_47 bitb_52_47 bitb_52_48 R_bl
Cb_52_47 bit_52_47 gnd C_bl
Cbb_52_47 bitb_52_47 gnd C_bl
Rb_52_48 bit_52_48 bit_52_49 R_bl
Rbb_52_48 bitb_52_48 bitb_52_49 R_bl
Cb_52_48 bit_52_48 gnd C_bl
Cbb_52_48 bitb_52_48 gnd C_bl
Rb_52_49 bit_52_49 bit_52_50 R_bl
Rbb_52_49 bitb_52_49 bitb_52_50 R_bl
Cb_52_49 bit_52_49 gnd C_bl
Cbb_52_49 bitb_52_49 gnd C_bl
Rb_52_50 bit_52_50 bit_52_51 R_bl
Rbb_52_50 bitb_52_50 bitb_52_51 R_bl
Cb_52_50 bit_52_50 gnd C_bl
Cbb_52_50 bitb_52_50 gnd C_bl
Rb_52_51 bit_52_51 bit_52_52 R_bl
Rbb_52_51 bitb_52_51 bitb_52_52 R_bl
Cb_52_51 bit_52_51 gnd C_bl
Cbb_52_51 bitb_52_51 gnd C_bl
Rb_52_52 bit_52_52 bit_52_53 R_bl
Rbb_52_52 bitb_52_52 bitb_52_53 R_bl
Cb_52_52 bit_52_52 gnd C_bl
Cbb_52_52 bitb_52_52 gnd C_bl
Rb_52_53 bit_52_53 bit_52_54 R_bl
Rbb_52_53 bitb_52_53 bitb_52_54 R_bl
Cb_52_53 bit_52_53 gnd C_bl
Cbb_52_53 bitb_52_53 gnd C_bl
Rb_52_54 bit_52_54 bit_52_55 R_bl
Rbb_52_54 bitb_52_54 bitb_52_55 R_bl
Cb_52_54 bit_52_54 gnd C_bl
Cbb_52_54 bitb_52_54 gnd C_bl
Rb_52_55 bit_52_55 bit_52_56 R_bl
Rbb_52_55 bitb_52_55 bitb_52_56 R_bl
Cb_52_55 bit_52_55 gnd C_bl
Cbb_52_55 bitb_52_55 gnd C_bl
Rb_52_56 bit_52_56 bit_52_57 R_bl
Rbb_52_56 bitb_52_56 bitb_52_57 R_bl
Cb_52_56 bit_52_56 gnd C_bl
Cbb_52_56 bitb_52_56 gnd C_bl
Rb_52_57 bit_52_57 bit_52_58 R_bl
Rbb_52_57 bitb_52_57 bitb_52_58 R_bl
Cb_52_57 bit_52_57 gnd C_bl
Cbb_52_57 bitb_52_57 gnd C_bl
Rb_52_58 bit_52_58 bit_52_59 R_bl
Rbb_52_58 bitb_52_58 bitb_52_59 R_bl
Cb_52_58 bit_52_58 gnd C_bl
Cbb_52_58 bitb_52_58 gnd C_bl
Rb_52_59 bit_52_59 bit_52_60 R_bl
Rbb_52_59 bitb_52_59 bitb_52_60 R_bl
Cb_52_59 bit_52_59 gnd C_bl
Cbb_52_59 bitb_52_59 gnd C_bl
Rb_52_60 bit_52_60 bit_52_61 R_bl
Rbb_52_60 bitb_52_60 bitb_52_61 R_bl
Cb_52_60 bit_52_60 gnd C_bl
Cbb_52_60 bitb_52_60 gnd C_bl
Rb_52_61 bit_52_61 bit_52_62 R_bl
Rbb_52_61 bitb_52_61 bitb_52_62 R_bl
Cb_52_61 bit_52_61 gnd C_bl
Cbb_52_61 bitb_52_61 gnd C_bl
Rb_52_62 bit_52_62 bit_52_63 R_bl
Rbb_52_62 bitb_52_62 bitb_52_63 R_bl
Cb_52_62 bit_52_62 gnd C_bl
Cbb_52_62 bitb_52_62 gnd C_bl
Rb_52_63 bit_52_63 bit_52_64 R_bl
Rbb_52_63 bitb_52_63 bitb_52_64 R_bl
Cb_52_63 bit_52_63 gnd C_bl
Cbb_52_63 bitb_52_63 gnd C_bl
Rb_52_64 bit_52_64 bit_52_65 R_bl
Rbb_52_64 bitb_52_64 bitb_52_65 R_bl
Cb_52_64 bit_52_64 gnd C_bl
Cbb_52_64 bitb_52_64 gnd C_bl
Rb_52_65 bit_52_65 bit_52_66 R_bl
Rbb_52_65 bitb_52_65 bitb_52_66 R_bl
Cb_52_65 bit_52_65 gnd C_bl
Cbb_52_65 bitb_52_65 gnd C_bl
Rb_52_66 bit_52_66 bit_52_67 R_bl
Rbb_52_66 bitb_52_66 bitb_52_67 R_bl
Cb_52_66 bit_52_66 gnd C_bl
Cbb_52_66 bitb_52_66 gnd C_bl
Rb_52_67 bit_52_67 bit_52_68 R_bl
Rbb_52_67 bitb_52_67 bitb_52_68 R_bl
Cb_52_67 bit_52_67 gnd C_bl
Cbb_52_67 bitb_52_67 gnd C_bl
Rb_52_68 bit_52_68 bit_52_69 R_bl
Rbb_52_68 bitb_52_68 bitb_52_69 R_bl
Cb_52_68 bit_52_68 gnd C_bl
Cbb_52_68 bitb_52_68 gnd C_bl
Rb_52_69 bit_52_69 bit_52_70 R_bl
Rbb_52_69 bitb_52_69 bitb_52_70 R_bl
Cb_52_69 bit_52_69 gnd C_bl
Cbb_52_69 bitb_52_69 gnd C_bl
Rb_52_70 bit_52_70 bit_52_71 R_bl
Rbb_52_70 bitb_52_70 bitb_52_71 R_bl
Cb_52_70 bit_52_70 gnd C_bl
Cbb_52_70 bitb_52_70 gnd C_bl
Rb_52_71 bit_52_71 bit_52_72 R_bl
Rbb_52_71 bitb_52_71 bitb_52_72 R_bl
Cb_52_71 bit_52_71 gnd C_bl
Cbb_52_71 bitb_52_71 gnd C_bl
Rb_52_72 bit_52_72 bit_52_73 R_bl
Rbb_52_72 bitb_52_72 bitb_52_73 R_bl
Cb_52_72 bit_52_72 gnd C_bl
Cbb_52_72 bitb_52_72 gnd C_bl
Rb_52_73 bit_52_73 bit_52_74 R_bl
Rbb_52_73 bitb_52_73 bitb_52_74 R_bl
Cb_52_73 bit_52_73 gnd C_bl
Cbb_52_73 bitb_52_73 gnd C_bl
Rb_52_74 bit_52_74 bit_52_75 R_bl
Rbb_52_74 bitb_52_74 bitb_52_75 R_bl
Cb_52_74 bit_52_74 gnd C_bl
Cbb_52_74 bitb_52_74 gnd C_bl
Rb_52_75 bit_52_75 bit_52_76 R_bl
Rbb_52_75 bitb_52_75 bitb_52_76 R_bl
Cb_52_75 bit_52_75 gnd C_bl
Cbb_52_75 bitb_52_75 gnd C_bl
Rb_52_76 bit_52_76 bit_52_77 R_bl
Rbb_52_76 bitb_52_76 bitb_52_77 R_bl
Cb_52_76 bit_52_76 gnd C_bl
Cbb_52_76 bitb_52_76 gnd C_bl
Rb_52_77 bit_52_77 bit_52_78 R_bl
Rbb_52_77 bitb_52_77 bitb_52_78 R_bl
Cb_52_77 bit_52_77 gnd C_bl
Cbb_52_77 bitb_52_77 gnd C_bl
Rb_52_78 bit_52_78 bit_52_79 R_bl
Rbb_52_78 bitb_52_78 bitb_52_79 R_bl
Cb_52_78 bit_52_78 gnd C_bl
Cbb_52_78 bitb_52_78 gnd C_bl
Rb_52_79 bit_52_79 bit_52_80 R_bl
Rbb_52_79 bitb_52_79 bitb_52_80 R_bl
Cb_52_79 bit_52_79 gnd C_bl
Cbb_52_79 bitb_52_79 gnd C_bl
Rb_52_80 bit_52_80 bit_52_81 R_bl
Rbb_52_80 bitb_52_80 bitb_52_81 R_bl
Cb_52_80 bit_52_80 gnd C_bl
Cbb_52_80 bitb_52_80 gnd C_bl
Rb_52_81 bit_52_81 bit_52_82 R_bl
Rbb_52_81 bitb_52_81 bitb_52_82 R_bl
Cb_52_81 bit_52_81 gnd C_bl
Cbb_52_81 bitb_52_81 gnd C_bl
Rb_52_82 bit_52_82 bit_52_83 R_bl
Rbb_52_82 bitb_52_82 bitb_52_83 R_bl
Cb_52_82 bit_52_82 gnd C_bl
Cbb_52_82 bitb_52_82 gnd C_bl
Rb_52_83 bit_52_83 bit_52_84 R_bl
Rbb_52_83 bitb_52_83 bitb_52_84 R_bl
Cb_52_83 bit_52_83 gnd C_bl
Cbb_52_83 bitb_52_83 gnd C_bl
Rb_52_84 bit_52_84 bit_52_85 R_bl
Rbb_52_84 bitb_52_84 bitb_52_85 R_bl
Cb_52_84 bit_52_84 gnd C_bl
Cbb_52_84 bitb_52_84 gnd C_bl
Rb_52_85 bit_52_85 bit_52_86 R_bl
Rbb_52_85 bitb_52_85 bitb_52_86 R_bl
Cb_52_85 bit_52_85 gnd C_bl
Cbb_52_85 bitb_52_85 gnd C_bl
Rb_52_86 bit_52_86 bit_52_87 R_bl
Rbb_52_86 bitb_52_86 bitb_52_87 R_bl
Cb_52_86 bit_52_86 gnd C_bl
Cbb_52_86 bitb_52_86 gnd C_bl
Rb_52_87 bit_52_87 bit_52_88 R_bl
Rbb_52_87 bitb_52_87 bitb_52_88 R_bl
Cb_52_87 bit_52_87 gnd C_bl
Cbb_52_87 bitb_52_87 gnd C_bl
Rb_52_88 bit_52_88 bit_52_89 R_bl
Rbb_52_88 bitb_52_88 bitb_52_89 R_bl
Cb_52_88 bit_52_88 gnd C_bl
Cbb_52_88 bitb_52_88 gnd C_bl
Rb_52_89 bit_52_89 bit_52_90 R_bl
Rbb_52_89 bitb_52_89 bitb_52_90 R_bl
Cb_52_89 bit_52_89 gnd C_bl
Cbb_52_89 bitb_52_89 gnd C_bl
Rb_52_90 bit_52_90 bit_52_91 R_bl
Rbb_52_90 bitb_52_90 bitb_52_91 R_bl
Cb_52_90 bit_52_90 gnd C_bl
Cbb_52_90 bitb_52_90 gnd C_bl
Rb_52_91 bit_52_91 bit_52_92 R_bl
Rbb_52_91 bitb_52_91 bitb_52_92 R_bl
Cb_52_91 bit_52_91 gnd C_bl
Cbb_52_91 bitb_52_91 gnd C_bl
Rb_52_92 bit_52_92 bit_52_93 R_bl
Rbb_52_92 bitb_52_92 bitb_52_93 R_bl
Cb_52_92 bit_52_92 gnd C_bl
Cbb_52_92 bitb_52_92 gnd C_bl
Rb_52_93 bit_52_93 bit_52_94 R_bl
Rbb_52_93 bitb_52_93 bitb_52_94 R_bl
Cb_52_93 bit_52_93 gnd C_bl
Cbb_52_93 bitb_52_93 gnd C_bl
Rb_52_94 bit_52_94 bit_52_95 R_bl
Rbb_52_94 bitb_52_94 bitb_52_95 R_bl
Cb_52_94 bit_52_94 gnd C_bl
Cbb_52_94 bitb_52_94 gnd C_bl
Rb_52_95 bit_52_95 bit_52_96 R_bl
Rbb_52_95 bitb_52_95 bitb_52_96 R_bl
Cb_52_95 bit_52_95 gnd C_bl
Cbb_52_95 bitb_52_95 gnd C_bl
Rb_52_96 bit_52_96 bit_52_97 R_bl
Rbb_52_96 bitb_52_96 bitb_52_97 R_bl
Cb_52_96 bit_52_96 gnd C_bl
Cbb_52_96 bitb_52_96 gnd C_bl
Rb_52_97 bit_52_97 bit_52_98 R_bl
Rbb_52_97 bitb_52_97 bitb_52_98 R_bl
Cb_52_97 bit_52_97 gnd C_bl
Cbb_52_97 bitb_52_97 gnd C_bl
Rb_52_98 bit_52_98 bit_52_99 R_bl
Rbb_52_98 bitb_52_98 bitb_52_99 R_bl
Cb_52_98 bit_52_98 gnd C_bl
Cbb_52_98 bitb_52_98 gnd C_bl
Rb_52_99 bit_52_99 bit_52_100 R_bl
Rbb_52_99 bitb_52_99 bitb_52_100 R_bl
Cb_52_99 bit_52_99 gnd C_bl
Cbb_52_99 bitb_52_99 gnd C_bl
Rb_53_0 bit_53_0 bit_53_1 R_bl
Rbb_53_0 bitb_53_0 bitb_53_1 R_bl
Cb_53_0 bit_53_0 gnd C_bl
Cbb_53_0 bitb_53_0 gnd C_bl
Rb_53_1 bit_53_1 bit_53_2 R_bl
Rbb_53_1 bitb_53_1 bitb_53_2 R_bl
Cb_53_1 bit_53_1 gnd C_bl
Cbb_53_1 bitb_53_1 gnd C_bl
Rb_53_2 bit_53_2 bit_53_3 R_bl
Rbb_53_2 bitb_53_2 bitb_53_3 R_bl
Cb_53_2 bit_53_2 gnd C_bl
Cbb_53_2 bitb_53_2 gnd C_bl
Rb_53_3 bit_53_3 bit_53_4 R_bl
Rbb_53_3 bitb_53_3 bitb_53_4 R_bl
Cb_53_3 bit_53_3 gnd C_bl
Cbb_53_3 bitb_53_3 gnd C_bl
Rb_53_4 bit_53_4 bit_53_5 R_bl
Rbb_53_4 bitb_53_4 bitb_53_5 R_bl
Cb_53_4 bit_53_4 gnd C_bl
Cbb_53_4 bitb_53_4 gnd C_bl
Rb_53_5 bit_53_5 bit_53_6 R_bl
Rbb_53_5 bitb_53_5 bitb_53_6 R_bl
Cb_53_5 bit_53_5 gnd C_bl
Cbb_53_5 bitb_53_5 gnd C_bl
Rb_53_6 bit_53_6 bit_53_7 R_bl
Rbb_53_6 bitb_53_6 bitb_53_7 R_bl
Cb_53_6 bit_53_6 gnd C_bl
Cbb_53_6 bitb_53_6 gnd C_bl
Rb_53_7 bit_53_7 bit_53_8 R_bl
Rbb_53_7 bitb_53_7 bitb_53_8 R_bl
Cb_53_7 bit_53_7 gnd C_bl
Cbb_53_7 bitb_53_7 gnd C_bl
Rb_53_8 bit_53_8 bit_53_9 R_bl
Rbb_53_8 bitb_53_8 bitb_53_9 R_bl
Cb_53_8 bit_53_8 gnd C_bl
Cbb_53_8 bitb_53_8 gnd C_bl
Rb_53_9 bit_53_9 bit_53_10 R_bl
Rbb_53_9 bitb_53_9 bitb_53_10 R_bl
Cb_53_9 bit_53_9 gnd C_bl
Cbb_53_9 bitb_53_9 gnd C_bl
Rb_53_10 bit_53_10 bit_53_11 R_bl
Rbb_53_10 bitb_53_10 bitb_53_11 R_bl
Cb_53_10 bit_53_10 gnd C_bl
Cbb_53_10 bitb_53_10 gnd C_bl
Rb_53_11 bit_53_11 bit_53_12 R_bl
Rbb_53_11 bitb_53_11 bitb_53_12 R_bl
Cb_53_11 bit_53_11 gnd C_bl
Cbb_53_11 bitb_53_11 gnd C_bl
Rb_53_12 bit_53_12 bit_53_13 R_bl
Rbb_53_12 bitb_53_12 bitb_53_13 R_bl
Cb_53_12 bit_53_12 gnd C_bl
Cbb_53_12 bitb_53_12 gnd C_bl
Rb_53_13 bit_53_13 bit_53_14 R_bl
Rbb_53_13 bitb_53_13 bitb_53_14 R_bl
Cb_53_13 bit_53_13 gnd C_bl
Cbb_53_13 bitb_53_13 gnd C_bl
Rb_53_14 bit_53_14 bit_53_15 R_bl
Rbb_53_14 bitb_53_14 bitb_53_15 R_bl
Cb_53_14 bit_53_14 gnd C_bl
Cbb_53_14 bitb_53_14 gnd C_bl
Rb_53_15 bit_53_15 bit_53_16 R_bl
Rbb_53_15 bitb_53_15 bitb_53_16 R_bl
Cb_53_15 bit_53_15 gnd C_bl
Cbb_53_15 bitb_53_15 gnd C_bl
Rb_53_16 bit_53_16 bit_53_17 R_bl
Rbb_53_16 bitb_53_16 bitb_53_17 R_bl
Cb_53_16 bit_53_16 gnd C_bl
Cbb_53_16 bitb_53_16 gnd C_bl
Rb_53_17 bit_53_17 bit_53_18 R_bl
Rbb_53_17 bitb_53_17 bitb_53_18 R_bl
Cb_53_17 bit_53_17 gnd C_bl
Cbb_53_17 bitb_53_17 gnd C_bl
Rb_53_18 bit_53_18 bit_53_19 R_bl
Rbb_53_18 bitb_53_18 bitb_53_19 R_bl
Cb_53_18 bit_53_18 gnd C_bl
Cbb_53_18 bitb_53_18 gnd C_bl
Rb_53_19 bit_53_19 bit_53_20 R_bl
Rbb_53_19 bitb_53_19 bitb_53_20 R_bl
Cb_53_19 bit_53_19 gnd C_bl
Cbb_53_19 bitb_53_19 gnd C_bl
Rb_53_20 bit_53_20 bit_53_21 R_bl
Rbb_53_20 bitb_53_20 bitb_53_21 R_bl
Cb_53_20 bit_53_20 gnd C_bl
Cbb_53_20 bitb_53_20 gnd C_bl
Rb_53_21 bit_53_21 bit_53_22 R_bl
Rbb_53_21 bitb_53_21 bitb_53_22 R_bl
Cb_53_21 bit_53_21 gnd C_bl
Cbb_53_21 bitb_53_21 gnd C_bl
Rb_53_22 bit_53_22 bit_53_23 R_bl
Rbb_53_22 bitb_53_22 bitb_53_23 R_bl
Cb_53_22 bit_53_22 gnd C_bl
Cbb_53_22 bitb_53_22 gnd C_bl
Rb_53_23 bit_53_23 bit_53_24 R_bl
Rbb_53_23 bitb_53_23 bitb_53_24 R_bl
Cb_53_23 bit_53_23 gnd C_bl
Cbb_53_23 bitb_53_23 gnd C_bl
Rb_53_24 bit_53_24 bit_53_25 R_bl
Rbb_53_24 bitb_53_24 bitb_53_25 R_bl
Cb_53_24 bit_53_24 gnd C_bl
Cbb_53_24 bitb_53_24 gnd C_bl
Rb_53_25 bit_53_25 bit_53_26 R_bl
Rbb_53_25 bitb_53_25 bitb_53_26 R_bl
Cb_53_25 bit_53_25 gnd C_bl
Cbb_53_25 bitb_53_25 gnd C_bl
Rb_53_26 bit_53_26 bit_53_27 R_bl
Rbb_53_26 bitb_53_26 bitb_53_27 R_bl
Cb_53_26 bit_53_26 gnd C_bl
Cbb_53_26 bitb_53_26 gnd C_bl
Rb_53_27 bit_53_27 bit_53_28 R_bl
Rbb_53_27 bitb_53_27 bitb_53_28 R_bl
Cb_53_27 bit_53_27 gnd C_bl
Cbb_53_27 bitb_53_27 gnd C_bl
Rb_53_28 bit_53_28 bit_53_29 R_bl
Rbb_53_28 bitb_53_28 bitb_53_29 R_bl
Cb_53_28 bit_53_28 gnd C_bl
Cbb_53_28 bitb_53_28 gnd C_bl
Rb_53_29 bit_53_29 bit_53_30 R_bl
Rbb_53_29 bitb_53_29 bitb_53_30 R_bl
Cb_53_29 bit_53_29 gnd C_bl
Cbb_53_29 bitb_53_29 gnd C_bl
Rb_53_30 bit_53_30 bit_53_31 R_bl
Rbb_53_30 bitb_53_30 bitb_53_31 R_bl
Cb_53_30 bit_53_30 gnd C_bl
Cbb_53_30 bitb_53_30 gnd C_bl
Rb_53_31 bit_53_31 bit_53_32 R_bl
Rbb_53_31 bitb_53_31 bitb_53_32 R_bl
Cb_53_31 bit_53_31 gnd C_bl
Cbb_53_31 bitb_53_31 gnd C_bl
Rb_53_32 bit_53_32 bit_53_33 R_bl
Rbb_53_32 bitb_53_32 bitb_53_33 R_bl
Cb_53_32 bit_53_32 gnd C_bl
Cbb_53_32 bitb_53_32 gnd C_bl
Rb_53_33 bit_53_33 bit_53_34 R_bl
Rbb_53_33 bitb_53_33 bitb_53_34 R_bl
Cb_53_33 bit_53_33 gnd C_bl
Cbb_53_33 bitb_53_33 gnd C_bl
Rb_53_34 bit_53_34 bit_53_35 R_bl
Rbb_53_34 bitb_53_34 bitb_53_35 R_bl
Cb_53_34 bit_53_34 gnd C_bl
Cbb_53_34 bitb_53_34 gnd C_bl
Rb_53_35 bit_53_35 bit_53_36 R_bl
Rbb_53_35 bitb_53_35 bitb_53_36 R_bl
Cb_53_35 bit_53_35 gnd C_bl
Cbb_53_35 bitb_53_35 gnd C_bl
Rb_53_36 bit_53_36 bit_53_37 R_bl
Rbb_53_36 bitb_53_36 bitb_53_37 R_bl
Cb_53_36 bit_53_36 gnd C_bl
Cbb_53_36 bitb_53_36 gnd C_bl
Rb_53_37 bit_53_37 bit_53_38 R_bl
Rbb_53_37 bitb_53_37 bitb_53_38 R_bl
Cb_53_37 bit_53_37 gnd C_bl
Cbb_53_37 bitb_53_37 gnd C_bl
Rb_53_38 bit_53_38 bit_53_39 R_bl
Rbb_53_38 bitb_53_38 bitb_53_39 R_bl
Cb_53_38 bit_53_38 gnd C_bl
Cbb_53_38 bitb_53_38 gnd C_bl
Rb_53_39 bit_53_39 bit_53_40 R_bl
Rbb_53_39 bitb_53_39 bitb_53_40 R_bl
Cb_53_39 bit_53_39 gnd C_bl
Cbb_53_39 bitb_53_39 gnd C_bl
Rb_53_40 bit_53_40 bit_53_41 R_bl
Rbb_53_40 bitb_53_40 bitb_53_41 R_bl
Cb_53_40 bit_53_40 gnd C_bl
Cbb_53_40 bitb_53_40 gnd C_bl
Rb_53_41 bit_53_41 bit_53_42 R_bl
Rbb_53_41 bitb_53_41 bitb_53_42 R_bl
Cb_53_41 bit_53_41 gnd C_bl
Cbb_53_41 bitb_53_41 gnd C_bl
Rb_53_42 bit_53_42 bit_53_43 R_bl
Rbb_53_42 bitb_53_42 bitb_53_43 R_bl
Cb_53_42 bit_53_42 gnd C_bl
Cbb_53_42 bitb_53_42 gnd C_bl
Rb_53_43 bit_53_43 bit_53_44 R_bl
Rbb_53_43 bitb_53_43 bitb_53_44 R_bl
Cb_53_43 bit_53_43 gnd C_bl
Cbb_53_43 bitb_53_43 gnd C_bl
Rb_53_44 bit_53_44 bit_53_45 R_bl
Rbb_53_44 bitb_53_44 bitb_53_45 R_bl
Cb_53_44 bit_53_44 gnd C_bl
Cbb_53_44 bitb_53_44 gnd C_bl
Rb_53_45 bit_53_45 bit_53_46 R_bl
Rbb_53_45 bitb_53_45 bitb_53_46 R_bl
Cb_53_45 bit_53_45 gnd C_bl
Cbb_53_45 bitb_53_45 gnd C_bl
Rb_53_46 bit_53_46 bit_53_47 R_bl
Rbb_53_46 bitb_53_46 bitb_53_47 R_bl
Cb_53_46 bit_53_46 gnd C_bl
Cbb_53_46 bitb_53_46 gnd C_bl
Rb_53_47 bit_53_47 bit_53_48 R_bl
Rbb_53_47 bitb_53_47 bitb_53_48 R_bl
Cb_53_47 bit_53_47 gnd C_bl
Cbb_53_47 bitb_53_47 gnd C_bl
Rb_53_48 bit_53_48 bit_53_49 R_bl
Rbb_53_48 bitb_53_48 bitb_53_49 R_bl
Cb_53_48 bit_53_48 gnd C_bl
Cbb_53_48 bitb_53_48 gnd C_bl
Rb_53_49 bit_53_49 bit_53_50 R_bl
Rbb_53_49 bitb_53_49 bitb_53_50 R_bl
Cb_53_49 bit_53_49 gnd C_bl
Cbb_53_49 bitb_53_49 gnd C_bl
Rb_53_50 bit_53_50 bit_53_51 R_bl
Rbb_53_50 bitb_53_50 bitb_53_51 R_bl
Cb_53_50 bit_53_50 gnd C_bl
Cbb_53_50 bitb_53_50 gnd C_bl
Rb_53_51 bit_53_51 bit_53_52 R_bl
Rbb_53_51 bitb_53_51 bitb_53_52 R_bl
Cb_53_51 bit_53_51 gnd C_bl
Cbb_53_51 bitb_53_51 gnd C_bl
Rb_53_52 bit_53_52 bit_53_53 R_bl
Rbb_53_52 bitb_53_52 bitb_53_53 R_bl
Cb_53_52 bit_53_52 gnd C_bl
Cbb_53_52 bitb_53_52 gnd C_bl
Rb_53_53 bit_53_53 bit_53_54 R_bl
Rbb_53_53 bitb_53_53 bitb_53_54 R_bl
Cb_53_53 bit_53_53 gnd C_bl
Cbb_53_53 bitb_53_53 gnd C_bl
Rb_53_54 bit_53_54 bit_53_55 R_bl
Rbb_53_54 bitb_53_54 bitb_53_55 R_bl
Cb_53_54 bit_53_54 gnd C_bl
Cbb_53_54 bitb_53_54 gnd C_bl
Rb_53_55 bit_53_55 bit_53_56 R_bl
Rbb_53_55 bitb_53_55 bitb_53_56 R_bl
Cb_53_55 bit_53_55 gnd C_bl
Cbb_53_55 bitb_53_55 gnd C_bl
Rb_53_56 bit_53_56 bit_53_57 R_bl
Rbb_53_56 bitb_53_56 bitb_53_57 R_bl
Cb_53_56 bit_53_56 gnd C_bl
Cbb_53_56 bitb_53_56 gnd C_bl
Rb_53_57 bit_53_57 bit_53_58 R_bl
Rbb_53_57 bitb_53_57 bitb_53_58 R_bl
Cb_53_57 bit_53_57 gnd C_bl
Cbb_53_57 bitb_53_57 gnd C_bl
Rb_53_58 bit_53_58 bit_53_59 R_bl
Rbb_53_58 bitb_53_58 bitb_53_59 R_bl
Cb_53_58 bit_53_58 gnd C_bl
Cbb_53_58 bitb_53_58 gnd C_bl
Rb_53_59 bit_53_59 bit_53_60 R_bl
Rbb_53_59 bitb_53_59 bitb_53_60 R_bl
Cb_53_59 bit_53_59 gnd C_bl
Cbb_53_59 bitb_53_59 gnd C_bl
Rb_53_60 bit_53_60 bit_53_61 R_bl
Rbb_53_60 bitb_53_60 bitb_53_61 R_bl
Cb_53_60 bit_53_60 gnd C_bl
Cbb_53_60 bitb_53_60 gnd C_bl
Rb_53_61 bit_53_61 bit_53_62 R_bl
Rbb_53_61 bitb_53_61 bitb_53_62 R_bl
Cb_53_61 bit_53_61 gnd C_bl
Cbb_53_61 bitb_53_61 gnd C_bl
Rb_53_62 bit_53_62 bit_53_63 R_bl
Rbb_53_62 bitb_53_62 bitb_53_63 R_bl
Cb_53_62 bit_53_62 gnd C_bl
Cbb_53_62 bitb_53_62 gnd C_bl
Rb_53_63 bit_53_63 bit_53_64 R_bl
Rbb_53_63 bitb_53_63 bitb_53_64 R_bl
Cb_53_63 bit_53_63 gnd C_bl
Cbb_53_63 bitb_53_63 gnd C_bl
Rb_53_64 bit_53_64 bit_53_65 R_bl
Rbb_53_64 bitb_53_64 bitb_53_65 R_bl
Cb_53_64 bit_53_64 gnd C_bl
Cbb_53_64 bitb_53_64 gnd C_bl
Rb_53_65 bit_53_65 bit_53_66 R_bl
Rbb_53_65 bitb_53_65 bitb_53_66 R_bl
Cb_53_65 bit_53_65 gnd C_bl
Cbb_53_65 bitb_53_65 gnd C_bl
Rb_53_66 bit_53_66 bit_53_67 R_bl
Rbb_53_66 bitb_53_66 bitb_53_67 R_bl
Cb_53_66 bit_53_66 gnd C_bl
Cbb_53_66 bitb_53_66 gnd C_bl
Rb_53_67 bit_53_67 bit_53_68 R_bl
Rbb_53_67 bitb_53_67 bitb_53_68 R_bl
Cb_53_67 bit_53_67 gnd C_bl
Cbb_53_67 bitb_53_67 gnd C_bl
Rb_53_68 bit_53_68 bit_53_69 R_bl
Rbb_53_68 bitb_53_68 bitb_53_69 R_bl
Cb_53_68 bit_53_68 gnd C_bl
Cbb_53_68 bitb_53_68 gnd C_bl
Rb_53_69 bit_53_69 bit_53_70 R_bl
Rbb_53_69 bitb_53_69 bitb_53_70 R_bl
Cb_53_69 bit_53_69 gnd C_bl
Cbb_53_69 bitb_53_69 gnd C_bl
Rb_53_70 bit_53_70 bit_53_71 R_bl
Rbb_53_70 bitb_53_70 bitb_53_71 R_bl
Cb_53_70 bit_53_70 gnd C_bl
Cbb_53_70 bitb_53_70 gnd C_bl
Rb_53_71 bit_53_71 bit_53_72 R_bl
Rbb_53_71 bitb_53_71 bitb_53_72 R_bl
Cb_53_71 bit_53_71 gnd C_bl
Cbb_53_71 bitb_53_71 gnd C_bl
Rb_53_72 bit_53_72 bit_53_73 R_bl
Rbb_53_72 bitb_53_72 bitb_53_73 R_bl
Cb_53_72 bit_53_72 gnd C_bl
Cbb_53_72 bitb_53_72 gnd C_bl
Rb_53_73 bit_53_73 bit_53_74 R_bl
Rbb_53_73 bitb_53_73 bitb_53_74 R_bl
Cb_53_73 bit_53_73 gnd C_bl
Cbb_53_73 bitb_53_73 gnd C_bl
Rb_53_74 bit_53_74 bit_53_75 R_bl
Rbb_53_74 bitb_53_74 bitb_53_75 R_bl
Cb_53_74 bit_53_74 gnd C_bl
Cbb_53_74 bitb_53_74 gnd C_bl
Rb_53_75 bit_53_75 bit_53_76 R_bl
Rbb_53_75 bitb_53_75 bitb_53_76 R_bl
Cb_53_75 bit_53_75 gnd C_bl
Cbb_53_75 bitb_53_75 gnd C_bl
Rb_53_76 bit_53_76 bit_53_77 R_bl
Rbb_53_76 bitb_53_76 bitb_53_77 R_bl
Cb_53_76 bit_53_76 gnd C_bl
Cbb_53_76 bitb_53_76 gnd C_bl
Rb_53_77 bit_53_77 bit_53_78 R_bl
Rbb_53_77 bitb_53_77 bitb_53_78 R_bl
Cb_53_77 bit_53_77 gnd C_bl
Cbb_53_77 bitb_53_77 gnd C_bl
Rb_53_78 bit_53_78 bit_53_79 R_bl
Rbb_53_78 bitb_53_78 bitb_53_79 R_bl
Cb_53_78 bit_53_78 gnd C_bl
Cbb_53_78 bitb_53_78 gnd C_bl
Rb_53_79 bit_53_79 bit_53_80 R_bl
Rbb_53_79 bitb_53_79 bitb_53_80 R_bl
Cb_53_79 bit_53_79 gnd C_bl
Cbb_53_79 bitb_53_79 gnd C_bl
Rb_53_80 bit_53_80 bit_53_81 R_bl
Rbb_53_80 bitb_53_80 bitb_53_81 R_bl
Cb_53_80 bit_53_80 gnd C_bl
Cbb_53_80 bitb_53_80 gnd C_bl
Rb_53_81 bit_53_81 bit_53_82 R_bl
Rbb_53_81 bitb_53_81 bitb_53_82 R_bl
Cb_53_81 bit_53_81 gnd C_bl
Cbb_53_81 bitb_53_81 gnd C_bl
Rb_53_82 bit_53_82 bit_53_83 R_bl
Rbb_53_82 bitb_53_82 bitb_53_83 R_bl
Cb_53_82 bit_53_82 gnd C_bl
Cbb_53_82 bitb_53_82 gnd C_bl
Rb_53_83 bit_53_83 bit_53_84 R_bl
Rbb_53_83 bitb_53_83 bitb_53_84 R_bl
Cb_53_83 bit_53_83 gnd C_bl
Cbb_53_83 bitb_53_83 gnd C_bl
Rb_53_84 bit_53_84 bit_53_85 R_bl
Rbb_53_84 bitb_53_84 bitb_53_85 R_bl
Cb_53_84 bit_53_84 gnd C_bl
Cbb_53_84 bitb_53_84 gnd C_bl
Rb_53_85 bit_53_85 bit_53_86 R_bl
Rbb_53_85 bitb_53_85 bitb_53_86 R_bl
Cb_53_85 bit_53_85 gnd C_bl
Cbb_53_85 bitb_53_85 gnd C_bl
Rb_53_86 bit_53_86 bit_53_87 R_bl
Rbb_53_86 bitb_53_86 bitb_53_87 R_bl
Cb_53_86 bit_53_86 gnd C_bl
Cbb_53_86 bitb_53_86 gnd C_bl
Rb_53_87 bit_53_87 bit_53_88 R_bl
Rbb_53_87 bitb_53_87 bitb_53_88 R_bl
Cb_53_87 bit_53_87 gnd C_bl
Cbb_53_87 bitb_53_87 gnd C_bl
Rb_53_88 bit_53_88 bit_53_89 R_bl
Rbb_53_88 bitb_53_88 bitb_53_89 R_bl
Cb_53_88 bit_53_88 gnd C_bl
Cbb_53_88 bitb_53_88 gnd C_bl
Rb_53_89 bit_53_89 bit_53_90 R_bl
Rbb_53_89 bitb_53_89 bitb_53_90 R_bl
Cb_53_89 bit_53_89 gnd C_bl
Cbb_53_89 bitb_53_89 gnd C_bl
Rb_53_90 bit_53_90 bit_53_91 R_bl
Rbb_53_90 bitb_53_90 bitb_53_91 R_bl
Cb_53_90 bit_53_90 gnd C_bl
Cbb_53_90 bitb_53_90 gnd C_bl
Rb_53_91 bit_53_91 bit_53_92 R_bl
Rbb_53_91 bitb_53_91 bitb_53_92 R_bl
Cb_53_91 bit_53_91 gnd C_bl
Cbb_53_91 bitb_53_91 gnd C_bl
Rb_53_92 bit_53_92 bit_53_93 R_bl
Rbb_53_92 bitb_53_92 bitb_53_93 R_bl
Cb_53_92 bit_53_92 gnd C_bl
Cbb_53_92 bitb_53_92 gnd C_bl
Rb_53_93 bit_53_93 bit_53_94 R_bl
Rbb_53_93 bitb_53_93 bitb_53_94 R_bl
Cb_53_93 bit_53_93 gnd C_bl
Cbb_53_93 bitb_53_93 gnd C_bl
Rb_53_94 bit_53_94 bit_53_95 R_bl
Rbb_53_94 bitb_53_94 bitb_53_95 R_bl
Cb_53_94 bit_53_94 gnd C_bl
Cbb_53_94 bitb_53_94 gnd C_bl
Rb_53_95 bit_53_95 bit_53_96 R_bl
Rbb_53_95 bitb_53_95 bitb_53_96 R_bl
Cb_53_95 bit_53_95 gnd C_bl
Cbb_53_95 bitb_53_95 gnd C_bl
Rb_53_96 bit_53_96 bit_53_97 R_bl
Rbb_53_96 bitb_53_96 bitb_53_97 R_bl
Cb_53_96 bit_53_96 gnd C_bl
Cbb_53_96 bitb_53_96 gnd C_bl
Rb_53_97 bit_53_97 bit_53_98 R_bl
Rbb_53_97 bitb_53_97 bitb_53_98 R_bl
Cb_53_97 bit_53_97 gnd C_bl
Cbb_53_97 bitb_53_97 gnd C_bl
Rb_53_98 bit_53_98 bit_53_99 R_bl
Rbb_53_98 bitb_53_98 bitb_53_99 R_bl
Cb_53_98 bit_53_98 gnd C_bl
Cbb_53_98 bitb_53_98 gnd C_bl
Rb_53_99 bit_53_99 bit_53_100 R_bl
Rbb_53_99 bitb_53_99 bitb_53_100 R_bl
Cb_53_99 bit_53_99 gnd C_bl
Cbb_53_99 bitb_53_99 gnd C_bl
Rb_54_0 bit_54_0 bit_54_1 R_bl
Rbb_54_0 bitb_54_0 bitb_54_1 R_bl
Cb_54_0 bit_54_0 gnd C_bl
Cbb_54_0 bitb_54_0 gnd C_bl
Rb_54_1 bit_54_1 bit_54_2 R_bl
Rbb_54_1 bitb_54_1 bitb_54_2 R_bl
Cb_54_1 bit_54_1 gnd C_bl
Cbb_54_1 bitb_54_1 gnd C_bl
Rb_54_2 bit_54_2 bit_54_3 R_bl
Rbb_54_2 bitb_54_2 bitb_54_3 R_bl
Cb_54_2 bit_54_2 gnd C_bl
Cbb_54_2 bitb_54_2 gnd C_bl
Rb_54_3 bit_54_3 bit_54_4 R_bl
Rbb_54_3 bitb_54_3 bitb_54_4 R_bl
Cb_54_3 bit_54_3 gnd C_bl
Cbb_54_3 bitb_54_3 gnd C_bl
Rb_54_4 bit_54_4 bit_54_5 R_bl
Rbb_54_4 bitb_54_4 bitb_54_5 R_bl
Cb_54_4 bit_54_4 gnd C_bl
Cbb_54_4 bitb_54_4 gnd C_bl
Rb_54_5 bit_54_5 bit_54_6 R_bl
Rbb_54_5 bitb_54_5 bitb_54_6 R_bl
Cb_54_5 bit_54_5 gnd C_bl
Cbb_54_5 bitb_54_5 gnd C_bl
Rb_54_6 bit_54_6 bit_54_7 R_bl
Rbb_54_6 bitb_54_6 bitb_54_7 R_bl
Cb_54_6 bit_54_6 gnd C_bl
Cbb_54_6 bitb_54_6 gnd C_bl
Rb_54_7 bit_54_7 bit_54_8 R_bl
Rbb_54_7 bitb_54_7 bitb_54_8 R_bl
Cb_54_7 bit_54_7 gnd C_bl
Cbb_54_7 bitb_54_7 gnd C_bl
Rb_54_8 bit_54_8 bit_54_9 R_bl
Rbb_54_8 bitb_54_8 bitb_54_9 R_bl
Cb_54_8 bit_54_8 gnd C_bl
Cbb_54_8 bitb_54_8 gnd C_bl
Rb_54_9 bit_54_9 bit_54_10 R_bl
Rbb_54_9 bitb_54_9 bitb_54_10 R_bl
Cb_54_9 bit_54_9 gnd C_bl
Cbb_54_9 bitb_54_9 gnd C_bl
Rb_54_10 bit_54_10 bit_54_11 R_bl
Rbb_54_10 bitb_54_10 bitb_54_11 R_bl
Cb_54_10 bit_54_10 gnd C_bl
Cbb_54_10 bitb_54_10 gnd C_bl
Rb_54_11 bit_54_11 bit_54_12 R_bl
Rbb_54_11 bitb_54_11 bitb_54_12 R_bl
Cb_54_11 bit_54_11 gnd C_bl
Cbb_54_11 bitb_54_11 gnd C_bl
Rb_54_12 bit_54_12 bit_54_13 R_bl
Rbb_54_12 bitb_54_12 bitb_54_13 R_bl
Cb_54_12 bit_54_12 gnd C_bl
Cbb_54_12 bitb_54_12 gnd C_bl
Rb_54_13 bit_54_13 bit_54_14 R_bl
Rbb_54_13 bitb_54_13 bitb_54_14 R_bl
Cb_54_13 bit_54_13 gnd C_bl
Cbb_54_13 bitb_54_13 gnd C_bl
Rb_54_14 bit_54_14 bit_54_15 R_bl
Rbb_54_14 bitb_54_14 bitb_54_15 R_bl
Cb_54_14 bit_54_14 gnd C_bl
Cbb_54_14 bitb_54_14 gnd C_bl
Rb_54_15 bit_54_15 bit_54_16 R_bl
Rbb_54_15 bitb_54_15 bitb_54_16 R_bl
Cb_54_15 bit_54_15 gnd C_bl
Cbb_54_15 bitb_54_15 gnd C_bl
Rb_54_16 bit_54_16 bit_54_17 R_bl
Rbb_54_16 bitb_54_16 bitb_54_17 R_bl
Cb_54_16 bit_54_16 gnd C_bl
Cbb_54_16 bitb_54_16 gnd C_bl
Rb_54_17 bit_54_17 bit_54_18 R_bl
Rbb_54_17 bitb_54_17 bitb_54_18 R_bl
Cb_54_17 bit_54_17 gnd C_bl
Cbb_54_17 bitb_54_17 gnd C_bl
Rb_54_18 bit_54_18 bit_54_19 R_bl
Rbb_54_18 bitb_54_18 bitb_54_19 R_bl
Cb_54_18 bit_54_18 gnd C_bl
Cbb_54_18 bitb_54_18 gnd C_bl
Rb_54_19 bit_54_19 bit_54_20 R_bl
Rbb_54_19 bitb_54_19 bitb_54_20 R_bl
Cb_54_19 bit_54_19 gnd C_bl
Cbb_54_19 bitb_54_19 gnd C_bl
Rb_54_20 bit_54_20 bit_54_21 R_bl
Rbb_54_20 bitb_54_20 bitb_54_21 R_bl
Cb_54_20 bit_54_20 gnd C_bl
Cbb_54_20 bitb_54_20 gnd C_bl
Rb_54_21 bit_54_21 bit_54_22 R_bl
Rbb_54_21 bitb_54_21 bitb_54_22 R_bl
Cb_54_21 bit_54_21 gnd C_bl
Cbb_54_21 bitb_54_21 gnd C_bl
Rb_54_22 bit_54_22 bit_54_23 R_bl
Rbb_54_22 bitb_54_22 bitb_54_23 R_bl
Cb_54_22 bit_54_22 gnd C_bl
Cbb_54_22 bitb_54_22 gnd C_bl
Rb_54_23 bit_54_23 bit_54_24 R_bl
Rbb_54_23 bitb_54_23 bitb_54_24 R_bl
Cb_54_23 bit_54_23 gnd C_bl
Cbb_54_23 bitb_54_23 gnd C_bl
Rb_54_24 bit_54_24 bit_54_25 R_bl
Rbb_54_24 bitb_54_24 bitb_54_25 R_bl
Cb_54_24 bit_54_24 gnd C_bl
Cbb_54_24 bitb_54_24 gnd C_bl
Rb_54_25 bit_54_25 bit_54_26 R_bl
Rbb_54_25 bitb_54_25 bitb_54_26 R_bl
Cb_54_25 bit_54_25 gnd C_bl
Cbb_54_25 bitb_54_25 gnd C_bl
Rb_54_26 bit_54_26 bit_54_27 R_bl
Rbb_54_26 bitb_54_26 bitb_54_27 R_bl
Cb_54_26 bit_54_26 gnd C_bl
Cbb_54_26 bitb_54_26 gnd C_bl
Rb_54_27 bit_54_27 bit_54_28 R_bl
Rbb_54_27 bitb_54_27 bitb_54_28 R_bl
Cb_54_27 bit_54_27 gnd C_bl
Cbb_54_27 bitb_54_27 gnd C_bl
Rb_54_28 bit_54_28 bit_54_29 R_bl
Rbb_54_28 bitb_54_28 bitb_54_29 R_bl
Cb_54_28 bit_54_28 gnd C_bl
Cbb_54_28 bitb_54_28 gnd C_bl
Rb_54_29 bit_54_29 bit_54_30 R_bl
Rbb_54_29 bitb_54_29 bitb_54_30 R_bl
Cb_54_29 bit_54_29 gnd C_bl
Cbb_54_29 bitb_54_29 gnd C_bl
Rb_54_30 bit_54_30 bit_54_31 R_bl
Rbb_54_30 bitb_54_30 bitb_54_31 R_bl
Cb_54_30 bit_54_30 gnd C_bl
Cbb_54_30 bitb_54_30 gnd C_bl
Rb_54_31 bit_54_31 bit_54_32 R_bl
Rbb_54_31 bitb_54_31 bitb_54_32 R_bl
Cb_54_31 bit_54_31 gnd C_bl
Cbb_54_31 bitb_54_31 gnd C_bl
Rb_54_32 bit_54_32 bit_54_33 R_bl
Rbb_54_32 bitb_54_32 bitb_54_33 R_bl
Cb_54_32 bit_54_32 gnd C_bl
Cbb_54_32 bitb_54_32 gnd C_bl
Rb_54_33 bit_54_33 bit_54_34 R_bl
Rbb_54_33 bitb_54_33 bitb_54_34 R_bl
Cb_54_33 bit_54_33 gnd C_bl
Cbb_54_33 bitb_54_33 gnd C_bl
Rb_54_34 bit_54_34 bit_54_35 R_bl
Rbb_54_34 bitb_54_34 bitb_54_35 R_bl
Cb_54_34 bit_54_34 gnd C_bl
Cbb_54_34 bitb_54_34 gnd C_bl
Rb_54_35 bit_54_35 bit_54_36 R_bl
Rbb_54_35 bitb_54_35 bitb_54_36 R_bl
Cb_54_35 bit_54_35 gnd C_bl
Cbb_54_35 bitb_54_35 gnd C_bl
Rb_54_36 bit_54_36 bit_54_37 R_bl
Rbb_54_36 bitb_54_36 bitb_54_37 R_bl
Cb_54_36 bit_54_36 gnd C_bl
Cbb_54_36 bitb_54_36 gnd C_bl
Rb_54_37 bit_54_37 bit_54_38 R_bl
Rbb_54_37 bitb_54_37 bitb_54_38 R_bl
Cb_54_37 bit_54_37 gnd C_bl
Cbb_54_37 bitb_54_37 gnd C_bl
Rb_54_38 bit_54_38 bit_54_39 R_bl
Rbb_54_38 bitb_54_38 bitb_54_39 R_bl
Cb_54_38 bit_54_38 gnd C_bl
Cbb_54_38 bitb_54_38 gnd C_bl
Rb_54_39 bit_54_39 bit_54_40 R_bl
Rbb_54_39 bitb_54_39 bitb_54_40 R_bl
Cb_54_39 bit_54_39 gnd C_bl
Cbb_54_39 bitb_54_39 gnd C_bl
Rb_54_40 bit_54_40 bit_54_41 R_bl
Rbb_54_40 bitb_54_40 bitb_54_41 R_bl
Cb_54_40 bit_54_40 gnd C_bl
Cbb_54_40 bitb_54_40 gnd C_bl
Rb_54_41 bit_54_41 bit_54_42 R_bl
Rbb_54_41 bitb_54_41 bitb_54_42 R_bl
Cb_54_41 bit_54_41 gnd C_bl
Cbb_54_41 bitb_54_41 gnd C_bl
Rb_54_42 bit_54_42 bit_54_43 R_bl
Rbb_54_42 bitb_54_42 bitb_54_43 R_bl
Cb_54_42 bit_54_42 gnd C_bl
Cbb_54_42 bitb_54_42 gnd C_bl
Rb_54_43 bit_54_43 bit_54_44 R_bl
Rbb_54_43 bitb_54_43 bitb_54_44 R_bl
Cb_54_43 bit_54_43 gnd C_bl
Cbb_54_43 bitb_54_43 gnd C_bl
Rb_54_44 bit_54_44 bit_54_45 R_bl
Rbb_54_44 bitb_54_44 bitb_54_45 R_bl
Cb_54_44 bit_54_44 gnd C_bl
Cbb_54_44 bitb_54_44 gnd C_bl
Rb_54_45 bit_54_45 bit_54_46 R_bl
Rbb_54_45 bitb_54_45 bitb_54_46 R_bl
Cb_54_45 bit_54_45 gnd C_bl
Cbb_54_45 bitb_54_45 gnd C_bl
Rb_54_46 bit_54_46 bit_54_47 R_bl
Rbb_54_46 bitb_54_46 bitb_54_47 R_bl
Cb_54_46 bit_54_46 gnd C_bl
Cbb_54_46 bitb_54_46 gnd C_bl
Rb_54_47 bit_54_47 bit_54_48 R_bl
Rbb_54_47 bitb_54_47 bitb_54_48 R_bl
Cb_54_47 bit_54_47 gnd C_bl
Cbb_54_47 bitb_54_47 gnd C_bl
Rb_54_48 bit_54_48 bit_54_49 R_bl
Rbb_54_48 bitb_54_48 bitb_54_49 R_bl
Cb_54_48 bit_54_48 gnd C_bl
Cbb_54_48 bitb_54_48 gnd C_bl
Rb_54_49 bit_54_49 bit_54_50 R_bl
Rbb_54_49 bitb_54_49 bitb_54_50 R_bl
Cb_54_49 bit_54_49 gnd C_bl
Cbb_54_49 bitb_54_49 gnd C_bl
Rb_54_50 bit_54_50 bit_54_51 R_bl
Rbb_54_50 bitb_54_50 bitb_54_51 R_bl
Cb_54_50 bit_54_50 gnd C_bl
Cbb_54_50 bitb_54_50 gnd C_bl
Rb_54_51 bit_54_51 bit_54_52 R_bl
Rbb_54_51 bitb_54_51 bitb_54_52 R_bl
Cb_54_51 bit_54_51 gnd C_bl
Cbb_54_51 bitb_54_51 gnd C_bl
Rb_54_52 bit_54_52 bit_54_53 R_bl
Rbb_54_52 bitb_54_52 bitb_54_53 R_bl
Cb_54_52 bit_54_52 gnd C_bl
Cbb_54_52 bitb_54_52 gnd C_bl
Rb_54_53 bit_54_53 bit_54_54 R_bl
Rbb_54_53 bitb_54_53 bitb_54_54 R_bl
Cb_54_53 bit_54_53 gnd C_bl
Cbb_54_53 bitb_54_53 gnd C_bl
Rb_54_54 bit_54_54 bit_54_55 R_bl
Rbb_54_54 bitb_54_54 bitb_54_55 R_bl
Cb_54_54 bit_54_54 gnd C_bl
Cbb_54_54 bitb_54_54 gnd C_bl
Rb_54_55 bit_54_55 bit_54_56 R_bl
Rbb_54_55 bitb_54_55 bitb_54_56 R_bl
Cb_54_55 bit_54_55 gnd C_bl
Cbb_54_55 bitb_54_55 gnd C_bl
Rb_54_56 bit_54_56 bit_54_57 R_bl
Rbb_54_56 bitb_54_56 bitb_54_57 R_bl
Cb_54_56 bit_54_56 gnd C_bl
Cbb_54_56 bitb_54_56 gnd C_bl
Rb_54_57 bit_54_57 bit_54_58 R_bl
Rbb_54_57 bitb_54_57 bitb_54_58 R_bl
Cb_54_57 bit_54_57 gnd C_bl
Cbb_54_57 bitb_54_57 gnd C_bl
Rb_54_58 bit_54_58 bit_54_59 R_bl
Rbb_54_58 bitb_54_58 bitb_54_59 R_bl
Cb_54_58 bit_54_58 gnd C_bl
Cbb_54_58 bitb_54_58 gnd C_bl
Rb_54_59 bit_54_59 bit_54_60 R_bl
Rbb_54_59 bitb_54_59 bitb_54_60 R_bl
Cb_54_59 bit_54_59 gnd C_bl
Cbb_54_59 bitb_54_59 gnd C_bl
Rb_54_60 bit_54_60 bit_54_61 R_bl
Rbb_54_60 bitb_54_60 bitb_54_61 R_bl
Cb_54_60 bit_54_60 gnd C_bl
Cbb_54_60 bitb_54_60 gnd C_bl
Rb_54_61 bit_54_61 bit_54_62 R_bl
Rbb_54_61 bitb_54_61 bitb_54_62 R_bl
Cb_54_61 bit_54_61 gnd C_bl
Cbb_54_61 bitb_54_61 gnd C_bl
Rb_54_62 bit_54_62 bit_54_63 R_bl
Rbb_54_62 bitb_54_62 bitb_54_63 R_bl
Cb_54_62 bit_54_62 gnd C_bl
Cbb_54_62 bitb_54_62 gnd C_bl
Rb_54_63 bit_54_63 bit_54_64 R_bl
Rbb_54_63 bitb_54_63 bitb_54_64 R_bl
Cb_54_63 bit_54_63 gnd C_bl
Cbb_54_63 bitb_54_63 gnd C_bl
Rb_54_64 bit_54_64 bit_54_65 R_bl
Rbb_54_64 bitb_54_64 bitb_54_65 R_bl
Cb_54_64 bit_54_64 gnd C_bl
Cbb_54_64 bitb_54_64 gnd C_bl
Rb_54_65 bit_54_65 bit_54_66 R_bl
Rbb_54_65 bitb_54_65 bitb_54_66 R_bl
Cb_54_65 bit_54_65 gnd C_bl
Cbb_54_65 bitb_54_65 gnd C_bl
Rb_54_66 bit_54_66 bit_54_67 R_bl
Rbb_54_66 bitb_54_66 bitb_54_67 R_bl
Cb_54_66 bit_54_66 gnd C_bl
Cbb_54_66 bitb_54_66 gnd C_bl
Rb_54_67 bit_54_67 bit_54_68 R_bl
Rbb_54_67 bitb_54_67 bitb_54_68 R_bl
Cb_54_67 bit_54_67 gnd C_bl
Cbb_54_67 bitb_54_67 gnd C_bl
Rb_54_68 bit_54_68 bit_54_69 R_bl
Rbb_54_68 bitb_54_68 bitb_54_69 R_bl
Cb_54_68 bit_54_68 gnd C_bl
Cbb_54_68 bitb_54_68 gnd C_bl
Rb_54_69 bit_54_69 bit_54_70 R_bl
Rbb_54_69 bitb_54_69 bitb_54_70 R_bl
Cb_54_69 bit_54_69 gnd C_bl
Cbb_54_69 bitb_54_69 gnd C_bl
Rb_54_70 bit_54_70 bit_54_71 R_bl
Rbb_54_70 bitb_54_70 bitb_54_71 R_bl
Cb_54_70 bit_54_70 gnd C_bl
Cbb_54_70 bitb_54_70 gnd C_bl
Rb_54_71 bit_54_71 bit_54_72 R_bl
Rbb_54_71 bitb_54_71 bitb_54_72 R_bl
Cb_54_71 bit_54_71 gnd C_bl
Cbb_54_71 bitb_54_71 gnd C_bl
Rb_54_72 bit_54_72 bit_54_73 R_bl
Rbb_54_72 bitb_54_72 bitb_54_73 R_bl
Cb_54_72 bit_54_72 gnd C_bl
Cbb_54_72 bitb_54_72 gnd C_bl
Rb_54_73 bit_54_73 bit_54_74 R_bl
Rbb_54_73 bitb_54_73 bitb_54_74 R_bl
Cb_54_73 bit_54_73 gnd C_bl
Cbb_54_73 bitb_54_73 gnd C_bl
Rb_54_74 bit_54_74 bit_54_75 R_bl
Rbb_54_74 bitb_54_74 bitb_54_75 R_bl
Cb_54_74 bit_54_74 gnd C_bl
Cbb_54_74 bitb_54_74 gnd C_bl
Rb_54_75 bit_54_75 bit_54_76 R_bl
Rbb_54_75 bitb_54_75 bitb_54_76 R_bl
Cb_54_75 bit_54_75 gnd C_bl
Cbb_54_75 bitb_54_75 gnd C_bl
Rb_54_76 bit_54_76 bit_54_77 R_bl
Rbb_54_76 bitb_54_76 bitb_54_77 R_bl
Cb_54_76 bit_54_76 gnd C_bl
Cbb_54_76 bitb_54_76 gnd C_bl
Rb_54_77 bit_54_77 bit_54_78 R_bl
Rbb_54_77 bitb_54_77 bitb_54_78 R_bl
Cb_54_77 bit_54_77 gnd C_bl
Cbb_54_77 bitb_54_77 gnd C_bl
Rb_54_78 bit_54_78 bit_54_79 R_bl
Rbb_54_78 bitb_54_78 bitb_54_79 R_bl
Cb_54_78 bit_54_78 gnd C_bl
Cbb_54_78 bitb_54_78 gnd C_bl
Rb_54_79 bit_54_79 bit_54_80 R_bl
Rbb_54_79 bitb_54_79 bitb_54_80 R_bl
Cb_54_79 bit_54_79 gnd C_bl
Cbb_54_79 bitb_54_79 gnd C_bl
Rb_54_80 bit_54_80 bit_54_81 R_bl
Rbb_54_80 bitb_54_80 bitb_54_81 R_bl
Cb_54_80 bit_54_80 gnd C_bl
Cbb_54_80 bitb_54_80 gnd C_bl
Rb_54_81 bit_54_81 bit_54_82 R_bl
Rbb_54_81 bitb_54_81 bitb_54_82 R_bl
Cb_54_81 bit_54_81 gnd C_bl
Cbb_54_81 bitb_54_81 gnd C_bl
Rb_54_82 bit_54_82 bit_54_83 R_bl
Rbb_54_82 bitb_54_82 bitb_54_83 R_bl
Cb_54_82 bit_54_82 gnd C_bl
Cbb_54_82 bitb_54_82 gnd C_bl
Rb_54_83 bit_54_83 bit_54_84 R_bl
Rbb_54_83 bitb_54_83 bitb_54_84 R_bl
Cb_54_83 bit_54_83 gnd C_bl
Cbb_54_83 bitb_54_83 gnd C_bl
Rb_54_84 bit_54_84 bit_54_85 R_bl
Rbb_54_84 bitb_54_84 bitb_54_85 R_bl
Cb_54_84 bit_54_84 gnd C_bl
Cbb_54_84 bitb_54_84 gnd C_bl
Rb_54_85 bit_54_85 bit_54_86 R_bl
Rbb_54_85 bitb_54_85 bitb_54_86 R_bl
Cb_54_85 bit_54_85 gnd C_bl
Cbb_54_85 bitb_54_85 gnd C_bl
Rb_54_86 bit_54_86 bit_54_87 R_bl
Rbb_54_86 bitb_54_86 bitb_54_87 R_bl
Cb_54_86 bit_54_86 gnd C_bl
Cbb_54_86 bitb_54_86 gnd C_bl
Rb_54_87 bit_54_87 bit_54_88 R_bl
Rbb_54_87 bitb_54_87 bitb_54_88 R_bl
Cb_54_87 bit_54_87 gnd C_bl
Cbb_54_87 bitb_54_87 gnd C_bl
Rb_54_88 bit_54_88 bit_54_89 R_bl
Rbb_54_88 bitb_54_88 bitb_54_89 R_bl
Cb_54_88 bit_54_88 gnd C_bl
Cbb_54_88 bitb_54_88 gnd C_bl
Rb_54_89 bit_54_89 bit_54_90 R_bl
Rbb_54_89 bitb_54_89 bitb_54_90 R_bl
Cb_54_89 bit_54_89 gnd C_bl
Cbb_54_89 bitb_54_89 gnd C_bl
Rb_54_90 bit_54_90 bit_54_91 R_bl
Rbb_54_90 bitb_54_90 bitb_54_91 R_bl
Cb_54_90 bit_54_90 gnd C_bl
Cbb_54_90 bitb_54_90 gnd C_bl
Rb_54_91 bit_54_91 bit_54_92 R_bl
Rbb_54_91 bitb_54_91 bitb_54_92 R_bl
Cb_54_91 bit_54_91 gnd C_bl
Cbb_54_91 bitb_54_91 gnd C_bl
Rb_54_92 bit_54_92 bit_54_93 R_bl
Rbb_54_92 bitb_54_92 bitb_54_93 R_bl
Cb_54_92 bit_54_92 gnd C_bl
Cbb_54_92 bitb_54_92 gnd C_bl
Rb_54_93 bit_54_93 bit_54_94 R_bl
Rbb_54_93 bitb_54_93 bitb_54_94 R_bl
Cb_54_93 bit_54_93 gnd C_bl
Cbb_54_93 bitb_54_93 gnd C_bl
Rb_54_94 bit_54_94 bit_54_95 R_bl
Rbb_54_94 bitb_54_94 bitb_54_95 R_bl
Cb_54_94 bit_54_94 gnd C_bl
Cbb_54_94 bitb_54_94 gnd C_bl
Rb_54_95 bit_54_95 bit_54_96 R_bl
Rbb_54_95 bitb_54_95 bitb_54_96 R_bl
Cb_54_95 bit_54_95 gnd C_bl
Cbb_54_95 bitb_54_95 gnd C_bl
Rb_54_96 bit_54_96 bit_54_97 R_bl
Rbb_54_96 bitb_54_96 bitb_54_97 R_bl
Cb_54_96 bit_54_96 gnd C_bl
Cbb_54_96 bitb_54_96 gnd C_bl
Rb_54_97 bit_54_97 bit_54_98 R_bl
Rbb_54_97 bitb_54_97 bitb_54_98 R_bl
Cb_54_97 bit_54_97 gnd C_bl
Cbb_54_97 bitb_54_97 gnd C_bl
Rb_54_98 bit_54_98 bit_54_99 R_bl
Rbb_54_98 bitb_54_98 bitb_54_99 R_bl
Cb_54_98 bit_54_98 gnd C_bl
Cbb_54_98 bitb_54_98 gnd C_bl
Rb_54_99 bit_54_99 bit_54_100 R_bl
Rbb_54_99 bitb_54_99 bitb_54_100 R_bl
Cb_54_99 bit_54_99 gnd C_bl
Cbb_54_99 bitb_54_99 gnd C_bl
Rb_55_0 bit_55_0 bit_55_1 R_bl
Rbb_55_0 bitb_55_0 bitb_55_1 R_bl
Cb_55_0 bit_55_0 gnd C_bl
Cbb_55_0 bitb_55_0 gnd C_bl
Rb_55_1 bit_55_1 bit_55_2 R_bl
Rbb_55_1 bitb_55_1 bitb_55_2 R_bl
Cb_55_1 bit_55_1 gnd C_bl
Cbb_55_1 bitb_55_1 gnd C_bl
Rb_55_2 bit_55_2 bit_55_3 R_bl
Rbb_55_2 bitb_55_2 bitb_55_3 R_bl
Cb_55_2 bit_55_2 gnd C_bl
Cbb_55_2 bitb_55_2 gnd C_bl
Rb_55_3 bit_55_3 bit_55_4 R_bl
Rbb_55_3 bitb_55_3 bitb_55_4 R_bl
Cb_55_3 bit_55_3 gnd C_bl
Cbb_55_3 bitb_55_3 gnd C_bl
Rb_55_4 bit_55_4 bit_55_5 R_bl
Rbb_55_4 bitb_55_4 bitb_55_5 R_bl
Cb_55_4 bit_55_4 gnd C_bl
Cbb_55_4 bitb_55_4 gnd C_bl
Rb_55_5 bit_55_5 bit_55_6 R_bl
Rbb_55_5 bitb_55_5 bitb_55_6 R_bl
Cb_55_5 bit_55_5 gnd C_bl
Cbb_55_5 bitb_55_5 gnd C_bl
Rb_55_6 bit_55_6 bit_55_7 R_bl
Rbb_55_6 bitb_55_6 bitb_55_7 R_bl
Cb_55_6 bit_55_6 gnd C_bl
Cbb_55_6 bitb_55_6 gnd C_bl
Rb_55_7 bit_55_7 bit_55_8 R_bl
Rbb_55_7 bitb_55_7 bitb_55_8 R_bl
Cb_55_7 bit_55_7 gnd C_bl
Cbb_55_7 bitb_55_7 gnd C_bl
Rb_55_8 bit_55_8 bit_55_9 R_bl
Rbb_55_8 bitb_55_8 bitb_55_9 R_bl
Cb_55_8 bit_55_8 gnd C_bl
Cbb_55_8 bitb_55_8 gnd C_bl
Rb_55_9 bit_55_9 bit_55_10 R_bl
Rbb_55_9 bitb_55_9 bitb_55_10 R_bl
Cb_55_9 bit_55_9 gnd C_bl
Cbb_55_9 bitb_55_9 gnd C_bl
Rb_55_10 bit_55_10 bit_55_11 R_bl
Rbb_55_10 bitb_55_10 bitb_55_11 R_bl
Cb_55_10 bit_55_10 gnd C_bl
Cbb_55_10 bitb_55_10 gnd C_bl
Rb_55_11 bit_55_11 bit_55_12 R_bl
Rbb_55_11 bitb_55_11 bitb_55_12 R_bl
Cb_55_11 bit_55_11 gnd C_bl
Cbb_55_11 bitb_55_11 gnd C_bl
Rb_55_12 bit_55_12 bit_55_13 R_bl
Rbb_55_12 bitb_55_12 bitb_55_13 R_bl
Cb_55_12 bit_55_12 gnd C_bl
Cbb_55_12 bitb_55_12 gnd C_bl
Rb_55_13 bit_55_13 bit_55_14 R_bl
Rbb_55_13 bitb_55_13 bitb_55_14 R_bl
Cb_55_13 bit_55_13 gnd C_bl
Cbb_55_13 bitb_55_13 gnd C_bl
Rb_55_14 bit_55_14 bit_55_15 R_bl
Rbb_55_14 bitb_55_14 bitb_55_15 R_bl
Cb_55_14 bit_55_14 gnd C_bl
Cbb_55_14 bitb_55_14 gnd C_bl
Rb_55_15 bit_55_15 bit_55_16 R_bl
Rbb_55_15 bitb_55_15 bitb_55_16 R_bl
Cb_55_15 bit_55_15 gnd C_bl
Cbb_55_15 bitb_55_15 gnd C_bl
Rb_55_16 bit_55_16 bit_55_17 R_bl
Rbb_55_16 bitb_55_16 bitb_55_17 R_bl
Cb_55_16 bit_55_16 gnd C_bl
Cbb_55_16 bitb_55_16 gnd C_bl
Rb_55_17 bit_55_17 bit_55_18 R_bl
Rbb_55_17 bitb_55_17 bitb_55_18 R_bl
Cb_55_17 bit_55_17 gnd C_bl
Cbb_55_17 bitb_55_17 gnd C_bl
Rb_55_18 bit_55_18 bit_55_19 R_bl
Rbb_55_18 bitb_55_18 bitb_55_19 R_bl
Cb_55_18 bit_55_18 gnd C_bl
Cbb_55_18 bitb_55_18 gnd C_bl
Rb_55_19 bit_55_19 bit_55_20 R_bl
Rbb_55_19 bitb_55_19 bitb_55_20 R_bl
Cb_55_19 bit_55_19 gnd C_bl
Cbb_55_19 bitb_55_19 gnd C_bl
Rb_55_20 bit_55_20 bit_55_21 R_bl
Rbb_55_20 bitb_55_20 bitb_55_21 R_bl
Cb_55_20 bit_55_20 gnd C_bl
Cbb_55_20 bitb_55_20 gnd C_bl
Rb_55_21 bit_55_21 bit_55_22 R_bl
Rbb_55_21 bitb_55_21 bitb_55_22 R_bl
Cb_55_21 bit_55_21 gnd C_bl
Cbb_55_21 bitb_55_21 gnd C_bl
Rb_55_22 bit_55_22 bit_55_23 R_bl
Rbb_55_22 bitb_55_22 bitb_55_23 R_bl
Cb_55_22 bit_55_22 gnd C_bl
Cbb_55_22 bitb_55_22 gnd C_bl
Rb_55_23 bit_55_23 bit_55_24 R_bl
Rbb_55_23 bitb_55_23 bitb_55_24 R_bl
Cb_55_23 bit_55_23 gnd C_bl
Cbb_55_23 bitb_55_23 gnd C_bl
Rb_55_24 bit_55_24 bit_55_25 R_bl
Rbb_55_24 bitb_55_24 bitb_55_25 R_bl
Cb_55_24 bit_55_24 gnd C_bl
Cbb_55_24 bitb_55_24 gnd C_bl
Rb_55_25 bit_55_25 bit_55_26 R_bl
Rbb_55_25 bitb_55_25 bitb_55_26 R_bl
Cb_55_25 bit_55_25 gnd C_bl
Cbb_55_25 bitb_55_25 gnd C_bl
Rb_55_26 bit_55_26 bit_55_27 R_bl
Rbb_55_26 bitb_55_26 bitb_55_27 R_bl
Cb_55_26 bit_55_26 gnd C_bl
Cbb_55_26 bitb_55_26 gnd C_bl
Rb_55_27 bit_55_27 bit_55_28 R_bl
Rbb_55_27 bitb_55_27 bitb_55_28 R_bl
Cb_55_27 bit_55_27 gnd C_bl
Cbb_55_27 bitb_55_27 gnd C_bl
Rb_55_28 bit_55_28 bit_55_29 R_bl
Rbb_55_28 bitb_55_28 bitb_55_29 R_bl
Cb_55_28 bit_55_28 gnd C_bl
Cbb_55_28 bitb_55_28 gnd C_bl
Rb_55_29 bit_55_29 bit_55_30 R_bl
Rbb_55_29 bitb_55_29 bitb_55_30 R_bl
Cb_55_29 bit_55_29 gnd C_bl
Cbb_55_29 bitb_55_29 gnd C_bl
Rb_55_30 bit_55_30 bit_55_31 R_bl
Rbb_55_30 bitb_55_30 bitb_55_31 R_bl
Cb_55_30 bit_55_30 gnd C_bl
Cbb_55_30 bitb_55_30 gnd C_bl
Rb_55_31 bit_55_31 bit_55_32 R_bl
Rbb_55_31 bitb_55_31 bitb_55_32 R_bl
Cb_55_31 bit_55_31 gnd C_bl
Cbb_55_31 bitb_55_31 gnd C_bl
Rb_55_32 bit_55_32 bit_55_33 R_bl
Rbb_55_32 bitb_55_32 bitb_55_33 R_bl
Cb_55_32 bit_55_32 gnd C_bl
Cbb_55_32 bitb_55_32 gnd C_bl
Rb_55_33 bit_55_33 bit_55_34 R_bl
Rbb_55_33 bitb_55_33 bitb_55_34 R_bl
Cb_55_33 bit_55_33 gnd C_bl
Cbb_55_33 bitb_55_33 gnd C_bl
Rb_55_34 bit_55_34 bit_55_35 R_bl
Rbb_55_34 bitb_55_34 bitb_55_35 R_bl
Cb_55_34 bit_55_34 gnd C_bl
Cbb_55_34 bitb_55_34 gnd C_bl
Rb_55_35 bit_55_35 bit_55_36 R_bl
Rbb_55_35 bitb_55_35 bitb_55_36 R_bl
Cb_55_35 bit_55_35 gnd C_bl
Cbb_55_35 bitb_55_35 gnd C_bl
Rb_55_36 bit_55_36 bit_55_37 R_bl
Rbb_55_36 bitb_55_36 bitb_55_37 R_bl
Cb_55_36 bit_55_36 gnd C_bl
Cbb_55_36 bitb_55_36 gnd C_bl
Rb_55_37 bit_55_37 bit_55_38 R_bl
Rbb_55_37 bitb_55_37 bitb_55_38 R_bl
Cb_55_37 bit_55_37 gnd C_bl
Cbb_55_37 bitb_55_37 gnd C_bl
Rb_55_38 bit_55_38 bit_55_39 R_bl
Rbb_55_38 bitb_55_38 bitb_55_39 R_bl
Cb_55_38 bit_55_38 gnd C_bl
Cbb_55_38 bitb_55_38 gnd C_bl
Rb_55_39 bit_55_39 bit_55_40 R_bl
Rbb_55_39 bitb_55_39 bitb_55_40 R_bl
Cb_55_39 bit_55_39 gnd C_bl
Cbb_55_39 bitb_55_39 gnd C_bl
Rb_55_40 bit_55_40 bit_55_41 R_bl
Rbb_55_40 bitb_55_40 bitb_55_41 R_bl
Cb_55_40 bit_55_40 gnd C_bl
Cbb_55_40 bitb_55_40 gnd C_bl
Rb_55_41 bit_55_41 bit_55_42 R_bl
Rbb_55_41 bitb_55_41 bitb_55_42 R_bl
Cb_55_41 bit_55_41 gnd C_bl
Cbb_55_41 bitb_55_41 gnd C_bl
Rb_55_42 bit_55_42 bit_55_43 R_bl
Rbb_55_42 bitb_55_42 bitb_55_43 R_bl
Cb_55_42 bit_55_42 gnd C_bl
Cbb_55_42 bitb_55_42 gnd C_bl
Rb_55_43 bit_55_43 bit_55_44 R_bl
Rbb_55_43 bitb_55_43 bitb_55_44 R_bl
Cb_55_43 bit_55_43 gnd C_bl
Cbb_55_43 bitb_55_43 gnd C_bl
Rb_55_44 bit_55_44 bit_55_45 R_bl
Rbb_55_44 bitb_55_44 bitb_55_45 R_bl
Cb_55_44 bit_55_44 gnd C_bl
Cbb_55_44 bitb_55_44 gnd C_bl
Rb_55_45 bit_55_45 bit_55_46 R_bl
Rbb_55_45 bitb_55_45 bitb_55_46 R_bl
Cb_55_45 bit_55_45 gnd C_bl
Cbb_55_45 bitb_55_45 gnd C_bl
Rb_55_46 bit_55_46 bit_55_47 R_bl
Rbb_55_46 bitb_55_46 bitb_55_47 R_bl
Cb_55_46 bit_55_46 gnd C_bl
Cbb_55_46 bitb_55_46 gnd C_bl
Rb_55_47 bit_55_47 bit_55_48 R_bl
Rbb_55_47 bitb_55_47 bitb_55_48 R_bl
Cb_55_47 bit_55_47 gnd C_bl
Cbb_55_47 bitb_55_47 gnd C_bl
Rb_55_48 bit_55_48 bit_55_49 R_bl
Rbb_55_48 bitb_55_48 bitb_55_49 R_bl
Cb_55_48 bit_55_48 gnd C_bl
Cbb_55_48 bitb_55_48 gnd C_bl
Rb_55_49 bit_55_49 bit_55_50 R_bl
Rbb_55_49 bitb_55_49 bitb_55_50 R_bl
Cb_55_49 bit_55_49 gnd C_bl
Cbb_55_49 bitb_55_49 gnd C_bl
Rb_55_50 bit_55_50 bit_55_51 R_bl
Rbb_55_50 bitb_55_50 bitb_55_51 R_bl
Cb_55_50 bit_55_50 gnd C_bl
Cbb_55_50 bitb_55_50 gnd C_bl
Rb_55_51 bit_55_51 bit_55_52 R_bl
Rbb_55_51 bitb_55_51 bitb_55_52 R_bl
Cb_55_51 bit_55_51 gnd C_bl
Cbb_55_51 bitb_55_51 gnd C_bl
Rb_55_52 bit_55_52 bit_55_53 R_bl
Rbb_55_52 bitb_55_52 bitb_55_53 R_bl
Cb_55_52 bit_55_52 gnd C_bl
Cbb_55_52 bitb_55_52 gnd C_bl
Rb_55_53 bit_55_53 bit_55_54 R_bl
Rbb_55_53 bitb_55_53 bitb_55_54 R_bl
Cb_55_53 bit_55_53 gnd C_bl
Cbb_55_53 bitb_55_53 gnd C_bl
Rb_55_54 bit_55_54 bit_55_55 R_bl
Rbb_55_54 bitb_55_54 bitb_55_55 R_bl
Cb_55_54 bit_55_54 gnd C_bl
Cbb_55_54 bitb_55_54 gnd C_bl
Rb_55_55 bit_55_55 bit_55_56 R_bl
Rbb_55_55 bitb_55_55 bitb_55_56 R_bl
Cb_55_55 bit_55_55 gnd C_bl
Cbb_55_55 bitb_55_55 gnd C_bl
Rb_55_56 bit_55_56 bit_55_57 R_bl
Rbb_55_56 bitb_55_56 bitb_55_57 R_bl
Cb_55_56 bit_55_56 gnd C_bl
Cbb_55_56 bitb_55_56 gnd C_bl
Rb_55_57 bit_55_57 bit_55_58 R_bl
Rbb_55_57 bitb_55_57 bitb_55_58 R_bl
Cb_55_57 bit_55_57 gnd C_bl
Cbb_55_57 bitb_55_57 gnd C_bl
Rb_55_58 bit_55_58 bit_55_59 R_bl
Rbb_55_58 bitb_55_58 bitb_55_59 R_bl
Cb_55_58 bit_55_58 gnd C_bl
Cbb_55_58 bitb_55_58 gnd C_bl
Rb_55_59 bit_55_59 bit_55_60 R_bl
Rbb_55_59 bitb_55_59 bitb_55_60 R_bl
Cb_55_59 bit_55_59 gnd C_bl
Cbb_55_59 bitb_55_59 gnd C_bl
Rb_55_60 bit_55_60 bit_55_61 R_bl
Rbb_55_60 bitb_55_60 bitb_55_61 R_bl
Cb_55_60 bit_55_60 gnd C_bl
Cbb_55_60 bitb_55_60 gnd C_bl
Rb_55_61 bit_55_61 bit_55_62 R_bl
Rbb_55_61 bitb_55_61 bitb_55_62 R_bl
Cb_55_61 bit_55_61 gnd C_bl
Cbb_55_61 bitb_55_61 gnd C_bl
Rb_55_62 bit_55_62 bit_55_63 R_bl
Rbb_55_62 bitb_55_62 bitb_55_63 R_bl
Cb_55_62 bit_55_62 gnd C_bl
Cbb_55_62 bitb_55_62 gnd C_bl
Rb_55_63 bit_55_63 bit_55_64 R_bl
Rbb_55_63 bitb_55_63 bitb_55_64 R_bl
Cb_55_63 bit_55_63 gnd C_bl
Cbb_55_63 bitb_55_63 gnd C_bl
Rb_55_64 bit_55_64 bit_55_65 R_bl
Rbb_55_64 bitb_55_64 bitb_55_65 R_bl
Cb_55_64 bit_55_64 gnd C_bl
Cbb_55_64 bitb_55_64 gnd C_bl
Rb_55_65 bit_55_65 bit_55_66 R_bl
Rbb_55_65 bitb_55_65 bitb_55_66 R_bl
Cb_55_65 bit_55_65 gnd C_bl
Cbb_55_65 bitb_55_65 gnd C_bl
Rb_55_66 bit_55_66 bit_55_67 R_bl
Rbb_55_66 bitb_55_66 bitb_55_67 R_bl
Cb_55_66 bit_55_66 gnd C_bl
Cbb_55_66 bitb_55_66 gnd C_bl
Rb_55_67 bit_55_67 bit_55_68 R_bl
Rbb_55_67 bitb_55_67 bitb_55_68 R_bl
Cb_55_67 bit_55_67 gnd C_bl
Cbb_55_67 bitb_55_67 gnd C_bl
Rb_55_68 bit_55_68 bit_55_69 R_bl
Rbb_55_68 bitb_55_68 bitb_55_69 R_bl
Cb_55_68 bit_55_68 gnd C_bl
Cbb_55_68 bitb_55_68 gnd C_bl
Rb_55_69 bit_55_69 bit_55_70 R_bl
Rbb_55_69 bitb_55_69 bitb_55_70 R_bl
Cb_55_69 bit_55_69 gnd C_bl
Cbb_55_69 bitb_55_69 gnd C_bl
Rb_55_70 bit_55_70 bit_55_71 R_bl
Rbb_55_70 bitb_55_70 bitb_55_71 R_bl
Cb_55_70 bit_55_70 gnd C_bl
Cbb_55_70 bitb_55_70 gnd C_bl
Rb_55_71 bit_55_71 bit_55_72 R_bl
Rbb_55_71 bitb_55_71 bitb_55_72 R_bl
Cb_55_71 bit_55_71 gnd C_bl
Cbb_55_71 bitb_55_71 gnd C_bl
Rb_55_72 bit_55_72 bit_55_73 R_bl
Rbb_55_72 bitb_55_72 bitb_55_73 R_bl
Cb_55_72 bit_55_72 gnd C_bl
Cbb_55_72 bitb_55_72 gnd C_bl
Rb_55_73 bit_55_73 bit_55_74 R_bl
Rbb_55_73 bitb_55_73 bitb_55_74 R_bl
Cb_55_73 bit_55_73 gnd C_bl
Cbb_55_73 bitb_55_73 gnd C_bl
Rb_55_74 bit_55_74 bit_55_75 R_bl
Rbb_55_74 bitb_55_74 bitb_55_75 R_bl
Cb_55_74 bit_55_74 gnd C_bl
Cbb_55_74 bitb_55_74 gnd C_bl
Rb_55_75 bit_55_75 bit_55_76 R_bl
Rbb_55_75 bitb_55_75 bitb_55_76 R_bl
Cb_55_75 bit_55_75 gnd C_bl
Cbb_55_75 bitb_55_75 gnd C_bl
Rb_55_76 bit_55_76 bit_55_77 R_bl
Rbb_55_76 bitb_55_76 bitb_55_77 R_bl
Cb_55_76 bit_55_76 gnd C_bl
Cbb_55_76 bitb_55_76 gnd C_bl
Rb_55_77 bit_55_77 bit_55_78 R_bl
Rbb_55_77 bitb_55_77 bitb_55_78 R_bl
Cb_55_77 bit_55_77 gnd C_bl
Cbb_55_77 bitb_55_77 gnd C_bl
Rb_55_78 bit_55_78 bit_55_79 R_bl
Rbb_55_78 bitb_55_78 bitb_55_79 R_bl
Cb_55_78 bit_55_78 gnd C_bl
Cbb_55_78 bitb_55_78 gnd C_bl
Rb_55_79 bit_55_79 bit_55_80 R_bl
Rbb_55_79 bitb_55_79 bitb_55_80 R_bl
Cb_55_79 bit_55_79 gnd C_bl
Cbb_55_79 bitb_55_79 gnd C_bl
Rb_55_80 bit_55_80 bit_55_81 R_bl
Rbb_55_80 bitb_55_80 bitb_55_81 R_bl
Cb_55_80 bit_55_80 gnd C_bl
Cbb_55_80 bitb_55_80 gnd C_bl
Rb_55_81 bit_55_81 bit_55_82 R_bl
Rbb_55_81 bitb_55_81 bitb_55_82 R_bl
Cb_55_81 bit_55_81 gnd C_bl
Cbb_55_81 bitb_55_81 gnd C_bl
Rb_55_82 bit_55_82 bit_55_83 R_bl
Rbb_55_82 bitb_55_82 bitb_55_83 R_bl
Cb_55_82 bit_55_82 gnd C_bl
Cbb_55_82 bitb_55_82 gnd C_bl
Rb_55_83 bit_55_83 bit_55_84 R_bl
Rbb_55_83 bitb_55_83 bitb_55_84 R_bl
Cb_55_83 bit_55_83 gnd C_bl
Cbb_55_83 bitb_55_83 gnd C_bl
Rb_55_84 bit_55_84 bit_55_85 R_bl
Rbb_55_84 bitb_55_84 bitb_55_85 R_bl
Cb_55_84 bit_55_84 gnd C_bl
Cbb_55_84 bitb_55_84 gnd C_bl
Rb_55_85 bit_55_85 bit_55_86 R_bl
Rbb_55_85 bitb_55_85 bitb_55_86 R_bl
Cb_55_85 bit_55_85 gnd C_bl
Cbb_55_85 bitb_55_85 gnd C_bl
Rb_55_86 bit_55_86 bit_55_87 R_bl
Rbb_55_86 bitb_55_86 bitb_55_87 R_bl
Cb_55_86 bit_55_86 gnd C_bl
Cbb_55_86 bitb_55_86 gnd C_bl
Rb_55_87 bit_55_87 bit_55_88 R_bl
Rbb_55_87 bitb_55_87 bitb_55_88 R_bl
Cb_55_87 bit_55_87 gnd C_bl
Cbb_55_87 bitb_55_87 gnd C_bl
Rb_55_88 bit_55_88 bit_55_89 R_bl
Rbb_55_88 bitb_55_88 bitb_55_89 R_bl
Cb_55_88 bit_55_88 gnd C_bl
Cbb_55_88 bitb_55_88 gnd C_bl
Rb_55_89 bit_55_89 bit_55_90 R_bl
Rbb_55_89 bitb_55_89 bitb_55_90 R_bl
Cb_55_89 bit_55_89 gnd C_bl
Cbb_55_89 bitb_55_89 gnd C_bl
Rb_55_90 bit_55_90 bit_55_91 R_bl
Rbb_55_90 bitb_55_90 bitb_55_91 R_bl
Cb_55_90 bit_55_90 gnd C_bl
Cbb_55_90 bitb_55_90 gnd C_bl
Rb_55_91 bit_55_91 bit_55_92 R_bl
Rbb_55_91 bitb_55_91 bitb_55_92 R_bl
Cb_55_91 bit_55_91 gnd C_bl
Cbb_55_91 bitb_55_91 gnd C_bl
Rb_55_92 bit_55_92 bit_55_93 R_bl
Rbb_55_92 bitb_55_92 bitb_55_93 R_bl
Cb_55_92 bit_55_92 gnd C_bl
Cbb_55_92 bitb_55_92 gnd C_bl
Rb_55_93 bit_55_93 bit_55_94 R_bl
Rbb_55_93 bitb_55_93 bitb_55_94 R_bl
Cb_55_93 bit_55_93 gnd C_bl
Cbb_55_93 bitb_55_93 gnd C_bl
Rb_55_94 bit_55_94 bit_55_95 R_bl
Rbb_55_94 bitb_55_94 bitb_55_95 R_bl
Cb_55_94 bit_55_94 gnd C_bl
Cbb_55_94 bitb_55_94 gnd C_bl
Rb_55_95 bit_55_95 bit_55_96 R_bl
Rbb_55_95 bitb_55_95 bitb_55_96 R_bl
Cb_55_95 bit_55_95 gnd C_bl
Cbb_55_95 bitb_55_95 gnd C_bl
Rb_55_96 bit_55_96 bit_55_97 R_bl
Rbb_55_96 bitb_55_96 bitb_55_97 R_bl
Cb_55_96 bit_55_96 gnd C_bl
Cbb_55_96 bitb_55_96 gnd C_bl
Rb_55_97 bit_55_97 bit_55_98 R_bl
Rbb_55_97 bitb_55_97 bitb_55_98 R_bl
Cb_55_97 bit_55_97 gnd C_bl
Cbb_55_97 bitb_55_97 gnd C_bl
Rb_55_98 bit_55_98 bit_55_99 R_bl
Rbb_55_98 bitb_55_98 bitb_55_99 R_bl
Cb_55_98 bit_55_98 gnd C_bl
Cbb_55_98 bitb_55_98 gnd C_bl
Rb_55_99 bit_55_99 bit_55_100 R_bl
Rbb_55_99 bitb_55_99 bitb_55_100 R_bl
Cb_55_99 bit_55_99 gnd C_bl
Cbb_55_99 bitb_55_99 gnd C_bl
Rb_56_0 bit_56_0 bit_56_1 R_bl
Rbb_56_0 bitb_56_0 bitb_56_1 R_bl
Cb_56_0 bit_56_0 gnd C_bl
Cbb_56_0 bitb_56_0 gnd C_bl
Rb_56_1 bit_56_1 bit_56_2 R_bl
Rbb_56_1 bitb_56_1 bitb_56_2 R_bl
Cb_56_1 bit_56_1 gnd C_bl
Cbb_56_1 bitb_56_1 gnd C_bl
Rb_56_2 bit_56_2 bit_56_3 R_bl
Rbb_56_2 bitb_56_2 bitb_56_3 R_bl
Cb_56_2 bit_56_2 gnd C_bl
Cbb_56_2 bitb_56_2 gnd C_bl
Rb_56_3 bit_56_3 bit_56_4 R_bl
Rbb_56_3 bitb_56_3 bitb_56_4 R_bl
Cb_56_3 bit_56_3 gnd C_bl
Cbb_56_3 bitb_56_3 gnd C_bl
Rb_56_4 bit_56_4 bit_56_5 R_bl
Rbb_56_4 bitb_56_4 bitb_56_5 R_bl
Cb_56_4 bit_56_4 gnd C_bl
Cbb_56_4 bitb_56_4 gnd C_bl
Rb_56_5 bit_56_5 bit_56_6 R_bl
Rbb_56_5 bitb_56_5 bitb_56_6 R_bl
Cb_56_5 bit_56_5 gnd C_bl
Cbb_56_5 bitb_56_5 gnd C_bl
Rb_56_6 bit_56_6 bit_56_7 R_bl
Rbb_56_6 bitb_56_6 bitb_56_7 R_bl
Cb_56_6 bit_56_6 gnd C_bl
Cbb_56_6 bitb_56_6 gnd C_bl
Rb_56_7 bit_56_7 bit_56_8 R_bl
Rbb_56_7 bitb_56_7 bitb_56_8 R_bl
Cb_56_7 bit_56_7 gnd C_bl
Cbb_56_7 bitb_56_7 gnd C_bl
Rb_56_8 bit_56_8 bit_56_9 R_bl
Rbb_56_8 bitb_56_8 bitb_56_9 R_bl
Cb_56_8 bit_56_8 gnd C_bl
Cbb_56_8 bitb_56_8 gnd C_bl
Rb_56_9 bit_56_9 bit_56_10 R_bl
Rbb_56_9 bitb_56_9 bitb_56_10 R_bl
Cb_56_9 bit_56_9 gnd C_bl
Cbb_56_9 bitb_56_9 gnd C_bl
Rb_56_10 bit_56_10 bit_56_11 R_bl
Rbb_56_10 bitb_56_10 bitb_56_11 R_bl
Cb_56_10 bit_56_10 gnd C_bl
Cbb_56_10 bitb_56_10 gnd C_bl
Rb_56_11 bit_56_11 bit_56_12 R_bl
Rbb_56_11 bitb_56_11 bitb_56_12 R_bl
Cb_56_11 bit_56_11 gnd C_bl
Cbb_56_11 bitb_56_11 gnd C_bl
Rb_56_12 bit_56_12 bit_56_13 R_bl
Rbb_56_12 bitb_56_12 bitb_56_13 R_bl
Cb_56_12 bit_56_12 gnd C_bl
Cbb_56_12 bitb_56_12 gnd C_bl
Rb_56_13 bit_56_13 bit_56_14 R_bl
Rbb_56_13 bitb_56_13 bitb_56_14 R_bl
Cb_56_13 bit_56_13 gnd C_bl
Cbb_56_13 bitb_56_13 gnd C_bl
Rb_56_14 bit_56_14 bit_56_15 R_bl
Rbb_56_14 bitb_56_14 bitb_56_15 R_bl
Cb_56_14 bit_56_14 gnd C_bl
Cbb_56_14 bitb_56_14 gnd C_bl
Rb_56_15 bit_56_15 bit_56_16 R_bl
Rbb_56_15 bitb_56_15 bitb_56_16 R_bl
Cb_56_15 bit_56_15 gnd C_bl
Cbb_56_15 bitb_56_15 gnd C_bl
Rb_56_16 bit_56_16 bit_56_17 R_bl
Rbb_56_16 bitb_56_16 bitb_56_17 R_bl
Cb_56_16 bit_56_16 gnd C_bl
Cbb_56_16 bitb_56_16 gnd C_bl
Rb_56_17 bit_56_17 bit_56_18 R_bl
Rbb_56_17 bitb_56_17 bitb_56_18 R_bl
Cb_56_17 bit_56_17 gnd C_bl
Cbb_56_17 bitb_56_17 gnd C_bl
Rb_56_18 bit_56_18 bit_56_19 R_bl
Rbb_56_18 bitb_56_18 bitb_56_19 R_bl
Cb_56_18 bit_56_18 gnd C_bl
Cbb_56_18 bitb_56_18 gnd C_bl
Rb_56_19 bit_56_19 bit_56_20 R_bl
Rbb_56_19 bitb_56_19 bitb_56_20 R_bl
Cb_56_19 bit_56_19 gnd C_bl
Cbb_56_19 bitb_56_19 gnd C_bl
Rb_56_20 bit_56_20 bit_56_21 R_bl
Rbb_56_20 bitb_56_20 bitb_56_21 R_bl
Cb_56_20 bit_56_20 gnd C_bl
Cbb_56_20 bitb_56_20 gnd C_bl
Rb_56_21 bit_56_21 bit_56_22 R_bl
Rbb_56_21 bitb_56_21 bitb_56_22 R_bl
Cb_56_21 bit_56_21 gnd C_bl
Cbb_56_21 bitb_56_21 gnd C_bl
Rb_56_22 bit_56_22 bit_56_23 R_bl
Rbb_56_22 bitb_56_22 bitb_56_23 R_bl
Cb_56_22 bit_56_22 gnd C_bl
Cbb_56_22 bitb_56_22 gnd C_bl
Rb_56_23 bit_56_23 bit_56_24 R_bl
Rbb_56_23 bitb_56_23 bitb_56_24 R_bl
Cb_56_23 bit_56_23 gnd C_bl
Cbb_56_23 bitb_56_23 gnd C_bl
Rb_56_24 bit_56_24 bit_56_25 R_bl
Rbb_56_24 bitb_56_24 bitb_56_25 R_bl
Cb_56_24 bit_56_24 gnd C_bl
Cbb_56_24 bitb_56_24 gnd C_bl
Rb_56_25 bit_56_25 bit_56_26 R_bl
Rbb_56_25 bitb_56_25 bitb_56_26 R_bl
Cb_56_25 bit_56_25 gnd C_bl
Cbb_56_25 bitb_56_25 gnd C_bl
Rb_56_26 bit_56_26 bit_56_27 R_bl
Rbb_56_26 bitb_56_26 bitb_56_27 R_bl
Cb_56_26 bit_56_26 gnd C_bl
Cbb_56_26 bitb_56_26 gnd C_bl
Rb_56_27 bit_56_27 bit_56_28 R_bl
Rbb_56_27 bitb_56_27 bitb_56_28 R_bl
Cb_56_27 bit_56_27 gnd C_bl
Cbb_56_27 bitb_56_27 gnd C_bl
Rb_56_28 bit_56_28 bit_56_29 R_bl
Rbb_56_28 bitb_56_28 bitb_56_29 R_bl
Cb_56_28 bit_56_28 gnd C_bl
Cbb_56_28 bitb_56_28 gnd C_bl
Rb_56_29 bit_56_29 bit_56_30 R_bl
Rbb_56_29 bitb_56_29 bitb_56_30 R_bl
Cb_56_29 bit_56_29 gnd C_bl
Cbb_56_29 bitb_56_29 gnd C_bl
Rb_56_30 bit_56_30 bit_56_31 R_bl
Rbb_56_30 bitb_56_30 bitb_56_31 R_bl
Cb_56_30 bit_56_30 gnd C_bl
Cbb_56_30 bitb_56_30 gnd C_bl
Rb_56_31 bit_56_31 bit_56_32 R_bl
Rbb_56_31 bitb_56_31 bitb_56_32 R_bl
Cb_56_31 bit_56_31 gnd C_bl
Cbb_56_31 bitb_56_31 gnd C_bl
Rb_56_32 bit_56_32 bit_56_33 R_bl
Rbb_56_32 bitb_56_32 bitb_56_33 R_bl
Cb_56_32 bit_56_32 gnd C_bl
Cbb_56_32 bitb_56_32 gnd C_bl
Rb_56_33 bit_56_33 bit_56_34 R_bl
Rbb_56_33 bitb_56_33 bitb_56_34 R_bl
Cb_56_33 bit_56_33 gnd C_bl
Cbb_56_33 bitb_56_33 gnd C_bl
Rb_56_34 bit_56_34 bit_56_35 R_bl
Rbb_56_34 bitb_56_34 bitb_56_35 R_bl
Cb_56_34 bit_56_34 gnd C_bl
Cbb_56_34 bitb_56_34 gnd C_bl
Rb_56_35 bit_56_35 bit_56_36 R_bl
Rbb_56_35 bitb_56_35 bitb_56_36 R_bl
Cb_56_35 bit_56_35 gnd C_bl
Cbb_56_35 bitb_56_35 gnd C_bl
Rb_56_36 bit_56_36 bit_56_37 R_bl
Rbb_56_36 bitb_56_36 bitb_56_37 R_bl
Cb_56_36 bit_56_36 gnd C_bl
Cbb_56_36 bitb_56_36 gnd C_bl
Rb_56_37 bit_56_37 bit_56_38 R_bl
Rbb_56_37 bitb_56_37 bitb_56_38 R_bl
Cb_56_37 bit_56_37 gnd C_bl
Cbb_56_37 bitb_56_37 gnd C_bl
Rb_56_38 bit_56_38 bit_56_39 R_bl
Rbb_56_38 bitb_56_38 bitb_56_39 R_bl
Cb_56_38 bit_56_38 gnd C_bl
Cbb_56_38 bitb_56_38 gnd C_bl
Rb_56_39 bit_56_39 bit_56_40 R_bl
Rbb_56_39 bitb_56_39 bitb_56_40 R_bl
Cb_56_39 bit_56_39 gnd C_bl
Cbb_56_39 bitb_56_39 gnd C_bl
Rb_56_40 bit_56_40 bit_56_41 R_bl
Rbb_56_40 bitb_56_40 bitb_56_41 R_bl
Cb_56_40 bit_56_40 gnd C_bl
Cbb_56_40 bitb_56_40 gnd C_bl
Rb_56_41 bit_56_41 bit_56_42 R_bl
Rbb_56_41 bitb_56_41 bitb_56_42 R_bl
Cb_56_41 bit_56_41 gnd C_bl
Cbb_56_41 bitb_56_41 gnd C_bl
Rb_56_42 bit_56_42 bit_56_43 R_bl
Rbb_56_42 bitb_56_42 bitb_56_43 R_bl
Cb_56_42 bit_56_42 gnd C_bl
Cbb_56_42 bitb_56_42 gnd C_bl
Rb_56_43 bit_56_43 bit_56_44 R_bl
Rbb_56_43 bitb_56_43 bitb_56_44 R_bl
Cb_56_43 bit_56_43 gnd C_bl
Cbb_56_43 bitb_56_43 gnd C_bl
Rb_56_44 bit_56_44 bit_56_45 R_bl
Rbb_56_44 bitb_56_44 bitb_56_45 R_bl
Cb_56_44 bit_56_44 gnd C_bl
Cbb_56_44 bitb_56_44 gnd C_bl
Rb_56_45 bit_56_45 bit_56_46 R_bl
Rbb_56_45 bitb_56_45 bitb_56_46 R_bl
Cb_56_45 bit_56_45 gnd C_bl
Cbb_56_45 bitb_56_45 gnd C_bl
Rb_56_46 bit_56_46 bit_56_47 R_bl
Rbb_56_46 bitb_56_46 bitb_56_47 R_bl
Cb_56_46 bit_56_46 gnd C_bl
Cbb_56_46 bitb_56_46 gnd C_bl
Rb_56_47 bit_56_47 bit_56_48 R_bl
Rbb_56_47 bitb_56_47 bitb_56_48 R_bl
Cb_56_47 bit_56_47 gnd C_bl
Cbb_56_47 bitb_56_47 gnd C_bl
Rb_56_48 bit_56_48 bit_56_49 R_bl
Rbb_56_48 bitb_56_48 bitb_56_49 R_bl
Cb_56_48 bit_56_48 gnd C_bl
Cbb_56_48 bitb_56_48 gnd C_bl
Rb_56_49 bit_56_49 bit_56_50 R_bl
Rbb_56_49 bitb_56_49 bitb_56_50 R_bl
Cb_56_49 bit_56_49 gnd C_bl
Cbb_56_49 bitb_56_49 gnd C_bl
Rb_56_50 bit_56_50 bit_56_51 R_bl
Rbb_56_50 bitb_56_50 bitb_56_51 R_bl
Cb_56_50 bit_56_50 gnd C_bl
Cbb_56_50 bitb_56_50 gnd C_bl
Rb_56_51 bit_56_51 bit_56_52 R_bl
Rbb_56_51 bitb_56_51 bitb_56_52 R_bl
Cb_56_51 bit_56_51 gnd C_bl
Cbb_56_51 bitb_56_51 gnd C_bl
Rb_56_52 bit_56_52 bit_56_53 R_bl
Rbb_56_52 bitb_56_52 bitb_56_53 R_bl
Cb_56_52 bit_56_52 gnd C_bl
Cbb_56_52 bitb_56_52 gnd C_bl
Rb_56_53 bit_56_53 bit_56_54 R_bl
Rbb_56_53 bitb_56_53 bitb_56_54 R_bl
Cb_56_53 bit_56_53 gnd C_bl
Cbb_56_53 bitb_56_53 gnd C_bl
Rb_56_54 bit_56_54 bit_56_55 R_bl
Rbb_56_54 bitb_56_54 bitb_56_55 R_bl
Cb_56_54 bit_56_54 gnd C_bl
Cbb_56_54 bitb_56_54 gnd C_bl
Rb_56_55 bit_56_55 bit_56_56 R_bl
Rbb_56_55 bitb_56_55 bitb_56_56 R_bl
Cb_56_55 bit_56_55 gnd C_bl
Cbb_56_55 bitb_56_55 gnd C_bl
Rb_56_56 bit_56_56 bit_56_57 R_bl
Rbb_56_56 bitb_56_56 bitb_56_57 R_bl
Cb_56_56 bit_56_56 gnd C_bl
Cbb_56_56 bitb_56_56 gnd C_bl
Rb_56_57 bit_56_57 bit_56_58 R_bl
Rbb_56_57 bitb_56_57 bitb_56_58 R_bl
Cb_56_57 bit_56_57 gnd C_bl
Cbb_56_57 bitb_56_57 gnd C_bl
Rb_56_58 bit_56_58 bit_56_59 R_bl
Rbb_56_58 bitb_56_58 bitb_56_59 R_bl
Cb_56_58 bit_56_58 gnd C_bl
Cbb_56_58 bitb_56_58 gnd C_bl
Rb_56_59 bit_56_59 bit_56_60 R_bl
Rbb_56_59 bitb_56_59 bitb_56_60 R_bl
Cb_56_59 bit_56_59 gnd C_bl
Cbb_56_59 bitb_56_59 gnd C_bl
Rb_56_60 bit_56_60 bit_56_61 R_bl
Rbb_56_60 bitb_56_60 bitb_56_61 R_bl
Cb_56_60 bit_56_60 gnd C_bl
Cbb_56_60 bitb_56_60 gnd C_bl
Rb_56_61 bit_56_61 bit_56_62 R_bl
Rbb_56_61 bitb_56_61 bitb_56_62 R_bl
Cb_56_61 bit_56_61 gnd C_bl
Cbb_56_61 bitb_56_61 gnd C_bl
Rb_56_62 bit_56_62 bit_56_63 R_bl
Rbb_56_62 bitb_56_62 bitb_56_63 R_bl
Cb_56_62 bit_56_62 gnd C_bl
Cbb_56_62 bitb_56_62 gnd C_bl
Rb_56_63 bit_56_63 bit_56_64 R_bl
Rbb_56_63 bitb_56_63 bitb_56_64 R_bl
Cb_56_63 bit_56_63 gnd C_bl
Cbb_56_63 bitb_56_63 gnd C_bl
Rb_56_64 bit_56_64 bit_56_65 R_bl
Rbb_56_64 bitb_56_64 bitb_56_65 R_bl
Cb_56_64 bit_56_64 gnd C_bl
Cbb_56_64 bitb_56_64 gnd C_bl
Rb_56_65 bit_56_65 bit_56_66 R_bl
Rbb_56_65 bitb_56_65 bitb_56_66 R_bl
Cb_56_65 bit_56_65 gnd C_bl
Cbb_56_65 bitb_56_65 gnd C_bl
Rb_56_66 bit_56_66 bit_56_67 R_bl
Rbb_56_66 bitb_56_66 bitb_56_67 R_bl
Cb_56_66 bit_56_66 gnd C_bl
Cbb_56_66 bitb_56_66 gnd C_bl
Rb_56_67 bit_56_67 bit_56_68 R_bl
Rbb_56_67 bitb_56_67 bitb_56_68 R_bl
Cb_56_67 bit_56_67 gnd C_bl
Cbb_56_67 bitb_56_67 gnd C_bl
Rb_56_68 bit_56_68 bit_56_69 R_bl
Rbb_56_68 bitb_56_68 bitb_56_69 R_bl
Cb_56_68 bit_56_68 gnd C_bl
Cbb_56_68 bitb_56_68 gnd C_bl
Rb_56_69 bit_56_69 bit_56_70 R_bl
Rbb_56_69 bitb_56_69 bitb_56_70 R_bl
Cb_56_69 bit_56_69 gnd C_bl
Cbb_56_69 bitb_56_69 gnd C_bl
Rb_56_70 bit_56_70 bit_56_71 R_bl
Rbb_56_70 bitb_56_70 bitb_56_71 R_bl
Cb_56_70 bit_56_70 gnd C_bl
Cbb_56_70 bitb_56_70 gnd C_bl
Rb_56_71 bit_56_71 bit_56_72 R_bl
Rbb_56_71 bitb_56_71 bitb_56_72 R_bl
Cb_56_71 bit_56_71 gnd C_bl
Cbb_56_71 bitb_56_71 gnd C_bl
Rb_56_72 bit_56_72 bit_56_73 R_bl
Rbb_56_72 bitb_56_72 bitb_56_73 R_bl
Cb_56_72 bit_56_72 gnd C_bl
Cbb_56_72 bitb_56_72 gnd C_bl
Rb_56_73 bit_56_73 bit_56_74 R_bl
Rbb_56_73 bitb_56_73 bitb_56_74 R_bl
Cb_56_73 bit_56_73 gnd C_bl
Cbb_56_73 bitb_56_73 gnd C_bl
Rb_56_74 bit_56_74 bit_56_75 R_bl
Rbb_56_74 bitb_56_74 bitb_56_75 R_bl
Cb_56_74 bit_56_74 gnd C_bl
Cbb_56_74 bitb_56_74 gnd C_bl
Rb_56_75 bit_56_75 bit_56_76 R_bl
Rbb_56_75 bitb_56_75 bitb_56_76 R_bl
Cb_56_75 bit_56_75 gnd C_bl
Cbb_56_75 bitb_56_75 gnd C_bl
Rb_56_76 bit_56_76 bit_56_77 R_bl
Rbb_56_76 bitb_56_76 bitb_56_77 R_bl
Cb_56_76 bit_56_76 gnd C_bl
Cbb_56_76 bitb_56_76 gnd C_bl
Rb_56_77 bit_56_77 bit_56_78 R_bl
Rbb_56_77 bitb_56_77 bitb_56_78 R_bl
Cb_56_77 bit_56_77 gnd C_bl
Cbb_56_77 bitb_56_77 gnd C_bl
Rb_56_78 bit_56_78 bit_56_79 R_bl
Rbb_56_78 bitb_56_78 bitb_56_79 R_bl
Cb_56_78 bit_56_78 gnd C_bl
Cbb_56_78 bitb_56_78 gnd C_bl
Rb_56_79 bit_56_79 bit_56_80 R_bl
Rbb_56_79 bitb_56_79 bitb_56_80 R_bl
Cb_56_79 bit_56_79 gnd C_bl
Cbb_56_79 bitb_56_79 gnd C_bl
Rb_56_80 bit_56_80 bit_56_81 R_bl
Rbb_56_80 bitb_56_80 bitb_56_81 R_bl
Cb_56_80 bit_56_80 gnd C_bl
Cbb_56_80 bitb_56_80 gnd C_bl
Rb_56_81 bit_56_81 bit_56_82 R_bl
Rbb_56_81 bitb_56_81 bitb_56_82 R_bl
Cb_56_81 bit_56_81 gnd C_bl
Cbb_56_81 bitb_56_81 gnd C_bl
Rb_56_82 bit_56_82 bit_56_83 R_bl
Rbb_56_82 bitb_56_82 bitb_56_83 R_bl
Cb_56_82 bit_56_82 gnd C_bl
Cbb_56_82 bitb_56_82 gnd C_bl
Rb_56_83 bit_56_83 bit_56_84 R_bl
Rbb_56_83 bitb_56_83 bitb_56_84 R_bl
Cb_56_83 bit_56_83 gnd C_bl
Cbb_56_83 bitb_56_83 gnd C_bl
Rb_56_84 bit_56_84 bit_56_85 R_bl
Rbb_56_84 bitb_56_84 bitb_56_85 R_bl
Cb_56_84 bit_56_84 gnd C_bl
Cbb_56_84 bitb_56_84 gnd C_bl
Rb_56_85 bit_56_85 bit_56_86 R_bl
Rbb_56_85 bitb_56_85 bitb_56_86 R_bl
Cb_56_85 bit_56_85 gnd C_bl
Cbb_56_85 bitb_56_85 gnd C_bl
Rb_56_86 bit_56_86 bit_56_87 R_bl
Rbb_56_86 bitb_56_86 bitb_56_87 R_bl
Cb_56_86 bit_56_86 gnd C_bl
Cbb_56_86 bitb_56_86 gnd C_bl
Rb_56_87 bit_56_87 bit_56_88 R_bl
Rbb_56_87 bitb_56_87 bitb_56_88 R_bl
Cb_56_87 bit_56_87 gnd C_bl
Cbb_56_87 bitb_56_87 gnd C_bl
Rb_56_88 bit_56_88 bit_56_89 R_bl
Rbb_56_88 bitb_56_88 bitb_56_89 R_bl
Cb_56_88 bit_56_88 gnd C_bl
Cbb_56_88 bitb_56_88 gnd C_bl
Rb_56_89 bit_56_89 bit_56_90 R_bl
Rbb_56_89 bitb_56_89 bitb_56_90 R_bl
Cb_56_89 bit_56_89 gnd C_bl
Cbb_56_89 bitb_56_89 gnd C_bl
Rb_56_90 bit_56_90 bit_56_91 R_bl
Rbb_56_90 bitb_56_90 bitb_56_91 R_bl
Cb_56_90 bit_56_90 gnd C_bl
Cbb_56_90 bitb_56_90 gnd C_bl
Rb_56_91 bit_56_91 bit_56_92 R_bl
Rbb_56_91 bitb_56_91 bitb_56_92 R_bl
Cb_56_91 bit_56_91 gnd C_bl
Cbb_56_91 bitb_56_91 gnd C_bl
Rb_56_92 bit_56_92 bit_56_93 R_bl
Rbb_56_92 bitb_56_92 bitb_56_93 R_bl
Cb_56_92 bit_56_92 gnd C_bl
Cbb_56_92 bitb_56_92 gnd C_bl
Rb_56_93 bit_56_93 bit_56_94 R_bl
Rbb_56_93 bitb_56_93 bitb_56_94 R_bl
Cb_56_93 bit_56_93 gnd C_bl
Cbb_56_93 bitb_56_93 gnd C_bl
Rb_56_94 bit_56_94 bit_56_95 R_bl
Rbb_56_94 bitb_56_94 bitb_56_95 R_bl
Cb_56_94 bit_56_94 gnd C_bl
Cbb_56_94 bitb_56_94 gnd C_bl
Rb_56_95 bit_56_95 bit_56_96 R_bl
Rbb_56_95 bitb_56_95 bitb_56_96 R_bl
Cb_56_95 bit_56_95 gnd C_bl
Cbb_56_95 bitb_56_95 gnd C_bl
Rb_56_96 bit_56_96 bit_56_97 R_bl
Rbb_56_96 bitb_56_96 bitb_56_97 R_bl
Cb_56_96 bit_56_96 gnd C_bl
Cbb_56_96 bitb_56_96 gnd C_bl
Rb_56_97 bit_56_97 bit_56_98 R_bl
Rbb_56_97 bitb_56_97 bitb_56_98 R_bl
Cb_56_97 bit_56_97 gnd C_bl
Cbb_56_97 bitb_56_97 gnd C_bl
Rb_56_98 bit_56_98 bit_56_99 R_bl
Rbb_56_98 bitb_56_98 bitb_56_99 R_bl
Cb_56_98 bit_56_98 gnd C_bl
Cbb_56_98 bitb_56_98 gnd C_bl
Rb_56_99 bit_56_99 bit_56_100 R_bl
Rbb_56_99 bitb_56_99 bitb_56_100 R_bl
Cb_56_99 bit_56_99 gnd C_bl
Cbb_56_99 bitb_56_99 gnd C_bl
Rb_57_0 bit_57_0 bit_57_1 R_bl
Rbb_57_0 bitb_57_0 bitb_57_1 R_bl
Cb_57_0 bit_57_0 gnd C_bl
Cbb_57_0 bitb_57_0 gnd C_bl
Rb_57_1 bit_57_1 bit_57_2 R_bl
Rbb_57_1 bitb_57_1 bitb_57_2 R_bl
Cb_57_1 bit_57_1 gnd C_bl
Cbb_57_1 bitb_57_1 gnd C_bl
Rb_57_2 bit_57_2 bit_57_3 R_bl
Rbb_57_2 bitb_57_2 bitb_57_3 R_bl
Cb_57_2 bit_57_2 gnd C_bl
Cbb_57_2 bitb_57_2 gnd C_bl
Rb_57_3 bit_57_3 bit_57_4 R_bl
Rbb_57_3 bitb_57_3 bitb_57_4 R_bl
Cb_57_3 bit_57_3 gnd C_bl
Cbb_57_3 bitb_57_3 gnd C_bl
Rb_57_4 bit_57_4 bit_57_5 R_bl
Rbb_57_4 bitb_57_4 bitb_57_5 R_bl
Cb_57_4 bit_57_4 gnd C_bl
Cbb_57_4 bitb_57_4 gnd C_bl
Rb_57_5 bit_57_5 bit_57_6 R_bl
Rbb_57_5 bitb_57_5 bitb_57_6 R_bl
Cb_57_5 bit_57_5 gnd C_bl
Cbb_57_5 bitb_57_5 gnd C_bl
Rb_57_6 bit_57_6 bit_57_7 R_bl
Rbb_57_6 bitb_57_6 bitb_57_7 R_bl
Cb_57_6 bit_57_6 gnd C_bl
Cbb_57_6 bitb_57_6 gnd C_bl
Rb_57_7 bit_57_7 bit_57_8 R_bl
Rbb_57_7 bitb_57_7 bitb_57_8 R_bl
Cb_57_7 bit_57_7 gnd C_bl
Cbb_57_7 bitb_57_7 gnd C_bl
Rb_57_8 bit_57_8 bit_57_9 R_bl
Rbb_57_8 bitb_57_8 bitb_57_9 R_bl
Cb_57_8 bit_57_8 gnd C_bl
Cbb_57_8 bitb_57_8 gnd C_bl
Rb_57_9 bit_57_9 bit_57_10 R_bl
Rbb_57_9 bitb_57_9 bitb_57_10 R_bl
Cb_57_9 bit_57_9 gnd C_bl
Cbb_57_9 bitb_57_9 gnd C_bl
Rb_57_10 bit_57_10 bit_57_11 R_bl
Rbb_57_10 bitb_57_10 bitb_57_11 R_bl
Cb_57_10 bit_57_10 gnd C_bl
Cbb_57_10 bitb_57_10 gnd C_bl
Rb_57_11 bit_57_11 bit_57_12 R_bl
Rbb_57_11 bitb_57_11 bitb_57_12 R_bl
Cb_57_11 bit_57_11 gnd C_bl
Cbb_57_11 bitb_57_11 gnd C_bl
Rb_57_12 bit_57_12 bit_57_13 R_bl
Rbb_57_12 bitb_57_12 bitb_57_13 R_bl
Cb_57_12 bit_57_12 gnd C_bl
Cbb_57_12 bitb_57_12 gnd C_bl
Rb_57_13 bit_57_13 bit_57_14 R_bl
Rbb_57_13 bitb_57_13 bitb_57_14 R_bl
Cb_57_13 bit_57_13 gnd C_bl
Cbb_57_13 bitb_57_13 gnd C_bl
Rb_57_14 bit_57_14 bit_57_15 R_bl
Rbb_57_14 bitb_57_14 bitb_57_15 R_bl
Cb_57_14 bit_57_14 gnd C_bl
Cbb_57_14 bitb_57_14 gnd C_bl
Rb_57_15 bit_57_15 bit_57_16 R_bl
Rbb_57_15 bitb_57_15 bitb_57_16 R_bl
Cb_57_15 bit_57_15 gnd C_bl
Cbb_57_15 bitb_57_15 gnd C_bl
Rb_57_16 bit_57_16 bit_57_17 R_bl
Rbb_57_16 bitb_57_16 bitb_57_17 R_bl
Cb_57_16 bit_57_16 gnd C_bl
Cbb_57_16 bitb_57_16 gnd C_bl
Rb_57_17 bit_57_17 bit_57_18 R_bl
Rbb_57_17 bitb_57_17 bitb_57_18 R_bl
Cb_57_17 bit_57_17 gnd C_bl
Cbb_57_17 bitb_57_17 gnd C_bl
Rb_57_18 bit_57_18 bit_57_19 R_bl
Rbb_57_18 bitb_57_18 bitb_57_19 R_bl
Cb_57_18 bit_57_18 gnd C_bl
Cbb_57_18 bitb_57_18 gnd C_bl
Rb_57_19 bit_57_19 bit_57_20 R_bl
Rbb_57_19 bitb_57_19 bitb_57_20 R_bl
Cb_57_19 bit_57_19 gnd C_bl
Cbb_57_19 bitb_57_19 gnd C_bl
Rb_57_20 bit_57_20 bit_57_21 R_bl
Rbb_57_20 bitb_57_20 bitb_57_21 R_bl
Cb_57_20 bit_57_20 gnd C_bl
Cbb_57_20 bitb_57_20 gnd C_bl
Rb_57_21 bit_57_21 bit_57_22 R_bl
Rbb_57_21 bitb_57_21 bitb_57_22 R_bl
Cb_57_21 bit_57_21 gnd C_bl
Cbb_57_21 bitb_57_21 gnd C_bl
Rb_57_22 bit_57_22 bit_57_23 R_bl
Rbb_57_22 bitb_57_22 bitb_57_23 R_bl
Cb_57_22 bit_57_22 gnd C_bl
Cbb_57_22 bitb_57_22 gnd C_bl
Rb_57_23 bit_57_23 bit_57_24 R_bl
Rbb_57_23 bitb_57_23 bitb_57_24 R_bl
Cb_57_23 bit_57_23 gnd C_bl
Cbb_57_23 bitb_57_23 gnd C_bl
Rb_57_24 bit_57_24 bit_57_25 R_bl
Rbb_57_24 bitb_57_24 bitb_57_25 R_bl
Cb_57_24 bit_57_24 gnd C_bl
Cbb_57_24 bitb_57_24 gnd C_bl
Rb_57_25 bit_57_25 bit_57_26 R_bl
Rbb_57_25 bitb_57_25 bitb_57_26 R_bl
Cb_57_25 bit_57_25 gnd C_bl
Cbb_57_25 bitb_57_25 gnd C_bl
Rb_57_26 bit_57_26 bit_57_27 R_bl
Rbb_57_26 bitb_57_26 bitb_57_27 R_bl
Cb_57_26 bit_57_26 gnd C_bl
Cbb_57_26 bitb_57_26 gnd C_bl
Rb_57_27 bit_57_27 bit_57_28 R_bl
Rbb_57_27 bitb_57_27 bitb_57_28 R_bl
Cb_57_27 bit_57_27 gnd C_bl
Cbb_57_27 bitb_57_27 gnd C_bl
Rb_57_28 bit_57_28 bit_57_29 R_bl
Rbb_57_28 bitb_57_28 bitb_57_29 R_bl
Cb_57_28 bit_57_28 gnd C_bl
Cbb_57_28 bitb_57_28 gnd C_bl
Rb_57_29 bit_57_29 bit_57_30 R_bl
Rbb_57_29 bitb_57_29 bitb_57_30 R_bl
Cb_57_29 bit_57_29 gnd C_bl
Cbb_57_29 bitb_57_29 gnd C_bl
Rb_57_30 bit_57_30 bit_57_31 R_bl
Rbb_57_30 bitb_57_30 bitb_57_31 R_bl
Cb_57_30 bit_57_30 gnd C_bl
Cbb_57_30 bitb_57_30 gnd C_bl
Rb_57_31 bit_57_31 bit_57_32 R_bl
Rbb_57_31 bitb_57_31 bitb_57_32 R_bl
Cb_57_31 bit_57_31 gnd C_bl
Cbb_57_31 bitb_57_31 gnd C_bl
Rb_57_32 bit_57_32 bit_57_33 R_bl
Rbb_57_32 bitb_57_32 bitb_57_33 R_bl
Cb_57_32 bit_57_32 gnd C_bl
Cbb_57_32 bitb_57_32 gnd C_bl
Rb_57_33 bit_57_33 bit_57_34 R_bl
Rbb_57_33 bitb_57_33 bitb_57_34 R_bl
Cb_57_33 bit_57_33 gnd C_bl
Cbb_57_33 bitb_57_33 gnd C_bl
Rb_57_34 bit_57_34 bit_57_35 R_bl
Rbb_57_34 bitb_57_34 bitb_57_35 R_bl
Cb_57_34 bit_57_34 gnd C_bl
Cbb_57_34 bitb_57_34 gnd C_bl
Rb_57_35 bit_57_35 bit_57_36 R_bl
Rbb_57_35 bitb_57_35 bitb_57_36 R_bl
Cb_57_35 bit_57_35 gnd C_bl
Cbb_57_35 bitb_57_35 gnd C_bl
Rb_57_36 bit_57_36 bit_57_37 R_bl
Rbb_57_36 bitb_57_36 bitb_57_37 R_bl
Cb_57_36 bit_57_36 gnd C_bl
Cbb_57_36 bitb_57_36 gnd C_bl
Rb_57_37 bit_57_37 bit_57_38 R_bl
Rbb_57_37 bitb_57_37 bitb_57_38 R_bl
Cb_57_37 bit_57_37 gnd C_bl
Cbb_57_37 bitb_57_37 gnd C_bl
Rb_57_38 bit_57_38 bit_57_39 R_bl
Rbb_57_38 bitb_57_38 bitb_57_39 R_bl
Cb_57_38 bit_57_38 gnd C_bl
Cbb_57_38 bitb_57_38 gnd C_bl
Rb_57_39 bit_57_39 bit_57_40 R_bl
Rbb_57_39 bitb_57_39 bitb_57_40 R_bl
Cb_57_39 bit_57_39 gnd C_bl
Cbb_57_39 bitb_57_39 gnd C_bl
Rb_57_40 bit_57_40 bit_57_41 R_bl
Rbb_57_40 bitb_57_40 bitb_57_41 R_bl
Cb_57_40 bit_57_40 gnd C_bl
Cbb_57_40 bitb_57_40 gnd C_bl
Rb_57_41 bit_57_41 bit_57_42 R_bl
Rbb_57_41 bitb_57_41 bitb_57_42 R_bl
Cb_57_41 bit_57_41 gnd C_bl
Cbb_57_41 bitb_57_41 gnd C_bl
Rb_57_42 bit_57_42 bit_57_43 R_bl
Rbb_57_42 bitb_57_42 bitb_57_43 R_bl
Cb_57_42 bit_57_42 gnd C_bl
Cbb_57_42 bitb_57_42 gnd C_bl
Rb_57_43 bit_57_43 bit_57_44 R_bl
Rbb_57_43 bitb_57_43 bitb_57_44 R_bl
Cb_57_43 bit_57_43 gnd C_bl
Cbb_57_43 bitb_57_43 gnd C_bl
Rb_57_44 bit_57_44 bit_57_45 R_bl
Rbb_57_44 bitb_57_44 bitb_57_45 R_bl
Cb_57_44 bit_57_44 gnd C_bl
Cbb_57_44 bitb_57_44 gnd C_bl
Rb_57_45 bit_57_45 bit_57_46 R_bl
Rbb_57_45 bitb_57_45 bitb_57_46 R_bl
Cb_57_45 bit_57_45 gnd C_bl
Cbb_57_45 bitb_57_45 gnd C_bl
Rb_57_46 bit_57_46 bit_57_47 R_bl
Rbb_57_46 bitb_57_46 bitb_57_47 R_bl
Cb_57_46 bit_57_46 gnd C_bl
Cbb_57_46 bitb_57_46 gnd C_bl
Rb_57_47 bit_57_47 bit_57_48 R_bl
Rbb_57_47 bitb_57_47 bitb_57_48 R_bl
Cb_57_47 bit_57_47 gnd C_bl
Cbb_57_47 bitb_57_47 gnd C_bl
Rb_57_48 bit_57_48 bit_57_49 R_bl
Rbb_57_48 bitb_57_48 bitb_57_49 R_bl
Cb_57_48 bit_57_48 gnd C_bl
Cbb_57_48 bitb_57_48 gnd C_bl
Rb_57_49 bit_57_49 bit_57_50 R_bl
Rbb_57_49 bitb_57_49 bitb_57_50 R_bl
Cb_57_49 bit_57_49 gnd C_bl
Cbb_57_49 bitb_57_49 gnd C_bl
Rb_57_50 bit_57_50 bit_57_51 R_bl
Rbb_57_50 bitb_57_50 bitb_57_51 R_bl
Cb_57_50 bit_57_50 gnd C_bl
Cbb_57_50 bitb_57_50 gnd C_bl
Rb_57_51 bit_57_51 bit_57_52 R_bl
Rbb_57_51 bitb_57_51 bitb_57_52 R_bl
Cb_57_51 bit_57_51 gnd C_bl
Cbb_57_51 bitb_57_51 gnd C_bl
Rb_57_52 bit_57_52 bit_57_53 R_bl
Rbb_57_52 bitb_57_52 bitb_57_53 R_bl
Cb_57_52 bit_57_52 gnd C_bl
Cbb_57_52 bitb_57_52 gnd C_bl
Rb_57_53 bit_57_53 bit_57_54 R_bl
Rbb_57_53 bitb_57_53 bitb_57_54 R_bl
Cb_57_53 bit_57_53 gnd C_bl
Cbb_57_53 bitb_57_53 gnd C_bl
Rb_57_54 bit_57_54 bit_57_55 R_bl
Rbb_57_54 bitb_57_54 bitb_57_55 R_bl
Cb_57_54 bit_57_54 gnd C_bl
Cbb_57_54 bitb_57_54 gnd C_bl
Rb_57_55 bit_57_55 bit_57_56 R_bl
Rbb_57_55 bitb_57_55 bitb_57_56 R_bl
Cb_57_55 bit_57_55 gnd C_bl
Cbb_57_55 bitb_57_55 gnd C_bl
Rb_57_56 bit_57_56 bit_57_57 R_bl
Rbb_57_56 bitb_57_56 bitb_57_57 R_bl
Cb_57_56 bit_57_56 gnd C_bl
Cbb_57_56 bitb_57_56 gnd C_bl
Rb_57_57 bit_57_57 bit_57_58 R_bl
Rbb_57_57 bitb_57_57 bitb_57_58 R_bl
Cb_57_57 bit_57_57 gnd C_bl
Cbb_57_57 bitb_57_57 gnd C_bl
Rb_57_58 bit_57_58 bit_57_59 R_bl
Rbb_57_58 bitb_57_58 bitb_57_59 R_bl
Cb_57_58 bit_57_58 gnd C_bl
Cbb_57_58 bitb_57_58 gnd C_bl
Rb_57_59 bit_57_59 bit_57_60 R_bl
Rbb_57_59 bitb_57_59 bitb_57_60 R_bl
Cb_57_59 bit_57_59 gnd C_bl
Cbb_57_59 bitb_57_59 gnd C_bl
Rb_57_60 bit_57_60 bit_57_61 R_bl
Rbb_57_60 bitb_57_60 bitb_57_61 R_bl
Cb_57_60 bit_57_60 gnd C_bl
Cbb_57_60 bitb_57_60 gnd C_bl
Rb_57_61 bit_57_61 bit_57_62 R_bl
Rbb_57_61 bitb_57_61 bitb_57_62 R_bl
Cb_57_61 bit_57_61 gnd C_bl
Cbb_57_61 bitb_57_61 gnd C_bl
Rb_57_62 bit_57_62 bit_57_63 R_bl
Rbb_57_62 bitb_57_62 bitb_57_63 R_bl
Cb_57_62 bit_57_62 gnd C_bl
Cbb_57_62 bitb_57_62 gnd C_bl
Rb_57_63 bit_57_63 bit_57_64 R_bl
Rbb_57_63 bitb_57_63 bitb_57_64 R_bl
Cb_57_63 bit_57_63 gnd C_bl
Cbb_57_63 bitb_57_63 gnd C_bl
Rb_57_64 bit_57_64 bit_57_65 R_bl
Rbb_57_64 bitb_57_64 bitb_57_65 R_bl
Cb_57_64 bit_57_64 gnd C_bl
Cbb_57_64 bitb_57_64 gnd C_bl
Rb_57_65 bit_57_65 bit_57_66 R_bl
Rbb_57_65 bitb_57_65 bitb_57_66 R_bl
Cb_57_65 bit_57_65 gnd C_bl
Cbb_57_65 bitb_57_65 gnd C_bl
Rb_57_66 bit_57_66 bit_57_67 R_bl
Rbb_57_66 bitb_57_66 bitb_57_67 R_bl
Cb_57_66 bit_57_66 gnd C_bl
Cbb_57_66 bitb_57_66 gnd C_bl
Rb_57_67 bit_57_67 bit_57_68 R_bl
Rbb_57_67 bitb_57_67 bitb_57_68 R_bl
Cb_57_67 bit_57_67 gnd C_bl
Cbb_57_67 bitb_57_67 gnd C_bl
Rb_57_68 bit_57_68 bit_57_69 R_bl
Rbb_57_68 bitb_57_68 bitb_57_69 R_bl
Cb_57_68 bit_57_68 gnd C_bl
Cbb_57_68 bitb_57_68 gnd C_bl
Rb_57_69 bit_57_69 bit_57_70 R_bl
Rbb_57_69 bitb_57_69 bitb_57_70 R_bl
Cb_57_69 bit_57_69 gnd C_bl
Cbb_57_69 bitb_57_69 gnd C_bl
Rb_57_70 bit_57_70 bit_57_71 R_bl
Rbb_57_70 bitb_57_70 bitb_57_71 R_bl
Cb_57_70 bit_57_70 gnd C_bl
Cbb_57_70 bitb_57_70 gnd C_bl
Rb_57_71 bit_57_71 bit_57_72 R_bl
Rbb_57_71 bitb_57_71 bitb_57_72 R_bl
Cb_57_71 bit_57_71 gnd C_bl
Cbb_57_71 bitb_57_71 gnd C_bl
Rb_57_72 bit_57_72 bit_57_73 R_bl
Rbb_57_72 bitb_57_72 bitb_57_73 R_bl
Cb_57_72 bit_57_72 gnd C_bl
Cbb_57_72 bitb_57_72 gnd C_bl
Rb_57_73 bit_57_73 bit_57_74 R_bl
Rbb_57_73 bitb_57_73 bitb_57_74 R_bl
Cb_57_73 bit_57_73 gnd C_bl
Cbb_57_73 bitb_57_73 gnd C_bl
Rb_57_74 bit_57_74 bit_57_75 R_bl
Rbb_57_74 bitb_57_74 bitb_57_75 R_bl
Cb_57_74 bit_57_74 gnd C_bl
Cbb_57_74 bitb_57_74 gnd C_bl
Rb_57_75 bit_57_75 bit_57_76 R_bl
Rbb_57_75 bitb_57_75 bitb_57_76 R_bl
Cb_57_75 bit_57_75 gnd C_bl
Cbb_57_75 bitb_57_75 gnd C_bl
Rb_57_76 bit_57_76 bit_57_77 R_bl
Rbb_57_76 bitb_57_76 bitb_57_77 R_bl
Cb_57_76 bit_57_76 gnd C_bl
Cbb_57_76 bitb_57_76 gnd C_bl
Rb_57_77 bit_57_77 bit_57_78 R_bl
Rbb_57_77 bitb_57_77 bitb_57_78 R_bl
Cb_57_77 bit_57_77 gnd C_bl
Cbb_57_77 bitb_57_77 gnd C_bl
Rb_57_78 bit_57_78 bit_57_79 R_bl
Rbb_57_78 bitb_57_78 bitb_57_79 R_bl
Cb_57_78 bit_57_78 gnd C_bl
Cbb_57_78 bitb_57_78 gnd C_bl
Rb_57_79 bit_57_79 bit_57_80 R_bl
Rbb_57_79 bitb_57_79 bitb_57_80 R_bl
Cb_57_79 bit_57_79 gnd C_bl
Cbb_57_79 bitb_57_79 gnd C_bl
Rb_57_80 bit_57_80 bit_57_81 R_bl
Rbb_57_80 bitb_57_80 bitb_57_81 R_bl
Cb_57_80 bit_57_80 gnd C_bl
Cbb_57_80 bitb_57_80 gnd C_bl
Rb_57_81 bit_57_81 bit_57_82 R_bl
Rbb_57_81 bitb_57_81 bitb_57_82 R_bl
Cb_57_81 bit_57_81 gnd C_bl
Cbb_57_81 bitb_57_81 gnd C_bl
Rb_57_82 bit_57_82 bit_57_83 R_bl
Rbb_57_82 bitb_57_82 bitb_57_83 R_bl
Cb_57_82 bit_57_82 gnd C_bl
Cbb_57_82 bitb_57_82 gnd C_bl
Rb_57_83 bit_57_83 bit_57_84 R_bl
Rbb_57_83 bitb_57_83 bitb_57_84 R_bl
Cb_57_83 bit_57_83 gnd C_bl
Cbb_57_83 bitb_57_83 gnd C_bl
Rb_57_84 bit_57_84 bit_57_85 R_bl
Rbb_57_84 bitb_57_84 bitb_57_85 R_bl
Cb_57_84 bit_57_84 gnd C_bl
Cbb_57_84 bitb_57_84 gnd C_bl
Rb_57_85 bit_57_85 bit_57_86 R_bl
Rbb_57_85 bitb_57_85 bitb_57_86 R_bl
Cb_57_85 bit_57_85 gnd C_bl
Cbb_57_85 bitb_57_85 gnd C_bl
Rb_57_86 bit_57_86 bit_57_87 R_bl
Rbb_57_86 bitb_57_86 bitb_57_87 R_bl
Cb_57_86 bit_57_86 gnd C_bl
Cbb_57_86 bitb_57_86 gnd C_bl
Rb_57_87 bit_57_87 bit_57_88 R_bl
Rbb_57_87 bitb_57_87 bitb_57_88 R_bl
Cb_57_87 bit_57_87 gnd C_bl
Cbb_57_87 bitb_57_87 gnd C_bl
Rb_57_88 bit_57_88 bit_57_89 R_bl
Rbb_57_88 bitb_57_88 bitb_57_89 R_bl
Cb_57_88 bit_57_88 gnd C_bl
Cbb_57_88 bitb_57_88 gnd C_bl
Rb_57_89 bit_57_89 bit_57_90 R_bl
Rbb_57_89 bitb_57_89 bitb_57_90 R_bl
Cb_57_89 bit_57_89 gnd C_bl
Cbb_57_89 bitb_57_89 gnd C_bl
Rb_57_90 bit_57_90 bit_57_91 R_bl
Rbb_57_90 bitb_57_90 bitb_57_91 R_bl
Cb_57_90 bit_57_90 gnd C_bl
Cbb_57_90 bitb_57_90 gnd C_bl
Rb_57_91 bit_57_91 bit_57_92 R_bl
Rbb_57_91 bitb_57_91 bitb_57_92 R_bl
Cb_57_91 bit_57_91 gnd C_bl
Cbb_57_91 bitb_57_91 gnd C_bl
Rb_57_92 bit_57_92 bit_57_93 R_bl
Rbb_57_92 bitb_57_92 bitb_57_93 R_bl
Cb_57_92 bit_57_92 gnd C_bl
Cbb_57_92 bitb_57_92 gnd C_bl
Rb_57_93 bit_57_93 bit_57_94 R_bl
Rbb_57_93 bitb_57_93 bitb_57_94 R_bl
Cb_57_93 bit_57_93 gnd C_bl
Cbb_57_93 bitb_57_93 gnd C_bl
Rb_57_94 bit_57_94 bit_57_95 R_bl
Rbb_57_94 bitb_57_94 bitb_57_95 R_bl
Cb_57_94 bit_57_94 gnd C_bl
Cbb_57_94 bitb_57_94 gnd C_bl
Rb_57_95 bit_57_95 bit_57_96 R_bl
Rbb_57_95 bitb_57_95 bitb_57_96 R_bl
Cb_57_95 bit_57_95 gnd C_bl
Cbb_57_95 bitb_57_95 gnd C_bl
Rb_57_96 bit_57_96 bit_57_97 R_bl
Rbb_57_96 bitb_57_96 bitb_57_97 R_bl
Cb_57_96 bit_57_96 gnd C_bl
Cbb_57_96 bitb_57_96 gnd C_bl
Rb_57_97 bit_57_97 bit_57_98 R_bl
Rbb_57_97 bitb_57_97 bitb_57_98 R_bl
Cb_57_97 bit_57_97 gnd C_bl
Cbb_57_97 bitb_57_97 gnd C_bl
Rb_57_98 bit_57_98 bit_57_99 R_bl
Rbb_57_98 bitb_57_98 bitb_57_99 R_bl
Cb_57_98 bit_57_98 gnd C_bl
Cbb_57_98 bitb_57_98 gnd C_bl
Rb_57_99 bit_57_99 bit_57_100 R_bl
Rbb_57_99 bitb_57_99 bitb_57_100 R_bl
Cb_57_99 bit_57_99 gnd C_bl
Cbb_57_99 bitb_57_99 gnd C_bl
Rb_58_0 bit_58_0 bit_58_1 R_bl
Rbb_58_0 bitb_58_0 bitb_58_1 R_bl
Cb_58_0 bit_58_0 gnd C_bl
Cbb_58_0 bitb_58_0 gnd C_bl
Rb_58_1 bit_58_1 bit_58_2 R_bl
Rbb_58_1 bitb_58_1 bitb_58_2 R_bl
Cb_58_1 bit_58_1 gnd C_bl
Cbb_58_1 bitb_58_1 gnd C_bl
Rb_58_2 bit_58_2 bit_58_3 R_bl
Rbb_58_2 bitb_58_2 bitb_58_3 R_bl
Cb_58_2 bit_58_2 gnd C_bl
Cbb_58_2 bitb_58_2 gnd C_bl
Rb_58_3 bit_58_3 bit_58_4 R_bl
Rbb_58_3 bitb_58_3 bitb_58_4 R_bl
Cb_58_3 bit_58_3 gnd C_bl
Cbb_58_3 bitb_58_3 gnd C_bl
Rb_58_4 bit_58_4 bit_58_5 R_bl
Rbb_58_4 bitb_58_4 bitb_58_5 R_bl
Cb_58_4 bit_58_4 gnd C_bl
Cbb_58_4 bitb_58_4 gnd C_bl
Rb_58_5 bit_58_5 bit_58_6 R_bl
Rbb_58_5 bitb_58_5 bitb_58_6 R_bl
Cb_58_5 bit_58_5 gnd C_bl
Cbb_58_5 bitb_58_5 gnd C_bl
Rb_58_6 bit_58_6 bit_58_7 R_bl
Rbb_58_6 bitb_58_6 bitb_58_7 R_bl
Cb_58_6 bit_58_6 gnd C_bl
Cbb_58_6 bitb_58_6 gnd C_bl
Rb_58_7 bit_58_7 bit_58_8 R_bl
Rbb_58_7 bitb_58_7 bitb_58_8 R_bl
Cb_58_7 bit_58_7 gnd C_bl
Cbb_58_7 bitb_58_7 gnd C_bl
Rb_58_8 bit_58_8 bit_58_9 R_bl
Rbb_58_8 bitb_58_8 bitb_58_9 R_bl
Cb_58_8 bit_58_8 gnd C_bl
Cbb_58_8 bitb_58_8 gnd C_bl
Rb_58_9 bit_58_9 bit_58_10 R_bl
Rbb_58_9 bitb_58_9 bitb_58_10 R_bl
Cb_58_9 bit_58_9 gnd C_bl
Cbb_58_9 bitb_58_9 gnd C_bl
Rb_58_10 bit_58_10 bit_58_11 R_bl
Rbb_58_10 bitb_58_10 bitb_58_11 R_bl
Cb_58_10 bit_58_10 gnd C_bl
Cbb_58_10 bitb_58_10 gnd C_bl
Rb_58_11 bit_58_11 bit_58_12 R_bl
Rbb_58_11 bitb_58_11 bitb_58_12 R_bl
Cb_58_11 bit_58_11 gnd C_bl
Cbb_58_11 bitb_58_11 gnd C_bl
Rb_58_12 bit_58_12 bit_58_13 R_bl
Rbb_58_12 bitb_58_12 bitb_58_13 R_bl
Cb_58_12 bit_58_12 gnd C_bl
Cbb_58_12 bitb_58_12 gnd C_bl
Rb_58_13 bit_58_13 bit_58_14 R_bl
Rbb_58_13 bitb_58_13 bitb_58_14 R_bl
Cb_58_13 bit_58_13 gnd C_bl
Cbb_58_13 bitb_58_13 gnd C_bl
Rb_58_14 bit_58_14 bit_58_15 R_bl
Rbb_58_14 bitb_58_14 bitb_58_15 R_bl
Cb_58_14 bit_58_14 gnd C_bl
Cbb_58_14 bitb_58_14 gnd C_bl
Rb_58_15 bit_58_15 bit_58_16 R_bl
Rbb_58_15 bitb_58_15 bitb_58_16 R_bl
Cb_58_15 bit_58_15 gnd C_bl
Cbb_58_15 bitb_58_15 gnd C_bl
Rb_58_16 bit_58_16 bit_58_17 R_bl
Rbb_58_16 bitb_58_16 bitb_58_17 R_bl
Cb_58_16 bit_58_16 gnd C_bl
Cbb_58_16 bitb_58_16 gnd C_bl
Rb_58_17 bit_58_17 bit_58_18 R_bl
Rbb_58_17 bitb_58_17 bitb_58_18 R_bl
Cb_58_17 bit_58_17 gnd C_bl
Cbb_58_17 bitb_58_17 gnd C_bl
Rb_58_18 bit_58_18 bit_58_19 R_bl
Rbb_58_18 bitb_58_18 bitb_58_19 R_bl
Cb_58_18 bit_58_18 gnd C_bl
Cbb_58_18 bitb_58_18 gnd C_bl
Rb_58_19 bit_58_19 bit_58_20 R_bl
Rbb_58_19 bitb_58_19 bitb_58_20 R_bl
Cb_58_19 bit_58_19 gnd C_bl
Cbb_58_19 bitb_58_19 gnd C_bl
Rb_58_20 bit_58_20 bit_58_21 R_bl
Rbb_58_20 bitb_58_20 bitb_58_21 R_bl
Cb_58_20 bit_58_20 gnd C_bl
Cbb_58_20 bitb_58_20 gnd C_bl
Rb_58_21 bit_58_21 bit_58_22 R_bl
Rbb_58_21 bitb_58_21 bitb_58_22 R_bl
Cb_58_21 bit_58_21 gnd C_bl
Cbb_58_21 bitb_58_21 gnd C_bl
Rb_58_22 bit_58_22 bit_58_23 R_bl
Rbb_58_22 bitb_58_22 bitb_58_23 R_bl
Cb_58_22 bit_58_22 gnd C_bl
Cbb_58_22 bitb_58_22 gnd C_bl
Rb_58_23 bit_58_23 bit_58_24 R_bl
Rbb_58_23 bitb_58_23 bitb_58_24 R_bl
Cb_58_23 bit_58_23 gnd C_bl
Cbb_58_23 bitb_58_23 gnd C_bl
Rb_58_24 bit_58_24 bit_58_25 R_bl
Rbb_58_24 bitb_58_24 bitb_58_25 R_bl
Cb_58_24 bit_58_24 gnd C_bl
Cbb_58_24 bitb_58_24 gnd C_bl
Rb_58_25 bit_58_25 bit_58_26 R_bl
Rbb_58_25 bitb_58_25 bitb_58_26 R_bl
Cb_58_25 bit_58_25 gnd C_bl
Cbb_58_25 bitb_58_25 gnd C_bl
Rb_58_26 bit_58_26 bit_58_27 R_bl
Rbb_58_26 bitb_58_26 bitb_58_27 R_bl
Cb_58_26 bit_58_26 gnd C_bl
Cbb_58_26 bitb_58_26 gnd C_bl
Rb_58_27 bit_58_27 bit_58_28 R_bl
Rbb_58_27 bitb_58_27 bitb_58_28 R_bl
Cb_58_27 bit_58_27 gnd C_bl
Cbb_58_27 bitb_58_27 gnd C_bl
Rb_58_28 bit_58_28 bit_58_29 R_bl
Rbb_58_28 bitb_58_28 bitb_58_29 R_bl
Cb_58_28 bit_58_28 gnd C_bl
Cbb_58_28 bitb_58_28 gnd C_bl
Rb_58_29 bit_58_29 bit_58_30 R_bl
Rbb_58_29 bitb_58_29 bitb_58_30 R_bl
Cb_58_29 bit_58_29 gnd C_bl
Cbb_58_29 bitb_58_29 gnd C_bl
Rb_58_30 bit_58_30 bit_58_31 R_bl
Rbb_58_30 bitb_58_30 bitb_58_31 R_bl
Cb_58_30 bit_58_30 gnd C_bl
Cbb_58_30 bitb_58_30 gnd C_bl
Rb_58_31 bit_58_31 bit_58_32 R_bl
Rbb_58_31 bitb_58_31 bitb_58_32 R_bl
Cb_58_31 bit_58_31 gnd C_bl
Cbb_58_31 bitb_58_31 gnd C_bl
Rb_58_32 bit_58_32 bit_58_33 R_bl
Rbb_58_32 bitb_58_32 bitb_58_33 R_bl
Cb_58_32 bit_58_32 gnd C_bl
Cbb_58_32 bitb_58_32 gnd C_bl
Rb_58_33 bit_58_33 bit_58_34 R_bl
Rbb_58_33 bitb_58_33 bitb_58_34 R_bl
Cb_58_33 bit_58_33 gnd C_bl
Cbb_58_33 bitb_58_33 gnd C_bl
Rb_58_34 bit_58_34 bit_58_35 R_bl
Rbb_58_34 bitb_58_34 bitb_58_35 R_bl
Cb_58_34 bit_58_34 gnd C_bl
Cbb_58_34 bitb_58_34 gnd C_bl
Rb_58_35 bit_58_35 bit_58_36 R_bl
Rbb_58_35 bitb_58_35 bitb_58_36 R_bl
Cb_58_35 bit_58_35 gnd C_bl
Cbb_58_35 bitb_58_35 gnd C_bl
Rb_58_36 bit_58_36 bit_58_37 R_bl
Rbb_58_36 bitb_58_36 bitb_58_37 R_bl
Cb_58_36 bit_58_36 gnd C_bl
Cbb_58_36 bitb_58_36 gnd C_bl
Rb_58_37 bit_58_37 bit_58_38 R_bl
Rbb_58_37 bitb_58_37 bitb_58_38 R_bl
Cb_58_37 bit_58_37 gnd C_bl
Cbb_58_37 bitb_58_37 gnd C_bl
Rb_58_38 bit_58_38 bit_58_39 R_bl
Rbb_58_38 bitb_58_38 bitb_58_39 R_bl
Cb_58_38 bit_58_38 gnd C_bl
Cbb_58_38 bitb_58_38 gnd C_bl
Rb_58_39 bit_58_39 bit_58_40 R_bl
Rbb_58_39 bitb_58_39 bitb_58_40 R_bl
Cb_58_39 bit_58_39 gnd C_bl
Cbb_58_39 bitb_58_39 gnd C_bl
Rb_58_40 bit_58_40 bit_58_41 R_bl
Rbb_58_40 bitb_58_40 bitb_58_41 R_bl
Cb_58_40 bit_58_40 gnd C_bl
Cbb_58_40 bitb_58_40 gnd C_bl
Rb_58_41 bit_58_41 bit_58_42 R_bl
Rbb_58_41 bitb_58_41 bitb_58_42 R_bl
Cb_58_41 bit_58_41 gnd C_bl
Cbb_58_41 bitb_58_41 gnd C_bl
Rb_58_42 bit_58_42 bit_58_43 R_bl
Rbb_58_42 bitb_58_42 bitb_58_43 R_bl
Cb_58_42 bit_58_42 gnd C_bl
Cbb_58_42 bitb_58_42 gnd C_bl
Rb_58_43 bit_58_43 bit_58_44 R_bl
Rbb_58_43 bitb_58_43 bitb_58_44 R_bl
Cb_58_43 bit_58_43 gnd C_bl
Cbb_58_43 bitb_58_43 gnd C_bl
Rb_58_44 bit_58_44 bit_58_45 R_bl
Rbb_58_44 bitb_58_44 bitb_58_45 R_bl
Cb_58_44 bit_58_44 gnd C_bl
Cbb_58_44 bitb_58_44 gnd C_bl
Rb_58_45 bit_58_45 bit_58_46 R_bl
Rbb_58_45 bitb_58_45 bitb_58_46 R_bl
Cb_58_45 bit_58_45 gnd C_bl
Cbb_58_45 bitb_58_45 gnd C_bl
Rb_58_46 bit_58_46 bit_58_47 R_bl
Rbb_58_46 bitb_58_46 bitb_58_47 R_bl
Cb_58_46 bit_58_46 gnd C_bl
Cbb_58_46 bitb_58_46 gnd C_bl
Rb_58_47 bit_58_47 bit_58_48 R_bl
Rbb_58_47 bitb_58_47 bitb_58_48 R_bl
Cb_58_47 bit_58_47 gnd C_bl
Cbb_58_47 bitb_58_47 gnd C_bl
Rb_58_48 bit_58_48 bit_58_49 R_bl
Rbb_58_48 bitb_58_48 bitb_58_49 R_bl
Cb_58_48 bit_58_48 gnd C_bl
Cbb_58_48 bitb_58_48 gnd C_bl
Rb_58_49 bit_58_49 bit_58_50 R_bl
Rbb_58_49 bitb_58_49 bitb_58_50 R_bl
Cb_58_49 bit_58_49 gnd C_bl
Cbb_58_49 bitb_58_49 gnd C_bl
Rb_58_50 bit_58_50 bit_58_51 R_bl
Rbb_58_50 bitb_58_50 bitb_58_51 R_bl
Cb_58_50 bit_58_50 gnd C_bl
Cbb_58_50 bitb_58_50 gnd C_bl
Rb_58_51 bit_58_51 bit_58_52 R_bl
Rbb_58_51 bitb_58_51 bitb_58_52 R_bl
Cb_58_51 bit_58_51 gnd C_bl
Cbb_58_51 bitb_58_51 gnd C_bl
Rb_58_52 bit_58_52 bit_58_53 R_bl
Rbb_58_52 bitb_58_52 bitb_58_53 R_bl
Cb_58_52 bit_58_52 gnd C_bl
Cbb_58_52 bitb_58_52 gnd C_bl
Rb_58_53 bit_58_53 bit_58_54 R_bl
Rbb_58_53 bitb_58_53 bitb_58_54 R_bl
Cb_58_53 bit_58_53 gnd C_bl
Cbb_58_53 bitb_58_53 gnd C_bl
Rb_58_54 bit_58_54 bit_58_55 R_bl
Rbb_58_54 bitb_58_54 bitb_58_55 R_bl
Cb_58_54 bit_58_54 gnd C_bl
Cbb_58_54 bitb_58_54 gnd C_bl
Rb_58_55 bit_58_55 bit_58_56 R_bl
Rbb_58_55 bitb_58_55 bitb_58_56 R_bl
Cb_58_55 bit_58_55 gnd C_bl
Cbb_58_55 bitb_58_55 gnd C_bl
Rb_58_56 bit_58_56 bit_58_57 R_bl
Rbb_58_56 bitb_58_56 bitb_58_57 R_bl
Cb_58_56 bit_58_56 gnd C_bl
Cbb_58_56 bitb_58_56 gnd C_bl
Rb_58_57 bit_58_57 bit_58_58 R_bl
Rbb_58_57 bitb_58_57 bitb_58_58 R_bl
Cb_58_57 bit_58_57 gnd C_bl
Cbb_58_57 bitb_58_57 gnd C_bl
Rb_58_58 bit_58_58 bit_58_59 R_bl
Rbb_58_58 bitb_58_58 bitb_58_59 R_bl
Cb_58_58 bit_58_58 gnd C_bl
Cbb_58_58 bitb_58_58 gnd C_bl
Rb_58_59 bit_58_59 bit_58_60 R_bl
Rbb_58_59 bitb_58_59 bitb_58_60 R_bl
Cb_58_59 bit_58_59 gnd C_bl
Cbb_58_59 bitb_58_59 gnd C_bl
Rb_58_60 bit_58_60 bit_58_61 R_bl
Rbb_58_60 bitb_58_60 bitb_58_61 R_bl
Cb_58_60 bit_58_60 gnd C_bl
Cbb_58_60 bitb_58_60 gnd C_bl
Rb_58_61 bit_58_61 bit_58_62 R_bl
Rbb_58_61 bitb_58_61 bitb_58_62 R_bl
Cb_58_61 bit_58_61 gnd C_bl
Cbb_58_61 bitb_58_61 gnd C_bl
Rb_58_62 bit_58_62 bit_58_63 R_bl
Rbb_58_62 bitb_58_62 bitb_58_63 R_bl
Cb_58_62 bit_58_62 gnd C_bl
Cbb_58_62 bitb_58_62 gnd C_bl
Rb_58_63 bit_58_63 bit_58_64 R_bl
Rbb_58_63 bitb_58_63 bitb_58_64 R_bl
Cb_58_63 bit_58_63 gnd C_bl
Cbb_58_63 bitb_58_63 gnd C_bl
Rb_58_64 bit_58_64 bit_58_65 R_bl
Rbb_58_64 bitb_58_64 bitb_58_65 R_bl
Cb_58_64 bit_58_64 gnd C_bl
Cbb_58_64 bitb_58_64 gnd C_bl
Rb_58_65 bit_58_65 bit_58_66 R_bl
Rbb_58_65 bitb_58_65 bitb_58_66 R_bl
Cb_58_65 bit_58_65 gnd C_bl
Cbb_58_65 bitb_58_65 gnd C_bl
Rb_58_66 bit_58_66 bit_58_67 R_bl
Rbb_58_66 bitb_58_66 bitb_58_67 R_bl
Cb_58_66 bit_58_66 gnd C_bl
Cbb_58_66 bitb_58_66 gnd C_bl
Rb_58_67 bit_58_67 bit_58_68 R_bl
Rbb_58_67 bitb_58_67 bitb_58_68 R_bl
Cb_58_67 bit_58_67 gnd C_bl
Cbb_58_67 bitb_58_67 gnd C_bl
Rb_58_68 bit_58_68 bit_58_69 R_bl
Rbb_58_68 bitb_58_68 bitb_58_69 R_bl
Cb_58_68 bit_58_68 gnd C_bl
Cbb_58_68 bitb_58_68 gnd C_bl
Rb_58_69 bit_58_69 bit_58_70 R_bl
Rbb_58_69 bitb_58_69 bitb_58_70 R_bl
Cb_58_69 bit_58_69 gnd C_bl
Cbb_58_69 bitb_58_69 gnd C_bl
Rb_58_70 bit_58_70 bit_58_71 R_bl
Rbb_58_70 bitb_58_70 bitb_58_71 R_bl
Cb_58_70 bit_58_70 gnd C_bl
Cbb_58_70 bitb_58_70 gnd C_bl
Rb_58_71 bit_58_71 bit_58_72 R_bl
Rbb_58_71 bitb_58_71 bitb_58_72 R_bl
Cb_58_71 bit_58_71 gnd C_bl
Cbb_58_71 bitb_58_71 gnd C_bl
Rb_58_72 bit_58_72 bit_58_73 R_bl
Rbb_58_72 bitb_58_72 bitb_58_73 R_bl
Cb_58_72 bit_58_72 gnd C_bl
Cbb_58_72 bitb_58_72 gnd C_bl
Rb_58_73 bit_58_73 bit_58_74 R_bl
Rbb_58_73 bitb_58_73 bitb_58_74 R_bl
Cb_58_73 bit_58_73 gnd C_bl
Cbb_58_73 bitb_58_73 gnd C_bl
Rb_58_74 bit_58_74 bit_58_75 R_bl
Rbb_58_74 bitb_58_74 bitb_58_75 R_bl
Cb_58_74 bit_58_74 gnd C_bl
Cbb_58_74 bitb_58_74 gnd C_bl
Rb_58_75 bit_58_75 bit_58_76 R_bl
Rbb_58_75 bitb_58_75 bitb_58_76 R_bl
Cb_58_75 bit_58_75 gnd C_bl
Cbb_58_75 bitb_58_75 gnd C_bl
Rb_58_76 bit_58_76 bit_58_77 R_bl
Rbb_58_76 bitb_58_76 bitb_58_77 R_bl
Cb_58_76 bit_58_76 gnd C_bl
Cbb_58_76 bitb_58_76 gnd C_bl
Rb_58_77 bit_58_77 bit_58_78 R_bl
Rbb_58_77 bitb_58_77 bitb_58_78 R_bl
Cb_58_77 bit_58_77 gnd C_bl
Cbb_58_77 bitb_58_77 gnd C_bl
Rb_58_78 bit_58_78 bit_58_79 R_bl
Rbb_58_78 bitb_58_78 bitb_58_79 R_bl
Cb_58_78 bit_58_78 gnd C_bl
Cbb_58_78 bitb_58_78 gnd C_bl
Rb_58_79 bit_58_79 bit_58_80 R_bl
Rbb_58_79 bitb_58_79 bitb_58_80 R_bl
Cb_58_79 bit_58_79 gnd C_bl
Cbb_58_79 bitb_58_79 gnd C_bl
Rb_58_80 bit_58_80 bit_58_81 R_bl
Rbb_58_80 bitb_58_80 bitb_58_81 R_bl
Cb_58_80 bit_58_80 gnd C_bl
Cbb_58_80 bitb_58_80 gnd C_bl
Rb_58_81 bit_58_81 bit_58_82 R_bl
Rbb_58_81 bitb_58_81 bitb_58_82 R_bl
Cb_58_81 bit_58_81 gnd C_bl
Cbb_58_81 bitb_58_81 gnd C_bl
Rb_58_82 bit_58_82 bit_58_83 R_bl
Rbb_58_82 bitb_58_82 bitb_58_83 R_bl
Cb_58_82 bit_58_82 gnd C_bl
Cbb_58_82 bitb_58_82 gnd C_bl
Rb_58_83 bit_58_83 bit_58_84 R_bl
Rbb_58_83 bitb_58_83 bitb_58_84 R_bl
Cb_58_83 bit_58_83 gnd C_bl
Cbb_58_83 bitb_58_83 gnd C_bl
Rb_58_84 bit_58_84 bit_58_85 R_bl
Rbb_58_84 bitb_58_84 bitb_58_85 R_bl
Cb_58_84 bit_58_84 gnd C_bl
Cbb_58_84 bitb_58_84 gnd C_bl
Rb_58_85 bit_58_85 bit_58_86 R_bl
Rbb_58_85 bitb_58_85 bitb_58_86 R_bl
Cb_58_85 bit_58_85 gnd C_bl
Cbb_58_85 bitb_58_85 gnd C_bl
Rb_58_86 bit_58_86 bit_58_87 R_bl
Rbb_58_86 bitb_58_86 bitb_58_87 R_bl
Cb_58_86 bit_58_86 gnd C_bl
Cbb_58_86 bitb_58_86 gnd C_bl
Rb_58_87 bit_58_87 bit_58_88 R_bl
Rbb_58_87 bitb_58_87 bitb_58_88 R_bl
Cb_58_87 bit_58_87 gnd C_bl
Cbb_58_87 bitb_58_87 gnd C_bl
Rb_58_88 bit_58_88 bit_58_89 R_bl
Rbb_58_88 bitb_58_88 bitb_58_89 R_bl
Cb_58_88 bit_58_88 gnd C_bl
Cbb_58_88 bitb_58_88 gnd C_bl
Rb_58_89 bit_58_89 bit_58_90 R_bl
Rbb_58_89 bitb_58_89 bitb_58_90 R_bl
Cb_58_89 bit_58_89 gnd C_bl
Cbb_58_89 bitb_58_89 gnd C_bl
Rb_58_90 bit_58_90 bit_58_91 R_bl
Rbb_58_90 bitb_58_90 bitb_58_91 R_bl
Cb_58_90 bit_58_90 gnd C_bl
Cbb_58_90 bitb_58_90 gnd C_bl
Rb_58_91 bit_58_91 bit_58_92 R_bl
Rbb_58_91 bitb_58_91 bitb_58_92 R_bl
Cb_58_91 bit_58_91 gnd C_bl
Cbb_58_91 bitb_58_91 gnd C_bl
Rb_58_92 bit_58_92 bit_58_93 R_bl
Rbb_58_92 bitb_58_92 bitb_58_93 R_bl
Cb_58_92 bit_58_92 gnd C_bl
Cbb_58_92 bitb_58_92 gnd C_bl
Rb_58_93 bit_58_93 bit_58_94 R_bl
Rbb_58_93 bitb_58_93 bitb_58_94 R_bl
Cb_58_93 bit_58_93 gnd C_bl
Cbb_58_93 bitb_58_93 gnd C_bl
Rb_58_94 bit_58_94 bit_58_95 R_bl
Rbb_58_94 bitb_58_94 bitb_58_95 R_bl
Cb_58_94 bit_58_94 gnd C_bl
Cbb_58_94 bitb_58_94 gnd C_bl
Rb_58_95 bit_58_95 bit_58_96 R_bl
Rbb_58_95 bitb_58_95 bitb_58_96 R_bl
Cb_58_95 bit_58_95 gnd C_bl
Cbb_58_95 bitb_58_95 gnd C_bl
Rb_58_96 bit_58_96 bit_58_97 R_bl
Rbb_58_96 bitb_58_96 bitb_58_97 R_bl
Cb_58_96 bit_58_96 gnd C_bl
Cbb_58_96 bitb_58_96 gnd C_bl
Rb_58_97 bit_58_97 bit_58_98 R_bl
Rbb_58_97 bitb_58_97 bitb_58_98 R_bl
Cb_58_97 bit_58_97 gnd C_bl
Cbb_58_97 bitb_58_97 gnd C_bl
Rb_58_98 bit_58_98 bit_58_99 R_bl
Rbb_58_98 bitb_58_98 bitb_58_99 R_bl
Cb_58_98 bit_58_98 gnd C_bl
Cbb_58_98 bitb_58_98 gnd C_bl
Rb_58_99 bit_58_99 bit_58_100 R_bl
Rbb_58_99 bitb_58_99 bitb_58_100 R_bl
Cb_58_99 bit_58_99 gnd C_bl
Cbb_58_99 bitb_58_99 gnd C_bl
Rb_59_0 bit_59_0 bit_59_1 R_bl
Rbb_59_0 bitb_59_0 bitb_59_1 R_bl
Cb_59_0 bit_59_0 gnd C_bl
Cbb_59_0 bitb_59_0 gnd C_bl
Rb_59_1 bit_59_1 bit_59_2 R_bl
Rbb_59_1 bitb_59_1 bitb_59_2 R_bl
Cb_59_1 bit_59_1 gnd C_bl
Cbb_59_1 bitb_59_1 gnd C_bl
Rb_59_2 bit_59_2 bit_59_3 R_bl
Rbb_59_2 bitb_59_2 bitb_59_3 R_bl
Cb_59_2 bit_59_2 gnd C_bl
Cbb_59_2 bitb_59_2 gnd C_bl
Rb_59_3 bit_59_3 bit_59_4 R_bl
Rbb_59_3 bitb_59_3 bitb_59_4 R_bl
Cb_59_3 bit_59_3 gnd C_bl
Cbb_59_3 bitb_59_3 gnd C_bl
Rb_59_4 bit_59_4 bit_59_5 R_bl
Rbb_59_4 bitb_59_4 bitb_59_5 R_bl
Cb_59_4 bit_59_4 gnd C_bl
Cbb_59_4 bitb_59_4 gnd C_bl
Rb_59_5 bit_59_5 bit_59_6 R_bl
Rbb_59_5 bitb_59_5 bitb_59_6 R_bl
Cb_59_5 bit_59_5 gnd C_bl
Cbb_59_5 bitb_59_5 gnd C_bl
Rb_59_6 bit_59_6 bit_59_7 R_bl
Rbb_59_6 bitb_59_6 bitb_59_7 R_bl
Cb_59_6 bit_59_6 gnd C_bl
Cbb_59_6 bitb_59_6 gnd C_bl
Rb_59_7 bit_59_7 bit_59_8 R_bl
Rbb_59_7 bitb_59_7 bitb_59_8 R_bl
Cb_59_7 bit_59_7 gnd C_bl
Cbb_59_7 bitb_59_7 gnd C_bl
Rb_59_8 bit_59_8 bit_59_9 R_bl
Rbb_59_8 bitb_59_8 bitb_59_9 R_bl
Cb_59_8 bit_59_8 gnd C_bl
Cbb_59_8 bitb_59_8 gnd C_bl
Rb_59_9 bit_59_9 bit_59_10 R_bl
Rbb_59_9 bitb_59_9 bitb_59_10 R_bl
Cb_59_9 bit_59_9 gnd C_bl
Cbb_59_9 bitb_59_9 gnd C_bl
Rb_59_10 bit_59_10 bit_59_11 R_bl
Rbb_59_10 bitb_59_10 bitb_59_11 R_bl
Cb_59_10 bit_59_10 gnd C_bl
Cbb_59_10 bitb_59_10 gnd C_bl
Rb_59_11 bit_59_11 bit_59_12 R_bl
Rbb_59_11 bitb_59_11 bitb_59_12 R_bl
Cb_59_11 bit_59_11 gnd C_bl
Cbb_59_11 bitb_59_11 gnd C_bl
Rb_59_12 bit_59_12 bit_59_13 R_bl
Rbb_59_12 bitb_59_12 bitb_59_13 R_bl
Cb_59_12 bit_59_12 gnd C_bl
Cbb_59_12 bitb_59_12 gnd C_bl
Rb_59_13 bit_59_13 bit_59_14 R_bl
Rbb_59_13 bitb_59_13 bitb_59_14 R_bl
Cb_59_13 bit_59_13 gnd C_bl
Cbb_59_13 bitb_59_13 gnd C_bl
Rb_59_14 bit_59_14 bit_59_15 R_bl
Rbb_59_14 bitb_59_14 bitb_59_15 R_bl
Cb_59_14 bit_59_14 gnd C_bl
Cbb_59_14 bitb_59_14 gnd C_bl
Rb_59_15 bit_59_15 bit_59_16 R_bl
Rbb_59_15 bitb_59_15 bitb_59_16 R_bl
Cb_59_15 bit_59_15 gnd C_bl
Cbb_59_15 bitb_59_15 gnd C_bl
Rb_59_16 bit_59_16 bit_59_17 R_bl
Rbb_59_16 bitb_59_16 bitb_59_17 R_bl
Cb_59_16 bit_59_16 gnd C_bl
Cbb_59_16 bitb_59_16 gnd C_bl
Rb_59_17 bit_59_17 bit_59_18 R_bl
Rbb_59_17 bitb_59_17 bitb_59_18 R_bl
Cb_59_17 bit_59_17 gnd C_bl
Cbb_59_17 bitb_59_17 gnd C_bl
Rb_59_18 bit_59_18 bit_59_19 R_bl
Rbb_59_18 bitb_59_18 bitb_59_19 R_bl
Cb_59_18 bit_59_18 gnd C_bl
Cbb_59_18 bitb_59_18 gnd C_bl
Rb_59_19 bit_59_19 bit_59_20 R_bl
Rbb_59_19 bitb_59_19 bitb_59_20 R_bl
Cb_59_19 bit_59_19 gnd C_bl
Cbb_59_19 bitb_59_19 gnd C_bl
Rb_59_20 bit_59_20 bit_59_21 R_bl
Rbb_59_20 bitb_59_20 bitb_59_21 R_bl
Cb_59_20 bit_59_20 gnd C_bl
Cbb_59_20 bitb_59_20 gnd C_bl
Rb_59_21 bit_59_21 bit_59_22 R_bl
Rbb_59_21 bitb_59_21 bitb_59_22 R_bl
Cb_59_21 bit_59_21 gnd C_bl
Cbb_59_21 bitb_59_21 gnd C_bl
Rb_59_22 bit_59_22 bit_59_23 R_bl
Rbb_59_22 bitb_59_22 bitb_59_23 R_bl
Cb_59_22 bit_59_22 gnd C_bl
Cbb_59_22 bitb_59_22 gnd C_bl
Rb_59_23 bit_59_23 bit_59_24 R_bl
Rbb_59_23 bitb_59_23 bitb_59_24 R_bl
Cb_59_23 bit_59_23 gnd C_bl
Cbb_59_23 bitb_59_23 gnd C_bl
Rb_59_24 bit_59_24 bit_59_25 R_bl
Rbb_59_24 bitb_59_24 bitb_59_25 R_bl
Cb_59_24 bit_59_24 gnd C_bl
Cbb_59_24 bitb_59_24 gnd C_bl
Rb_59_25 bit_59_25 bit_59_26 R_bl
Rbb_59_25 bitb_59_25 bitb_59_26 R_bl
Cb_59_25 bit_59_25 gnd C_bl
Cbb_59_25 bitb_59_25 gnd C_bl
Rb_59_26 bit_59_26 bit_59_27 R_bl
Rbb_59_26 bitb_59_26 bitb_59_27 R_bl
Cb_59_26 bit_59_26 gnd C_bl
Cbb_59_26 bitb_59_26 gnd C_bl
Rb_59_27 bit_59_27 bit_59_28 R_bl
Rbb_59_27 bitb_59_27 bitb_59_28 R_bl
Cb_59_27 bit_59_27 gnd C_bl
Cbb_59_27 bitb_59_27 gnd C_bl
Rb_59_28 bit_59_28 bit_59_29 R_bl
Rbb_59_28 bitb_59_28 bitb_59_29 R_bl
Cb_59_28 bit_59_28 gnd C_bl
Cbb_59_28 bitb_59_28 gnd C_bl
Rb_59_29 bit_59_29 bit_59_30 R_bl
Rbb_59_29 bitb_59_29 bitb_59_30 R_bl
Cb_59_29 bit_59_29 gnd C_bl
Cbb_59_29 bitb_59_29 gnd C_bl
Rb_59_30 bit_59_30 bit_59_31 R_bl
Rbb_59_30 bitb_59_30 bitb_59_31 R_bl
Cb_59_30 bit_59_30 gnd C_bl
Cbb_59_30 bitb_59_30 gnd C_bl
Rb_59_31 bit_59_31 bit_59_32 R_bl
Rbb_59_31 bitb_59_31 bitb_59_32 R_bl
Cb_59_31 bit_59_31 gnd C_bl
Cbb_59_31 bitb_59_31 gnd C_bl
Rb_59_32 bit_59_32 bit_59_33 R_bl
Rbb_59_32 bitb_59_32 bitb_59_33 R_bl
Cb_59_32 bit_59_32 gnd C_bl
Cbb_59_32 bitb_59_32 gnd C_bl
Rb_59_33 bit_59_33 bit_59_34 R_bl
Rbb_59_33 bitb_59_33 bitb_59_34 R_bl
Cb_59_33 bit_59_33 gnd C_bl
Cbb_59_33 bitb_59_33 gnd C_bl
Rb_59_34 bit_59_34 bit_59_35 R_bl
Rbb_59_34 bitb_59_34 bitb_59_35 R_bl
Cb_59_34 bit_59_34 gnd C_bl
Cbb_59_34 bitb_59_34 gnd C_bl
Rb_59_35 bit_59_35 bit_59_36 R_bl
Rbb_59_35 bitb_59_35 bitb_59_36 R_bl
Cb_59_35 bit_59_35 gnd C_bl
Cbb_59_35 bitb_59_35 gnd C_bl
Rb_59_36 bit_59_36 bit_59_37 R_bl
Rbb_59_36 bitb_59_36 bitb_59_37 R_bl
Cb_59_36 bit_59_36 gnd C_bl
Cbb_59_36 bitb_59_36 gnd C_bl
Rb_59_37 bit_59_37 bit_59_38 R_bl
Rbb_59_37 bitb_59_37 bitb_59_38 R_bl
Cb_59_37 bit_59_37 gnd C_bl
Cbb_59_37 bitb_59_37 gnd C_bl
Rb_59_38 bit_59_38 bit_59_39 R_bl
Rbb_59_38 bitb_59_38 bitb_59_39 R_bl
Cb_59_38 bit_59_38 gnd C_bl
Cbb_59_38 bitb_59_38 gnd C_bl
Rb_59_39 bit_59_39 bit_59_40 R_bl
Rbb_59_39 bitb_59_39 bitb_59_40 R_bl
Cb_59_39 bit_59_39 gnd C_bl
Cbb_59_39 bitb_59_39 gnd C_bl
Rb_59_40 bit_59_40 bit_59_41 R_bl
Rbb_59_40 bitb_59_40 bitb_59_41 R_bl
Cb_59_40 bit_59_40 gnd C_bl
Cbb_59_40 bitb_59_40 gnd C_bl
Rb_59_41 bit_59_41 bit_59_42 R_bl
Rbb_59_41 bitb_59_41 bitb_59_42 R_bl
Cb_59_41 bit_59_41 gnd C_bl
Cbb_59_41 bitb_59_41 gnd C_bl
Rb_59_42 bit_59_42 bit_59_43 R_bl
Rbb_59_42 bitb_59_42 bitb_59_43 R_bl
Cb_59_42 bit_59_42 gnd C_bl
Cbb_59_42 bitb_59_42 gnd C_bl
Rb_59_43 bit_59_43 bit_59_44 R_bl
Rbb_59_43 bitb_59_43 bitb_59_44 R_bl
Cb_59_43 bit_59_43 gnd C_bl
Cbb_59_43 bitb_59_43 gnd C_bl
Rb_59_44 bit_59_44 bit_59_45 R_bl
Rbb_59_44 bitb_59_44 bitb_59_45 R_bl
Cb_59_44 bit_59_44 gnd C_bl
Cbb_59_44 bitb_59_44 gnd C_bl
Rb_59_45 bit_59_45 bit_59_46 R_bl
Rbb_59_45 bitb_59_45 bitb_59_46 R_bl
Cb_59_45 bit_59_45 gnd C_bl
Cbb_59_45 bitb_59_45 gnd C_bl
Rb_59_46 bit_59_46 bit_59_47 R_bl
Rbb_59_46 bitb_59_46 bitb_59_47 R_bl
Cb_59_46 bit_59_46 gnd C_bl
Cbb_59_46 bitb_59_46 gnd C_bl
Rb_59_47 bit_59_47 bit_59_48 R_bl
Rbb_59_47 bitb_59_47 bitb_59_48 R_bl
Cb_59_47 bit_59_47 gnd C_bl
Cbb_59_47 bitb_59_47 gnd C_bl
Rb_59_48 bit_59_48 bit_59_49 R_bl
Rbb_59_48 bitb_59_48 bitb_59_49 R_bl
Cb_59_48 bit_59_48 gnd C_bl
Cbb_59_48 bitb_59_48 gnd C_bl
Rb_59_49 bit_59_49 bit_59_50 R_bl
Rbb_59_49 bitb_59_49 bitb_59_50 R_bl
Cb_59_49 bit_59_49 gnd C_bl
Cbb_59_49 bitb_59_49 gnd C_bl
Rb_59_50 bit_59_50 bit_59_51 R_bl
Rbb_59_50 bitb_59_50 bitb_59_51 R_bl
Cb_59_50 bit_59_50 gnd C_bl
Cbb_59_50 bitb_59_50 gnd C_bl
Rb_59_51 bit_59_51 bit_59_52 R_bl
Rbb_59_51 bitb_59_51 bitb_59_52 R_bl
Cb_59_51 bit_59_51 gnd C_bl
Cbb_59_51 bitb_59_51 gnd C_bl
Rb_59_52 bit_59_52 bit_59_53 R_bl
Rbb_59_52 bitb_59_52 bitb_59_53 R_bl
Cb_59_52 bit_59_52 gnd C_bl
Cbb_59_52 bitb_59_52 gnd C_bl
Rb_59_53 bit_59_53 bit_59_54 R_bl
Rbb_59_53 bitb_59_53 bitb_59_54 R_bl
Cb_59_53 bit_59_53 gnd C_bl
Cbb_59_53 bitb_59_53 gnd C_bl
Rb_59_54 bit_59_54 bit_59_55 R_bl
Rbb_59_54 bitb_59_54 bitb_59_55 R_bl
Cb_59_54 bit_59_54 gnd C_bl
Cbb_59_54 bitb_59_54 gnd C_bl
Rb_59_55 bit_59_55 bit_59_56 R_bl
Rbb_59_55 bitb_59_55 bitb_59_56 R_bl
Cb_59_55 bit_59_55 gnd C_bl
Cbb_59_55 bitb_59_55 gnd C_bl
Rb_59_56 bit_59_56 bit_59_57 R_bl
Rbb_59_56 bitb_59_56 bitb_59_57 R_bl
Cb_59_56 bit_59_56 gnd C_bl
Cbb_59_56 bitb_59_56 gnd C_bl
Rb_59_57 bit_59_57 bit_59_58 R_bl
Rbb_59_57 bitb_59_57 bitb_59_58 R_bl
Cb_59_57 bit_59_57 gnd C_bl
Cbb_59_57 bitb_59_57 gnd C_bl
Rb_59_58 bit_59_58 bit_59_59 R_bl
Rbb_59_58 bitb_59_58 bitb_59_59 R_bl
Cb_59_58 bit_59_58 gnd C_bl
Cbb_59_58 bitb_59_58 gnd C_bl
Rb_59_59 bit_59_59 bit_59_60 R_bl
Rbb_59_59 bitb_59_59 bitb_59_60 R_bl
Cb_59_59 bit_59_59 gnd C_bl
Cbb_59_59 bitb_59_59 gnd C_bl
Rb_59_60 bit_59_60 bit_59_61 R_bl
Rbb_59_60 bitb_59_60 bitb_59_61 R_bl
Cb_59_60 bit_59_60 gnd C_bl
Cbb_59_60 bitb_59_60 gnd C_bl
Rb_59_61 bit_59_61 bit_59_62 R_bl
Rbb_59_61 bitb_59_61 bitb_59_62 R_bl
Cb_59_61 bit_59_61 gnd C_bl
Cbb_59_61 bitb_59_61 gnd C_bl
Rb_59_62 bit_59_62 bit_59_63 R_bl
Rbb_59_62 bitb_59_62 bitb_59_63 R_bl
Cb_59_62 bit_59_62 gnd C_bl
Cbb_59_62 bitb_59_62 gnd C_bl
Rb_59_63 bit_59_63 bit_59_64 R_bl
Rbb_59_63 bitb_59_63 bitb_59_64 R_bl
Cb_59_63 bit_59_63 gnd C_bl
Cbb_59_63 bitb_59_63 gnd C_bl
Rb_59_64 bit_59_64 bit_59_65 R_bl
Rbb_59_64 bitb_59_64 bitb_59_65 R_bl
Cb_59_64 bit_59_64 gnd C_bl
Cbb_59_64 bitb_59_64 gnd C_bl
Rb_59_65 bit_59_65 bit_59_66 R_bl
Rbb_59_65 bitb_59_65 bitb_59_66 R_bl
Cb_59_65 bit_59_65 gnd C_bl
Cbb_59_65 bitb_59_65 gnd C_bl
Rb_59_66 bit_59_66 bit_59_67 R_bl
Rbb_59_66 bitb_59_66 bitb_59_67 R_bl
Cb_59_66 bit_59_66 gnd C_bl
Cbb_59_66 bitb_59_66 gnd C_bl
Rb_59_67 bit_59_67 bit_59_68 R_bl
Rbb_59_67 bitb_59_67 bitb_59_68 R_bl
Cb_59_67 bit_59_67 gnd C_bl
Cbb_59_67 bitb_59_67 gnd C_bl
Rb_59_68 bit_59_68 bit_59_69 R_bl
Rbb_59_68 bitb_59_68 bitb_59_69 R_bl
Cb_59_68 bit_59_68 gnd C_bl
Cbb_59_68 bitb_59_68 gnd C_bl
Rb_59_69 bit_59_69 bit_59_70 R_bl
Rbb_59_69 bitb_59_69 bitb_59_70 R_bl
Cb_59_69 bit_59_69 gnd C_bl
Cbb_59_69 bitb_59_69 gnd C_bl
Rb_59_70 bit_59_70 bit_59_71 R_bl
Rbb_59_70 bitb_59_70 bitb_59_71 R_bl
Cb_59_70 bit_59_70 gnd C_bl
Cbb_59_70 bitb_59_70 gnd C_bl
Rb_59_71 bit_59_71 bit_59_72 R_bl
Rbb_59_71 bitb_59_71 bitb_59_72 R_bl
Cb_59_71 bit_59_71 gnd C_bl
Cbb_59_71 bitb_59_71 gnd C_bl
Rb_59_72 bit_59_72 bit_59_73 R_bl
Rbb_59_72 bitb_59_72 bitb_59_73 R_bl
Cb_59_72 bit_59_72 gnd C_bl
Cbb_59_72 bitb_59_72 gnd C_bl
Rb_59_73 bit_59_73 bit_59_74 R_bl
Rbb_59_73 bitb_59_73 bitb_59_74 R_bl
Cb_59_73 bit_59_73 gnd C_bl
Cbb_59_73 bitb_59_73 gnd C_bl
Rb_59_74 bit_59_74 bit_59_75 R_bl
Rbb_59_74 bitb_59_74 bitb_59_75 R_bl
Cb_59_74 bit_59_74 gnd C_bl
Cbb_59_74 bitb_59_74 gnd C_bl
Rb_59_75 bit_59_75 bit_59_76 R_bl
Rbb_59_75 bitb_59_75 bitb_59_76 R_bl
Cb_59_75 bit_59_75 gnd C_bl
Cbb_59_75 bitb_59_75 gnd C_bl
Rb_59_76 bit_59_76 bit_59_77 R_bl
Rbb_59_76 bitb_59_76 bitb_59_77 R_bl
Cb_59_76 bit_59_76 gnd C_bl
Cbb_59_76 bitb_59_76 gnd C_bl
Rb_59_77 bit_59_77 bit_59_78 R_bl
Rbb_59_77 bitb_59_77 bitb_59_78 R_bl
Cb_59_77 bit_59_77 gnd C_bl
Cbb_59_77 bitb_59_77 gnd C_bl
Rb_59_78 bit_59_78 bit_59_79 R_bl
Rbb_59_78 bitb_59_78 bitb_59_79 R_bl
Cb_59_78 bit_59_78 gnd C_bl
Cbb_59_78 bitb_59_78 gnd C_bl
Rb_59_79 bit_59_79 bit_59_80 R_bl
Rbb_59_79 bitb_59_79 bitb_59_80 R_bl
Cb_59_79 bit_59_79 gnd C_bl
Cbb_59_79 bitb_59_79 gnd C_bl
Rb_59_80 bit_59_80 bit_59_81 R_bl
Rbb_59_80 bitb_59_80 bitb_59_81 R_bl
Cb_59_80 bit_59_80 gnd C_bl
Cbb_59_80 bitb_59_80 gnd C_bl
Rb_59_81 bit_59_81 bit_59_82 R_bl
Rbb_59_81 bitb_59_81 bitb_59_82 R_bl
Cb_59_81 bit_59_81 gnd C_bl
Cbb_59_81 bitb_59_81 gnd C_bl
Rb_59_82 bit_59_82 bit_59_83 R_bl
Rbb_59_82 bitb_59_82 bitb_59_83 R_bl
Cb_59_82 bit_59_82 gnd C_bl
Cbb_59_82 bitb_59_82 gnd C_bl
Rb_59_83 bit_59_83 bit_59_84 R_bl
Rbb_59_83 bitb_59_83 bitb_59_84 R_bl
Cb_59_83 bit_59_83 gnd C_bl
Cbb_59_83 bitb_59_83 gnd C_bl
Rb_59_84 bit_59_84 bit_59_85 R_bl
Rbb_59_84 bitb_59_84 bitb_59_85 R_bl
Cb_59_84 bit_59_84 gnd C_bl
Cbb_59_84 bitb_59_84 gnd C_bl
Rb_59_85 bit_59_85 bit_59_86 R_bl
Rbb_59_85 bitb_59_85 bitb_59_86 R_bl
Cb_59_85 bit_59_85 gnd C_bl
Cbb_59_85 bitb_59_85 gnd C_bl
Rb_59_86 bit_59_86 bit_59_87 R_bl
Rbb_59_86 bitb_59_86 bitb_59_87 R_bl
Cb_59_86 bit_59_86 gnd C_bl
Cbb_59_86 bitb_59_86 gnd C_bl
Rb_59_87 bit_59_87 bit_59_88 R_bl
Rbb_59_87 bitb_59_87 bitb_59_88 R_bl
Cb_59_87 bit_59_87 gnd C_bl
Cbb_59_87 bitb_59_87 gnd C_bl
Rb_59_88 bit_59_88 bit_59_89 R_bl
Rbb_59_88 bitb_59_88 bitb_59_89 R_bl
Cb_59_88 bit_59_88 gnd C_bl
Cbb_59_88 bitb_59_88 gnd C_bl
Rb_59_89 bit_59_89 bit_59_90 R_bl
Rbb_59_89 bitb_59_89 bitb_59_90 R_bl
Cb_59_89 bit_59_89 gnd C_bl
Cbb_59_89 bitb_59_89 gnd C_bl
Rb_59_90 bit_59_90 bit_59_91 R_bl
Rbb_59_90 bitb_59_90 bitb_59_91 R_bl
Cb_59_90 bit_59_90 gnd C_bl
Cbb_59_90 bitb_59_90 gnd C_bl
Rb_59_91 bit_59_91 bit_59_92 R_bl
Rbb_59_91 bitb_59_91 bitb_59_92 R_bl
Cb_59_91 bit_59_91 gnd C_bl
Cbb_59_91 bitb_59_91 gnd C_bl
Rb_59_92 bit_59_92 bit_59_93 R_bl
Rbb_59_92 bitb_59_92 bitb_59_93 R_bl
Cb_59_92 bit_59_92 gnd C_bl
Cbb_59_92 bitb_59_92 gnd C_bl
Rb_59_93 bit_59_93 bit_59_94 R_bl
Rbb_59_93 bitb_59_93 bitb_59_94 R_bl
Cb_59_93 bit_59_93 gnd C_bl
Cbb_59_93 bitb_59_93 gnd C_bl
Rb_59_94 bit_59_94 bit_59_95 R_bl
Rbb_59_94 bitb_59_94 bitb_59_95 R_bl
Cb_59_94 bit_59_94 gnd C_bl
Cbb_59_94 bitb_59_94 gnd C_bl
Rb_59_95 bit_59_95 bit_59_96 R_bl
Rbb_59_95 bitb_59_95 bitb_59_96 R_bl
Cb_59_95 bit_59_95 gnd C_bl
Cbb_59_95 bitb_59_95 gnd C_bl
Rb_59_96 bit_59_96 bit_59_97 R_bl
Rbb_59_96 bitb_59_96 bitb_59_97 R_bl
Cb_59_96 bit_59_96 gnd C_bl
Cbb_59_96 bitb_59_96 gnd C_bl
Rb_59_97 bit_59_97 bit_59_98 R_bl
Rbb_59_97 bitb_59_97 bitb_59_98 R_bl
Cb_59_97 bit_59_97 gnd C_bl
Cbb_59_97 bitb_59_97 gnd C_bl
Rb_59_98 bit_59_98 bit_59_99 R_bl
Rbb_59_98 bitb_59_98 bitb_59_99 R_bl
Cb_59_98 bit_59_98 gnd C_bl
Cbb_59_98 bitb_59_98 gnd C_bl
Rb_59_99 bit_59_99 bit_59_100 R_bl
Rbb_59_99 bitb_59_99 bitb_59_100 R_bl
Cb_59_99 bit_59_99 gnd C_bl
Cbb_59_99 bitb_59_99 gnd C_bl
Rb_60_0 bit_60_0 bit_60_1 R_bl
Rbb_60_0 bitb_60_0 bitb_60_1 R_bl
Cb_60_0 bit_60_0 gnd C_bl
Cbb_60_0 bitb_60_0 gnd C_bl
Rb_60_1 bit_60_1 bit_60_2 R_bl
Rbb_60_1 bitb_60_1 bitb_60_2 R_bl
Cb_60_1 bit_60_1 gnd C_bl
Cbb_60_1 bitb_60_1 gnd C_bl
Rb_60_2 bit_60_2 bit_60_3 R_bl
Rbb_60_2 bitb_60_2 bitb_60_3 R_bl
Cb_60_2 bit_60_2 gnd C_bl
Cbb_60_2 bitb_60_2 gnd C_bl
Rb_60_3 bit_60_3 bit_60_4 R_bl
Rbb_60_3 bitb_60_3 bitb_60_4 R_bl
Cb_60_3 bit_60_3 gnd C_bl
Cbb_60_3 bitb_60_3 gnd C_bl
Rb_60_4 bit_60_4 bit_60_5 R_bl
Rbb_60_4 bitb_60_4 bitb_60_5 R_bl
Cb_60_4 bit_60_4 gnd C_bl
Cbb_60_4 bitb_60_4 gnd C_bl
Rb_60_5 bit_60_5 bit_60_6 R_bl
Rbb_60_5 bitb_60_5 bitb_60_6 R_bl
Cb_60_5 bit_60_5 gnd C_bl
Cbb_60_5 bitb_60_5 gnd C_bl
Rb_60_6 bit_60_6 bit_60_7 R_bl
Rbb_60_6 bitb_60_6 bitb_60_7 R_bl
Cb_60_6 bit_60_6 gnd C_bl
Cbb_60_6 bitb_60_6 gnd C_bl
Rb_60_7 bit_60_7 bit_60_8 R_bl
Rbb_60_7 bitb_60_7 bitb_60_8 R_bl
Cb_60_7 bit_60_7 gnd C_bl
Cbb_60_7 bitb_60_7 gnd C_bl
Rb_60_8 bit_60_8 bit_60_9 R_bl
Rbb_60_8 bitb_60_8 bitb_60_9 R_bl
Cb_60_8 bit_60_8 gnd C_bl
Cbb_60_8 bitb_60_8 gnd C_bl
Rb_60_9 bit_60_9 bit_60_10 R_bl
Rbb_60_9 bitb_60_9 bitb_60_10 R_bl
Cb_60_9 bit_60_9 gnd C_bl
Cbb_60_9 bitb_60_9 gnd C_bl
Rb_60_10 bit_60_10 bit_60_11 R_bl
Rbb_60_10 bitb_60_10 bitb_60_11 R_bl
Cb_60_10 bit_60_10 gnd C_bl
Cbb_60_10 bitb_60_10 gnd C_bl
Rb_60_11 bit_60_11 bit_60_12 R_bl
Rbb_60_11 bitb_60_11 bitb_60_12 R_bl
Cb_60_11 bit_60_11 gnd C_bl
Cbb_60_11 bitb_60_11 gnd C_bl
Rb_60_12 bit_60_12 bit_60_13 R_bl
Rbb_60_12 bitb_60_12 bitb_60_13 R_bl
Cb_60_12 bit_60_12 gnd C_bl
Cbb_60_12 bitb_60_12 gnd C_bl
Rb_60_13 bit_60_13 bit_60_14 R_bl
Rbb_60_13 bitb_60_13 bitb_60_14 R_bl
Cb_60_13 bit_60_13 gnd C_bl
Cbb_60_13 bitb_60_13 gnd C_bl
Rb_60_14 bit_60_14 bit_60_15 R_bl
Rbb_60_14 bitb_60_14 bitb_60_15 R_bl
Cb_60_14 bit_60_14 gnd C_bl
Cbb_60_14 bitb_60_14 gnd C_bl
Rb_60_15 bit_60_15 bit_60_16 R_bl
Rbb_60_15 bitb_60_15 bitb_60_16 R_bl
Cb_60_15 bit_60_15 gnd C_bl
Cbb_60_15 bitb_60_15 gnd C_bl
Rb_60_16 bit_60_16 bit_60_17 R_bl
Rbb_60_16 bitb_60_16 bitb_60_17 R_bl
Cb_60_16 bit_60_16 gnd C_bl
Cbb_60_16 bitb_60_16 gnd C_bl
Rb_60_17 bit_60_17 bit_60_18 R_bl
Rbb_60_17 bitb_60_17 bitb_60_18 R_bl
Cb_60_17 bit_60_17 gnd C_bl
Cbb_60_17 bitb_60_17 gnd C_bl
Rb_60_18 bit_60_18 bit_60_19 R_bl
Rbb_60_18 bitb_60_18 bitb_60_19 R_bl
Cb_60_18 bit_60_18 gnd C_bl
Cbb_60_18 bitb_60_18 gnd C_bl
Rb_60_19 bit_60_19 bit_60_20 R_bl
Rbb_60_19 bitb_60_19 bitb_60_20 R_bl
Cb_60_19 bit_60_19 gnd C_bl
Cbb_60_19 bitb_60_19 gnd C_bl
Rb_60_20 bit_60_20 bit_60_21 R_bl
Rbb_60_20 bitb_60_20 bitb_60_21 R_bl
Cb_60_20 bit_60_20 gnd C_bl
Cbb_60_20 bitb_60_20 gnd C_bl
Rb_60_21 bit_60_21 bit_60_22 R_bl
Rbb_60_21 bitb_60_21 bitb_60_22 R_bl
Cb_60_21 bit_60_21 gnd C_bl
Cbb_60_21 bitb_60_21 gnd C_bl
Rb_60_22 bit_60_22 bit_60_23 R_bl
Rbb_60_22 bitb_60_22 bitb_60_23 R_bl
Cb_60_22 bit_60_22 gnd C_bl
Cbb_60_22 bitb_60_22 gnd C_bl
Rb_60_23 bit_60_23 bit_60_24 R_bl
Rbb_60_23 bitb_60_23 bitb_60_24 R_bl
Cb_60_23 bit_60_23 gnd C_bl
Cbb_60_23 bitb_60_23 gnd C_bl
Rb_60_24 bit_60_24 bit_60_25 R_bl
Rbb_60_24 bitb_60_24 bitb_60_25 R_bl
Cb_60_24 bit_60_24 gnd C_bl
Cbb_60_24 bitb_60_24 gnd C_bl
Rb_60_25 bit_60_25 bit_60_26 R_bl
Rbb_60_25 bitb_60_25 bitb_60_26 R_bl
Cb_60_25 bit_60_25 gnd C_bl
Cbb_60_25 bitb_60_25 gnd C_bl
Rb_60_26 bit_60_26 bit_60_27 R_bl
Rbb_60_26 bitb_60_26 bitb_60_27 R_bl
Cb_60_26 bit_60_26 gnd C_bl
Cbb_60_26 bitb_60_26 gnd C_bl
Rb_60_27 bit_60_27 bit_60_28 R_bl
Rbb_60_27 bitb_60_27 bitb_60_28 R_bl
Cb_60_27 bit_60_27 gnd C_bl
Cbb_60_27 bitb_60_27 gnd C_bl
Rb_60_28 bit_60_28 bit_60_29 R_bl
Rbb_60_28 bitb_60_28 bitb_60_29 R_bl
Cb_60_28 bit_60_28 gnd C_bl
Cbb_60_28 bitb_60_28 gnd C_bl
Rb_60_29 bit_60_29 bit_60_30 R_bl
Rbb_60_29 bitb_60_29 bitb_60_30 R_bl
Cb_60_29 bit_60_29 gnd C_bl
Cbb_60_29 bitb_60_29 gnd C_bl
Rb_60_30 bit_60_30 bit_60_31 R_bl
Rbb_60_30 bitb_60_30 bitb_60_31 R_bl
Cb_60_30 bit_60_30 gnd C_bl
Cbb_60_30 bitb_60_30 gnd C_bl
Rb_60_31 bit_60_31 bit_60_32 R_bl
Rbb_60_31 bitb_60_31 bitb_60_32 R_bl
Cb_60_31 bit_60_31 gnd C_bl
Cbb_60_31 bitb_60_31 gnd C_bl
Rb_60_32 bit_60_32 bit_60_33 R_bl
Rbb_60_32 bitb_60_32 bitb_60_33 R_bl
Cb_60_32 bit_60_32 gnd C_bl
Cbb_60_32 bitb_60_32 gnd C_bl
Rb_60_33 bit_60_33 bit_60_34 R_bl
Rbb_60_33 bitb_60_33 bitb_60_34 R_bl
Cb_60_33 bit_60_33 gnd C_bl
Cbb_60_33 bitb_60_33 gnd C_bl
Rb_60_34 bit_60_34 bit_60_35 R_bl
Rbb_60_34 bitb_60_34 bitb_60_35 R_bl
Cb_60_34 bit_60_34 gnd C_bl
Cbb_60_34 bitb_60_34 gnd C_bl
Rb_60_35 bit_60_35 bit_60_36 R_bl
Rbb_60_35 bitb_60_35 bitb_60_36 R_bl
Cb_60_35 bit_60_35 gnd C_bl
Cbb_60_35 bitb_60_35 gnd C_bl
Rb_60_36 bit_60_36 bit_60_37 R_bl
Rbb_60_36 bitb_60_36 bitb_60_37 R_bl
Cb_60_36 bit_60_36 gnd C_bl
Cbb_60_36 bitb_60_36 gnd C_bl
Rb_60_37 bit_60_37 bit_60_38 R_bl
Rbb_60_37 bitb_60_37 bitb_60_38 R_bl
Cb_60_37 bit_60_37 gnd C_bl
Cbb_60_37 bitb_60_37 gnd C_bl
Rb_60_38 bit_60_38 bit_60_39 R_bl
Rbb_60_38 bitb_60_38 bitb_60_39 R_bl
Cb_60_38 bit_60_38 gnd C_bl
Cbb_60_38 bitb_60_38 gnd C_bl
Rb_60_39 bit_60_39 bit_60_40 R_bl
Rbb_60_39 bitb_60_39 bitb_60_40 R_bl
Cb_60_39 bit_60_39 gnd C_bl
Cbb_60_39 bitb_60_39 gnd C_bl
Rb_60_40 bit_60_40 bit_60_41 R_bl
Rbb_60_40 bitb_60_40 bitb_60_41 R_bl
Cb_60_40 bit_60_40 gnd C_bl
Cbb_60_40 bitb_60_40 gnd C_bl
Rb_60_41 bit_60_41 bit_60_42 R_bl
Rbb_60_41 bitb_60_41 bitb_60_42 R_bl
Cb_60_41 bit_60_41 gnd C_bl
Cbb_60_41 bitb_60_41 gnd C_bl
Rb_60_42 bit_60_42 bit_60_43 R_bl
Rbb_60_42 bitb_60_42 bitb_60_43 R_bl
Cb_60_42 bit_60_42 gnd C_bl
Cbb_60_42 bitb_60_42 gnd C_bl
Rb_60_43 bit_60_43 bit_60_44 R_bl
Rbb_60_43 bitb_60_43 bitb_60_44 R_bl
Cb_60_43 bit_60_43 gnd C_bl
Cbb_60_43 bitb_60_43 gnd C_bl
Rb_60_44 bit_60_44 bit_60_45 R_bl
Rbb_60_44 bitb_60_44 bitb_60_45 R_bl
Cb_60_44 bit_60_44 gnd C_bl
Cbb_60_44 bitb_60_44 gnd C_bl
Rb_60_45 bit_60_45 bit_60_46 R_bl
Rbb_60_45 bitb_60_45 bitb_60_46 R_bl
Cb_60_45 bit_60_45 gnd C_bl
Cbb_60_45 bitb_60_45 gnd C_bl
Rb_60_46 bit_60_46 bit_60_47 R_bl
Rbb_60_46 bitb_60_46 bitb_60_47 R_bl
Cb_60_46 bit_60_46 gnd C_bl
Cbb_60_46 bitb_60_46 gnd C_bl
Rb_60_47 bit_60_47 bit_60_48 R_bl
Rbb_60_47 bitb_60_47 bitb_60_48 R_bl
Cb_60_47 bit_60_47 gnd C_bl
Cbb_60_47 bitb_60_47 gnd C_bl
Rb_60_48 bit_60_48 bit_60_49 R_bl
Rbb_60_48 bitb_60_48 bitb_60_49 R_bl
Cb_60_48 bit_60_48 gnd C_bl
Cbb_60_48 bitb_60_48 gnd C_bl
Rb_60_49 bit_60_49 bit_60_50 R_bl
Rbb_60_49 bitb_60_49 bitb_60_50 R_bl
Cb_60_49 bit_60_49 gnd C_bl
Cbb_60_49 bitb_60_49 gnd C_bl
Rb_60_50 bit_60_50 bit_60_51 R_bl
Rbb_60_50 bitb_60_50 bitb_60_51 R_bl
Cb_60_50 bit_60_50 gnd C_bl
Cbb_60_50 bitb_60_50 gnd C_bl
Rb_60_51 bit_60_51 bit_60_52 R_bl
Rbb_60_51 bitb_60_51 bitb_60_52 R_bl
Cb_60_51 bit_60_51 gnd C_bl
Cbb_60_51 bitb_60_51 gnd C_bl
Rb_60_52 bit_60_52 bit_60_53 R_bl
Rbb_60_52 bitb_60_52 bitb_60_53 R_bl
Cb_60_52 bit_60_52 gnd C_bl
Cbb_60_52 bitb_60_52 gnd C_bl
Rb_60_53 bit_60_53 bit_60_54 R_bl
Rbb_60_53 bitb_60_53 bitb_60_54 R_bl
Cb_60_53 bit_60_53 gnd C_bl
Cbb_60_53 bitb_60_53 gnd C_bl
Rb_60_54 bit_60_54 bit_60_55 R_bl
Rbb_60_54 bitb_60_54 bitb_60_55 R_bl
Cb_60_54 bit_60_54 gnd C_bl
Cbb_60_54 bitb_60_54 gnd C_bl
Rb_60_55 bit_60_55 bit_60_56 R_bl
Rbb_60_55 bitb_60_55 bitb_60_56 R_bl
Cb_60_55 bit_60_55 gnd C_bl
Cbb_60_55 bitb_60_55 gnd C_bl
Rb_60_56 bit_60_56 bit_60_57 R_bl
Rbb_60_56 bitb_60_56 bitb_60_57 R_bl
Cb_60_56 bit_60_56 gnd C_bl
Cbb_60_56 bitb_60_56 gnd C_bl
Rb_60_57 bit_60_57 bit_60_58 R_bl
Rbb_60_57 bitb_60_57 bitb_60_58 R_bl
Cb_60_57 bit_60_57 gnd C_bl
Cbb_60_57 bitb_60_57 gnd C_bl
Rb_60_58 bit_60_58 bit_60_59 R_bl
Rbb_60_58 bitb_60_58 bitb_60_59 R_bl
Cb_60_58 bit_60_58 gnd C_bl
Cbb_60_58 bitb_60_58 gnd C_bl
Rb_60_59 bit_60_59 bit_60_60 R_bl
Rbb_60_59 bitb_60_59 bitb_60_60 R_bl
Cb_60_59 bit_60_59 gnd C_bl
Cbb_60_59 bitb_60_59 gnd C_bl
Rb_60_60 bit_60_60 bit_60_61 R_bl
Rbb_60_60 bitb_60_60 bitb_60_61 R_bl
Cb_60_60 bit_60_60 gnd C_bl
Cbb_60_60 bitb_60_60 gnd C_bl
Rb_60_61 bit_60_61 bit_60_62 R_bl
Rbb_60_61 bitb_60_61 bitb_60_62 R_bl
Cb_60_61 bit_60_61 gnd C_bl
Cbb_60_61 bitb_60_61 gnd C_bl
Rb_60_62 bit_60_62 bit_60_63 R_bl
Rbb_60_62 bitb_60_62 bitb_60_63 R_bl
Cb_60_62 bit_60_62 gnd C_bl
Cbb_60_62 bitb_60_62 gnd C_bl
Rb_60_63 bit_60_63 bit_60_64 R_bl
Rbb_60_63 bitb_60_63 bitb_60_64 R_bl
Cb_60_63 bit_60_63 gnd C_bl
Cbb_60_63 bitb_60_63 gnd C_bl
Rb_60_64 bit_60_64 bit_60_65 R_bl
Rbb_60_64 bitb_60_64 bitb_60_65 R_bl
Cb_60_64 bit_60_64 gnd C_bl
Cbb_60_64 bitb_60_64 gnd C_bl
Rb_60_65 bit_60_65 bit_60_66 R_bl
Rbb_60_65 bitb_60_65 bitb_60_66 R_bl
Cb_60_65 bit_60_65 gnd C_bl
Cbb_60_65 bitb_60_65 gnd C_bl
Rb_60_66 bit_60_66 bit_60_67 R_bl
Rbb_60_66 bitb_60_66 bitb_60_67 R_bl
Cb_60_66 bit_60_66 gnd C_bl
Cbb_60_66 bitb_60_66 gnd C_bl
Rb_60_67 bit_60_67 bit_60_68 R_bl
Rbb_60_67 bitb_60_67 bitb_60_68 R_bl
Cb_60_67 bit_60_67 gnd C_bl
Cbb_60_67 bitb_60_67 gnd C_bl
Rb_60_68 bit_60_68 bit_60_69 R_bl
Rbb_60_68 bitb_60_68 bitb_60_69 R_bl
Cb_60_68 bit_60_68 gnd C_bl
Cbb_60_68 bitb_60_68 gnd C_bl
Rb_60_69 bit_60_69 bit_60_70 R_bl
Rbb_60_69 bitb_60_69 bitb_60_70 R_bl
Cb_60_69 bit_60_69 gnd C_bl
Cbb_60_69 bitb_60_69 gnd C_bl
Rb_60_70 bit_60_70 bit_60_71 R_bl
Rbb_60_70 bitb_60_70 bitb_60_71 R_bl
Cb_60_70 bit_60_70 gnd C_bl
Cbb_60_70 bitb_60_70 gnd C_bl
Rb_60_71 bit_60_71 bit_60_72 R_bl
Rbb_60_71 bitb_60_71 bitb_60_72 R_bl
Cb_60_71 bit_60_71 gnd C_bl
Cbb_60_71 bitb_60_71 gnd C_bl
Rb_60_72 bit_60_72 bit_60_73 R_bl
Rbb_60_72 bitb_60_72 bitb_60_73 R_bl
Cb_60_72 bit_60_72 gnd C_bl
Cbb_60_72 bitb_60_72 gnd C_bl
Rb_60_73 bit_60_73 bit_60_74 R_bl
Rbb_60_73 bitb_60_73 bitb_60_74 R_bl
Cb_60_73 bit_60_73 gnd C_bl
Cbb_60_73 bitb_60_73 gnd C_bl
Rb_60_74 bit_60_74 bit_60_75 R_bl
Rbb_60_74 bitb_60_74 bitb_60_75 R_bl
Cb_60_74 bit_60_74 gnd C_bl
Cbb_60_74 bitb_60_74 gnd C_bl
Rb_60_75 bit_60_75 bit_60_76 R_bl
Rbb_60_75 bitb_60_75 bitb_60_76 R_bl
Cb_60_75 bit_60_75 gnd C_bl
Cbb_60_75 bitb_60_75 gnd C_bl
Rb_60_76 bit_60_76 bit_60_77 R_bl
Rbb_60_76 bitb_60_76 bitb_60_77 R_bl
Cb_60_76 bit_60_76 gnd C_bl
Cbb_60_76 bitb_60_76 gnd C_bl
Rb_60_77 bit_60_77 bit_60_78 R_bl
Rbb_60_77 bitb_60_77 bitb_60_78 R_bl
Cb_60_77 bit_60_77 gnd C_bl
Cbb_60_77 bitb_60_77 gnd C_bl
Rb_60_78 bit_60_78 bit_60_79 R_bl
Rbb_60_78 bitb_60_78 bitb_60_79 R_bl
Cb_60_78 bit_60_78 gnd C_bl
Cbb_60_78 bitb_60_78 gnd C_bl
Rb_60_79 bit_60_79 bit_60_80 R_bl
Rbb_60_79 bitb_60_79 bitb_60_80 R_bl
Cb_60_79 bit_60_79 gnd C_bl
Cbb_60_79 bitb_60_79 gnd C_bl
Rb_60_80 bit_60_80 bit_60_81 R_bl
Rbb_60_80 bitb_60_80 bitb_60_81 R_bl
Cb_60_80 bit_60_80 gnd C_bl
Cbb_60_80 bitb_60_80 gnd C_bl
Rb_60_81 bit_60_81 bit_60_82 R_bl
Rbb_60_81 bitb_60_81 bitb_60_82 R_bl
Cb_60_81 bit_60_81 gnd C_bl
Cbb_60_81 bitb_60_81 gnd C_bl
Rb_60_82 bit_60_82 bit_60_83 R_bl
Rbb_60_82 bitb_60_82 bitb_60_83 R_bl
Cb_60_82 bit_60_82 gnd C_bl
Cbb_60_82 bitb_60_82 gnd C_bl
Rb_60_83 bit_60_83 bit_60_84 R_bl
Rbb_60_83 bitb_60_83 bitb_60_84 R_bl
Cb_60_83 bit_60_83 gnd C_bl
Cbb_60_83 bitb_60_83 gnd C_bl
Rb_60_84 bit_60_84 bit_60_85 R_bl
Rbb_60_84 bitb_60_84 bitb_60_85 R_bl
Cb_60_84 bit_60_84 gnd C_bl
Cbb_60_84 bitb_60_84 gnd C_bl
Rb_60_85 bit_60_85 bit_60_86 R_bl
Rbb_60_85 bitb_60_85 bitb_60_86 R_bl
Cb_60_85 bit_60_85 gnd C_bl
Cbb_60_85 bitb_60_85 gnd C_bl
Rb_60_86 bit_60_86 bit_60_87 R_bl
Rbb_60_86 bitb_60_86 bitb_60_87 R_bl
Cb_60_86 bit_60_86 gnd C_bl
Cbb_60_86 bitb_60_86 gnd C_bl
Rb_60_87 bit_60_87 bit_60_88 R_bl
Rbb_60_87 bitb_60_87 bitb_60_88 R_bl
Cb_60_87 bit_60_87 gnd C_bl
Cbb_60_87 bitb_60_87 gnd C_bl
Rb_60_88 bit_60_88 bit_60_89 R_bl
Rbb_60_88 bitb_60_88 bitb_60_89 R_bl
Cb_60_88 bit_60_88 gnd C_bl
Cbb_60_88 bitb_60_88 gnd C_bl
Rb_60_89 bit_60_89 bit_60_90 R_bl
Rbb_60_89 bitb_60_89 bitb_60_90 R_bl
Cb_60_89 bit_60_89 gnd C_bl
Cbb_60_89 bitb_60_89 gnd C_bl
Rb_60_90 bit_60_90 bit_60_91 R_bl
Rbb_60_90 bitb_60_90 bitb_60_91 R_bl
Cb_60_90 bit_60_90 gnd C_bl
Cbb_60_90 bitb_60_90 gnd C_bl
Rb_60_91 bit_60_91 bit_60_92 R_bl
Rbb_60_91 bitb_60_91 bitb_60_92 R_bl
Cb_60_91 bit_60_91 gnd C_bl
Cbb_60_91 bitb_60_91 gnd C_bl
Rb_60_92 bit_60_92 bit_60_93 R_bl
Rbb_60_92 bitb_60_92 bitb_60_93 R_bl
Cb_60_92 bit_60_92 gnd C_bl
Cbb_60_92 bitb_60_92 gnd C_bl
Rb_60_93 bit_60_93 bit_60_94 R_bl
Rbb_60_93 bitb_60_93 bitb_60_94 R_bl
Cb_60_93 bit_60_93 gnd C_bl
Cbb_60_93 bitb_60_93 gnd C_bl
Rb_60_94 bit_60_94 bit_60_95 R_bl
Rbb_60_94 bitb_60_94 bitb_60_95 R_bl
Cb_60_94 bit_60_94 gnd C_bl
Cbb_60_94 bitb_60_94 gnd C_bl
Rb_60_95 bit_60_95 bit_60_96 R_bl
Rbb_60_95 bitb_60_95 bitb_60_96 R_bl
Cb_60_95 bit_60_95 gnd C_bl
Cbb_60_95 bitb_60_95 gnd C_bl
Rb_60_96 bit_60_96 bit_60_97 R_bl
Rbb_60_96 bitb_60_96 bitb_60_97 R_bl
Cb_60_96 bit_60_96 gnd C_bl
Cbb_60_96 bitb_60_96 gnd C_bl
Rb_60_97 bit_60_97 bit_60_98 R_bl
Rbb_60_97 bitb_60_97 bitb_60_98 R_bl
Cb_60_97 bit_60_97 gnd C_bl
Cbb_60_97 bitb_60_97 gnd C_bl
Rb_60_98 bit_60_98 bit_60_99 R_bl
Rbb_60_98 bitb_60_98 bitb_60_99 R_bl
Cb_60_98 bit_60_98 gnd C_bl
Cbb_60_98 bitb_60_98 gnd C_bl
Rb_60_99 bit_60_99 bit_60_100 R_bl
Rbb_60_99 bitb_60_99 bitb_60_100 R_bl
Cb_60_99 bit_60_99 gnd C_bl
Cbb_60_99 bitb_60_99 gnd C_bl
Rb_61_0 bit_61_0 bit_61_1 R_bl
Rbb_61_0 bitb_61_0 bitb_61_1 R_bl
Cb_61_0 bit_61_0 gnd C_bl
Cbb_61_0 bitb_61_0 gnd C_bl
Rb_61_1 bit_61_1 bit_61_2 R_bl
Rbb_61_1 bitb_61_1 bitb_61_2 R_bl
Cb_61_1 bit_61_1 gnd C_bl
Cbb_61_1 bitb_61_1 gnd C_bl
Rb_61_2 bit_61_2 bit_61_3 R_bl
Rbb_61_2 bitb_61_2 bitb_61_3 R_bl
Cb_61_2 bit_61_2 gnd C_bl
Cbb_61_2 bitb_61_2 gnd C_bl
Rb_61_3 bit_61_3 bit_61_4 R_bl
Rbb_61_3 bitb_61_3 bitb_61_4 R_bl
Cb_61_3 bit_61_3 gnd C_bl
Cbb_61_3 bitb_61_3 gnd C_bl
Rb_61_4 bit_61_4 bit_61_5 R_bl
Rbb_61_4 bitb_61_4 bitb_61_5 R_bl
Cb_61_4 bit_61_4 gnd C_bl
Cbb_61_4 bitb_61_4 gnd C_bl
Rb_61_5 bit_61_5 bit_61_6 R_bl
Rbb_61_5 bitb_61_5 bitb_61_6 R_bl
Cb_61_5 bit_61_5 gnd C_bl
Cbb_61_5 bitb_61_5 gnd C_bl
Rb_61_6 bit_61_6 bit_61_7 R_bl
Rbb_61_6 bitb_61_6 bitb_61_7 R_bl
Cb_61_6 bit_61_6 gnd C_bl
Cbb_61_6 bitb_61_6 gnd C_bl
Rb_61_7 bit_61_7 bit_61_8 R_bl
Rbb_61_7 bitb_61_7 bitb_61_8 R_bl
Cb_61_7 bit_61_7 gnd C_bl
Cbb_61_7 bitb_61_7 gnd C_bl
Rb_61_8 bit_61_8 bit_61_9 R_bl
Rbb_61_8 bitb_61_8 bitb_61_9 R_bl
Cb_61_8 bit_61_8 gnd C_bl
Cbb_61_8 bitb_61_8 gnd C_bl
Rb_61_9 bit_61_9 bit_61_10 R_bl
Rbb_61_9 bitb_61_9 bitb_61_10 R_bl
Cb_61_9 bit_61_9 gnd C_bl
Cbb_61_9 bitb_61_9 gnd C_bl
Rb_61_10 bit_61_10 bit_61_11 R_bl
Rbb_61_10 bitb_61_10 bitb_61_11 R_bl
Cb_61_10 bit_61_10 gnd C_bl
Cbb_61_10 bitb_61_10 gnd C_bl
Rb_61_11 bit_61_11 bit_61_12 R_bl
Rbb_61_11 bitb_61_11 bitb_61_12 R_bl
Cb_61_11 bit_61_11 gnd C_bl
Cbb_61_11 bitb_61_11 gnd C_bl
Rb_61_12 bit_61_12 bit_61_13 R_bl
Rbb_61_12 bitb_61_12 bitb_61_13 R_bl
Cb_61_12 bit_61_12 gnd C_bl
Cbb_61_12 bitb_61_12 gnd C_bl
Rb_61_13 bit_61_13 bit_61_14 R_bl
Rbb_61_13 bitb_61_13 bitb_61_14 R_bl
Cb_61_13 bit_61_13 gnd C_bl
Cbb_61_13 bitb_61_13 gnd C_bl
Rb_61_14 bit_61_14 bit_61_15 R_bl
Rbb_61_14 bitb_61_14 bitb_61_15 R_bl
Cb_61_14 bit_61_14 gnd C_bl
Cbb_61_14 bitb_61_14 gnd C_bl
Rb_61_15 bit_61_15 bit_61_16 R_bl
Rbb_61_15 bitb_61_15 bitb_61_16 R_bl
Cb_61_15 bit_61_15 gnd C_bl
Cbb_61_15 bitb_61_15 gnd C_bl
Rb_61_16 bit_61_16 bit_61_17 R_bl
Rbb_61_16 bitb_61_16 bitb_61_17 R_bl
Cb_61_16 bit_61_16 gnd C_bl
Cbb_61_16 bitb_61_16 gnd C_bl
Rb_61_17 bit_61_17 bit_61_18 R_bl
Rbb_61_17 bitb_61_17 bitb_61_18 R_bl
Cb_61_17 bit_61_17 gnd C_bl
Cbb_61_17 bitb_61_17 gnd C_bl
Rb_61_18 bit_61_18 bit_61_19 R_bl
Rbb_61_18 bitb_61_18 bitb_61_19 R_bl
Cb_61_18 bit_61_18 gnd C_bl
Cbb_61_18 bitb_61_18 gnd C_bl
Rb_61_19 bit_61_19 bit_61_20 R_bl
Rbb_61_19 bitb_61_19 bitb_61_20 R_bl
Cb_61_19 bit_61_19 gnd C_bl
Cbb_61_19 bitb_61_19 gnd C_bl
Rb_61_20 bit_61_20 bit_61_21 R_bl
Rbb_61_20 bitb_61_20 bitb_61_21 R_bl
Cb_61_20 bit_61_20 gnd C_bl
Cbb_61_20 bitb_61_20 gnd C_bl
Rb_61_21 bit_61_21 bit_61_22 R_bl
Rbb_61_21 bitb_61_21 bitb_61_22 R_bl
Cb_61_21 bit_61_21 gnd C_bl
Cbb_61_21 bitb_61_21 gnd C_bl
Rb_61_22 bit_61_22 bit_61_23 R_bl
Rbb_61_22 bitb_61_22 bitb_61_23 R_bl
Cb_61_22 bit_61_22 gnd C_bl
Cbb_61_22 bitb_61_22 gnd C_bl
Rb_61_23 bit_61_23 bit_61_24 R_bl
Rbb_61_23 bitb_61_23 bitb_61_24 R_bl
Cb_61_23 bit_61_23 gnd C_bl
Cbb_61_23 bitb_61_23 gnd C_bl
Rb_61_24 bit_61_24 bit_61_25 R_bl
Rbb_61_24 bitb_61_24 bitb_61_25 R_bl
Cb_61_24 bit_61_24 gnd C_bl
Cbb_61_24 bitb_61_24 gnd C_bl
Rb_61_25 bit_61_25 bit_61_26 R_bl
Rbb_61_25 bitb_61_25 bitb_61_26 R_bl
Cb_61_25 bit_61_25 gnd C_bl
Cbb_61_25 bitb_61_25 gnd C_bl
Rb_61_26 bit_61_26 bit_61_27 R_bl
Rbb_61_26 bitb_61_26 bitb_61_27 R_bl
Cb_61_26 bit_61_26 gnd C_bl
Cbb_61_26 bitb_61_26 gnd C_bl
Rb_61_27 bit_61_27 bit_61_28 R_bl
Rbb_61_27 bitb_61_27 bitb_61_28 R_bl
Cb_61_27 bit_61_27 gnd C_bl
Cbb_61_27 bitb_61_27 gnd C_bl
Rb_61_28 bit_61_28 bit_61_29 R_bl
Rbb_61_28 bitb_61_28 bitb_61_29 R_bl
Cb_61_28 bit_61_28 gnd C_bl
Cbb_61_28 bitb_61_28 gnd C_bl
Rb_61_29 bit_61_29 bit_61_30 R_bl
Rbb_61_29 bitb_61_29 bitb_61_30 R_bl
Cb_61_29 bit_61_29 gnd C_bl
Cbb_61_29 bitb_61_29 gnd C_bl
Rb_61_30 bit_61_30 bit_61_31 R_bl
Rbb_61_30 bitb_61_30 bitb_61_31 R_bl
Cb_61_30 bit_61_30 gnd C_bl
Cbb_61_30 bitb_61_30 gnd C_bl
Rb_61_31 bit_61_31 bit_61_32 R_bl
Rbb_61_31 bitb_61_31 bitb_61_32 R_bl
Cb_61_31 bit_61_31 gnd C_bl
Cbb_61_31 bitb_61_31 gnd C_bl
Rb_61_32 bit_61_32 bit_61_33 R_bl
Rbb_61_32 bitb_61_32 bitb_61_33 R_bl
Cb_61_32 bit_61_32 gnd C_bl
Cbb_61_32 bitb_61_32 gnd C_bl
Rb_61_33 bit_61_33 bit_61_34 R_bl
Rbb_61_33 bitb_61_33 bitb_61_34 R_bl
Cb_61_33 bit_61_33 gnd C_bl
Cbb_61_33 bitb_61_33 gnd C_bl
Rb_61_34 bit_61_34 bit_61_35 R_bl
Rbb_61_34 bitb_61_34 bitb_61_35 R_bl
Cb_61_34 bit_61_34 gnd C_bl
Cbb_61_34 bitb_61_34 gnd C_bl
Rb_61_35 bit_61_35 bit_61_36 R_bl
Rbb_61_35 bitb_61_35 bitb_61_36 R_bl
Cb_61_35 bit_61_35 gnd C_bl
Cbb_61_35 bitb_61_35 gnd C_bl
Rb_61_36 bit_61_36 bit_61_37 R_bl
Rbb_61_36 bitb_61_36 bitb_61_37 R_bl
Cb_61_36 bit_61_36 gnd C_bl
Cbb_61_36 bitb_61_36 gnd C_bl
Rb_61_37 bit_61_37 bit_61_38 R_bl
Rbb_61_37 bitb_61_37 bitb_61_38 R_bl
Cb_61_37 bit_61_37 gnd C_bl
Cbb_61_37 bitb_61_37 gnd C_bl
Rb_61_38 bit_61_38 bit_61_39 R_bl
Rbb_61_38 bitb_61_38 bitb_61_39 R_bl
Cb_61_38 bit_61_38 gnd C_bl
Cbb_61_38 bitb_61_38 gnd C_bl
Rb_61_39 bit_61_39 bit_61_40 R_bl
Rbb_61_39 bitb_61_39 bitb_61_40 R_bl
Cb_61_39 bit_61_39 gnd C_bl
Cbb_61_39 bitb_61_39 gnd C_bl
Rb_61_40 bit_61_40 bit_61_41 R_bl
Rbb_61_40 bitb_61_40 bitb_61_41 R_bl
Cb_61_40 bit_61_40 gnd C_bl
Cbb_61_40 bitb_61_40 gnd C_bl
Rb_61_41 bit_61_41 bit_61_42 R_bl
Rbb_61_41 bitb_61_41 bitb_61_42 R_bl
Cb_61_41 bit_61_41 gnd C_bl
Cbb_61_41 bitb_61_41 gnd C_bl
Rb_61_42 bit_61_42 bit_61_43 R_bl
Rbb_61_42 bitb_61_42 bitb_61_43 R_bl
Cb_61_42 bit_61_42 gnd C_bl
Cbb_61_42 bitb_61_42 gnd C_bl
Rb_61_43 bit_61_43 bit_61_44 R_bl
Rbb_61_43 bitb_61_43 bitb_61_44 R_bl
Cb_61_43 bit_61_43 gnd C_bl
Cbb_61_43 bitb_61_43 gnd C_bl
Rb_61_44 bit_61_44 bit_61_45 R_bl
Rbb_61_44 bitb_61_44 bitb_61_45 R_bl
Cb_61_44 bit_61_44 gnd C_bl
Cbb_61_44 bitb_61_44 gnd C_bl
Rb_61_45 bit_61_45 bit_61_46 R_bl
Rbb_61_45 bitb_61_45 bitb_61_46 R_bl
Cb_61_45 bit_61_45 gnd C_bl
Cbb_61_45 bitb_61_45 gnd C_bl
Rb_61_46 bit_61_46 bit_61_47 R_bl
Rbb_61_46 bitb_61_46 bitb_61_47 R_bl
Cb_61_46 bit_61_46 gnd C_bl
Cbb_61_46 bitb_61_46 gnd C_bl
Rb_61_47 bit_61_47 bit_61_48 R_bl
Rbb_61_47 bitb_61_47 bitb_61_48 R_bl
Cb_61_47 bit_61_47 gnd C_bl
Cbb_61_47 bitb_61_47 gnd C_bl
Rb_61_48 bit_61_48 bit_61_49 R_bl
Rbb_61_48 bitb_61_48 bitb_61_49 R_bl
Cb_61_48 bit_61_48 gnd C_bl
Cbb_61_48 bitb_61_48 gnd C_bl
Rb_61_49 bit_61_49 bit_61_50 R_bl
Rbb_61_49 bitb_61_49 bitb_61_50 R_bl
Cb_61_49 bit_61_49 gnd C_bl
Cbb_61_49 bitb_61_49 gnd C_bl
Rb_61_50 bit_61_50 bit_61_51 R_bl
Rbb_61_50 bitb_61_50 bitb_61_51 R_bl
Cb_61_50 bit_61_50 gnd C_bl
Cbb_61_50 bitb_61_50 gnd C_bl
Rb_61_51 bit_61_51 bit_61_52 R_bl
Rbb_61_51 bitb_61_51 bitb_61_52 R_bl
Cb_61_51 bit_61_51 gnd C_bl
Cbb_61_51 bitb_61_51 gnd C_bl
Rb_61_52 bit_61_52 bit_61_53 R_bl
Rbb_61_52 bitb_61_52 bitb_61_53 R_bl
Cb_61_52 bit_61_52 gnd C_bl
Cbb_61_52 bitb_61_52 gnd C_bl
Rb_61_53 bit_61_53 bit_61_54 R_bl
Rbb_61_53 bitb_61_53 bitb_61_54 R_bl
Cb_61_53 bit_61_53 gnd C_bl
Cbb_61_53 bitb_61_53 gnd C_bl
Rb_61_54 bit_61_54 bit_61_55 R_bl
Rbb_61_54 bitb_61_54 bitb_61_55 R_bl
Cb_61_54 bit_61_54 gnd C_bl
Cbb_61_54 bitb_61_54 gnd C_bl
Rb_61_55 bit_61_55 bit_61_56 R_bl
Rbb_61_55 bitb_61_55 bitb_61_56 R_bl
Cb_61_55 bit_61_55 gnd C_bl
Cbb_61_55 bitb_61_55 gnd C_bl
Rb_61_56 bit_61_56 bit_61_57 R_bl
Rbb_61_56 bitb_61_56 bitb_61_57 R_bl
Cb_61_56 bit_61_56 gnd C_bl
Cbb_61_56 bitb_61_56 gnd C_bl
Rb_61_57 bit_61_57 bit_61_58 R_bl
Rbb_61_57 bitb_61_57 bitb_61_58 R_bl
Cb_61_57 bit_61_57 gnd C_bl
Cbb_61_57 bitb_61_57 gnd C_bl
Rb_61_58 bit_61_58 bit_61_59 R_bl
Rbb_61_58 bitb_61_58 bitb_61_59 R_bl
Cb_61_58 bit_61_58 gnd C_bl
Cbb_61_58 bitb_61_58 gnd C_bl
Rb_61_59 bit_61_59 bit_61_60 R_bl
Rbb_61_59 bitb_61_59 bitb_61_60 R_bl
Cb_61_59 bit_61_59 gnd C_bl
Cbb_61_59 bitb_61_59 gnd C_bl
Rb_61_60 bit_61_60 bit_61_61 R_bl
Rbb_61_60 bitb_61_60 bitb_61_61 R_bl
Cb_61_60 bit_61_60 gnd C_bl
Cbb_61_60 bitb_61_60 gnd C_bl
Rb_61_61 bit_61_61 bit_61_62 R_bl
Rbb_61_61 bitb_61_61 bitb_61_62 R_bl
Cb_61_61 bit_61_61 gnd C_bl
Cbb_61_61 bitb_61_61 gnd C_bl
Rb_61_62 bit_61_62 bit_61_63 R_bl
Rbb_61_62 bitb_61_62 bitb_61_63 R_bl
Cb_61_62 bit_61_62 gnd C_bl
Cbb_61_62 bitb_61_62 gnd C_bl
Rb_61_63 bit_61_63 bit_61_64 R_bl
Rbb_61_63 bitb_61_63 bitb_61_64 R_bl
Cb_61_63 bit_61_63 gnd C_bl
Cbb_61_63 bitb_61_63 gnd C_bl
Rb_61_64 bit_61_64 bit_61_65 R_bl
Rbb_61_64 bitb_61_64 bitb_61_65 R_bl
Cb_61_64 bit_61_64 gnd C_bl
Cbb_61_64 bitb_61_64 gnd C_bl
Rb_61_65 bit_61_65 bit_61_66 R_bl
Rbb_61_65 bitb_61_65 bitb_61_66 R_bl
Cb_61_65 bit_61_65 gnd C_bl
Cbb_61_65 bitb_61_65 gnd C_bl
Rb_61_66 bit_61_66 bit_61_67 R_bl
Rbb_61_66 bitb_61_66 bitb_61_67 R_bl
Cb_61_66 bit_61_66 gnd C_bl
Cbb_61_66 bitb_61_66 gnd C_bl
Rb_61_67 bit_61_67 bit_61_68 R_bl
Rbb_61_67 bitb_61_67 bitb_61_68 R_bl
Cb_61_67 bit_61_67 gnd C_bl
Cbb_61_67 bitb_61_67 gnd C_bl
Rb_61_68 bit_61_68 bit_61_69 R_bl
Rbb_61_68 bitb_61_68 bitb_61_69 R_bl
Cb_61_68 bit_61_68 gnd C_bl
Cbb_61_68 bitb_61_68 gnd C_bl
Rb_61_69 bit_61_69 bit_61_70 R_bl
Rbb_61_69 bitb_61_69 bitb_61_70 R_bl
Cb_61_69 bit_61_69 gnd C_bl
Cbb_61_69 bitb_61_69 gnd C_bl
Rb_61_70 bit_61_70 bit_61_71 R_bl
Rbb_61_70 bitb_61_70 bitb_61_71 R_bl
Cb_61_70 bit_61_70 gnd C_bl
Cbb_61_70 bitb_61_70 gnd C_bl
Rb_61_71 bit_61_71 bit_61_72 R_bl
Rbb_61_71 bitb_61_71 bitb_61_72 R_bl
Cb_61_71 bit_61_71 gnd C_bl
Cbb_61_71 bitb_61_71 gnd C_bl
Rb_61_72 bit_61_72 bit_61_73 R_bl
Rbb_61_72 bitb_61_72 bitb_61_73 R_bl
Cb_61_72 bit_61_72 gnd C_bl
Cbb_61_72 bitb_61_72 gnd C_bl
Rb_61_73 bit_61_73 bit_61_74 R_bl
Rbb_61_73 bitb_61_73 bitb_61_74 R_bl
Cb_61_73 bit_61_73 gnd C_bl
Cbb_61_73 bitb_61_73 gnd C_bl
Rb_61_74 bit_61_74 bit_61_75 R_bl
Rbb_61_74 bitb_61_74 bitb_61_75 R_bl
Cb_61_74 bit_61_74 gnd C_bl
Cbb_61_74 bitb_61_74 gnd C_bl
Rb_61_75 bit_61_75 bit_61_76 R_bl
Rbb_61_75 bitb_61_75 bitb_61_76 R_bl
Cb_61_75 bit_61_75 gnd C_bl
Cbb_61_75 bitb_61_75 gnd C_bl
Rb_61_76 bit_61_76 bit_61_77 R_bl
Rbb_61_76 bitb_61_76 bitb_61_77 R_bl
Cb_61_76 bit_61_76 gnd C_bl
Cbb_61_76 bitb_61_76 gnd C_bl
Rb_61_77 bit_61_77 bit_61_78 R_bl
Rbb_61_77 bitb_61_77 bitb_61_78 R_bl
Cb_61_77 bit_61_77 gnd C_bl
Cbb_61_77 bitb_61_77 gnd C_bl
Rb_61_78 bit_61_78 bit_61_79 R_bl
Rbb_61_78 bitb_61_78 bitb_61_79 R_bl
Cb_61_78 bit_61_78 gnd C_bl
Cbb_61_78 bitb_61_78 gnd C_bl
Rb_61_79 bit_61_79 bit_61_80 R_bl
Rbb_61_79 bitb_61_79 bitb_61_80 R_bl
Cb_61_79 bit_61_79 gnd C_bl
Cbb_61_79 bitb_61_79 gnd C_bl
Rb_61_80 bit_61_80 bit_61_81 R_bl
Rbb_61_80 bitb_61_80 bitb_61_81 R_bl
Cb_61_80 bit_61_80 gnd C_bl
Cbb_61_80 bitb_61_80 gnd C_bl
Rb_61_81 bit_61_81 bit_61_82 R_bl
Rbb_61_81 bitb_61_81 bitb_61_82 R_bl
Cb_61_81 bit_61_81 gnd C_bl
Cbb_61_81 bitb_61_81 gnd C_bl
Rb_61_82 bit_61_82 bit_61_83 R_bl
Rbb_61_82 bitb_61_82 bitb_61_83 R_bl
Cb_61_82 bit_61_82 gnd C_bl
Cbb_61_82 bitb_61_82 gnd C_bl
Rb_61_83 bit_61_83 bit_61_84 R_bl
Rbb_61_83 bitb_61_83 bitb_61_84 R_bl
Cb_61_83 bit_61_83 gnd C_bl
Cbb_61_83 bitb_61_83 gnd C_bl
Rb_61_84 bit_61_84 bit_61_85 R_bl
Rbb_61_84 bitb_61_84 bitb_61_85 R_bl
Cb_61_84 bit_61_84 gnd C_bl
Cbb_61_84 bitb_61_84 gnd C_bl
Rb_61_85 bit_61_85 bit_61_86 R_bl
Rbb_61_85 bitb_61_85 bitb_61_86 R_bl
Cb_61_85 bit_61_85 gnd C_bl
Cbb_61_85 bitb_61_85 gnd C_bl
Rb_61_86 bit_61_86 bit_61_87 R_bl
Rbb_61_86 bitb_61_86 bitb_61_87 R_bl
Cb_61_86 bit_61_86 gnd C_bl
Cbb_61_86 bitb_61_86 gnd C_bl
Rb_61_87 bit_61_87 bit_61_88 R_bl
Rbb_61_87 bitb_61_87 bitb_61_88 R_bl
Cb_61_87 bit_61_87 gnd C_bl
Cbb_61_87 bitb_61_87 gnd C_bl
Rb_61_88 bit_61_88 bit_61_89 R_bl
Rbb_61_88 bitb_61_88 bitb_61_89 R_bl
Cb_61_88 bit_61_88 gnd C_bl
Cbb_61_88 bitb_61_88 gnd C_bl
Rb_61_89 bit_61_89 bit_61_90 R_bl
Rbb_61_89 bitb_61_89 bitb_61_90 R_bl
Cb_61_89 bit_61_89 gnd C_bl
Cbb_61_89 bitb_61_89 gnd C_bl
Rb_61_90 bit_61_90 bit_61_91 R_bl
Rbb_61_90 bitb_61_90 bitb_61_91 R_bl
Cb_61_90 bit_61_90 gnd C_bl
Cbb_61_90 bitb_61_90 gnd C_bl
Rb_61_91 bit_61_91 bit_61_92 R_bl
Rbb_61_91 bitb_61_91 bitb_61_92 R_bl
Cb_61_91 bit_61_91 gnd C_bl
Cbb_61_91 bitb_61_91 gnd C_bl
Rb_61_92 bit_61_92 bit_61_93 R_bl
Rbb_61_92 bitb_61_92 bitb_61_93 R_bl
Cb_61_92 bit_61_92 gnd C_bl
Cbb_61_92 bitb_61_92 gnd C_bl
Rb_61_93 bit_61_93 bit_61_94 R_bl
Rbb_61_93 bitb_61_93 bitb_61_94 R_bl
Cb_61_93 bit_61_93 gnd C_bl
Cbb_61_93 bitb_61_93 gnd C_bl
Rb_61_94 bit_61_94 bit_61_95 R_bl
Rbb_61_94 bitb_61_94 bitb_61_95 R_bl
Cb_61_94 bit_61_94 gnd C_bl
Cbb_61_94 bitb_61_94 gnd C_bl
Rb_61_95 bit_61_95 bit_61_96 R_bl
Rbb_61_95 bitb_61_95 bitb_61_96 R_bl
Cb_61_95 bit_61_95 gnd C_bl
Cbb_61_95 bitb_61_95 gnd C_bl
Rb_61_96 bit_61_96 bit_61_97 R_bl
Rbb_61_96 bitb_61_96 bitb_61_97 R_bl
Cb_61_96 bit_61_96 gnd C_bl
Cbb_61_96 bitb_61_96 gnd C_bl
Rb_61_97 bit_61_97 bit_61_98 R_bl
Rbb_61_97 bitb_61_97 bitb_61_98 R_bl
Cb_61_97 bit_61_97 gnd C_bl
Cbb_61_97 bitb_61_97 gnd C_bl
Rb_61_98 bit_61_98 bit_61_99 R_bl
Rbb_61_98 bitb_61_98 bitb_61_99 R_bl
Cb_61_98 bit_61_98 gnd C_bl
Cbb_61_98 bitb_61_98 gnd C_bl
Rb_61_99 bit_61_99 bit_61_100 R_bl
Rbb_61_99 bitb_61_99 bitb_61_100 R_bl
Cb_61_99 bit_61_99 gnd C_bl
Cbb_61_99 bitb_61_99 gnd C_bl
Rb_62_0 bit_62_0 bit_62_1 R_bl
Rbb_62_0 bitb_62_0 bitb_62_1 R_bl
Cb_62_0 bit_62_0 gnd C_bl
Cbb_62_0 bitb_62_0 gnd C_bl
Rb_62_1 bit_62_1 bit_62_2 R_bl
Rbb_62_1 bitb_62_1 bitb_62_2 R_bl
Cb_62_1 bit_62_1 gnd C_bl
Cbb_62_1 bitb_62_1 gnd C_bl
Rb_62_2 bit_62_2 bit_62_3 R_bl
Rbb_62_2 bitb_62_2 bitb_62_3 R_bl
Cb_62_2 bit_62_2 gnd C_bl
Cbb_62_2 bitb_62_2 gnd C_bl
Rb_62_3 bit_62_3 bit_62_4 R_bl
Rbb_62_3 bitb_62_3 bitb_62_4 R_bl
Cb_62_3 bit_62_3 gnd C_bl
Cbb_62_3 bitb_62_3 gnd C_bl
Rb_62_4 bit_62_4 bit_62_5 R_bl
Rbb_62_4 bitb_62_4 bitb_62_5 R_bl
Cb_62_4 bit_62_4 gnd C_bl
Cbb_62_4 bitb_62_4 gnd C_bl
Rb_62_5 bit_62_5 bit_62_6 R_bl
Rbb_62_5 bitb_62_5 bitb_62_6 R_bl
Cb_62_5 bit_62_5 gnd C_bl
Cbb_62_5 bitb_62_5 gnd C_bl
Rb_62_6 bit_62_6 bit_62_7 R_bl
Rbb_62_6 bitb_62_6 bitb_62_7 R_bl
Cb_62_6 bit_62_6 gnd C_bl
Cbb_62_6 bitb_62_6 gnd C_bl
Rb_62_7 bit_62_7 bit_62_8 R_bl
Rbb_62_7 bitb_62_7 bitb_62_8 R_bl
Cb_62_7 bit_62_7 gnd C_bl
Cbb_62_7 bitb_62_7 gnd C_bl
Rb_62_8 bit_62_8 bit_62_9 R_bl
Rbb_62_8 bitb_62_8 bitb_62_9 R_bl
Cb_62_8 bit_62_8 gnd C_bl
Cbb_62_8 bitb_62_8 gnd C_bl
Rb_62_9 bit_62_9 bit_62_10 R_bl
Rbb_62_9 bitb_62_9 bitb_62_10 R_bl
Cb_62_9 bit_62_9 gnd C_bl
Cbb_62_9 bitb_62_9 gnd C_bl
Rb_62_10 bit_62_10 bit_62_11 R_bl
Rbb_62_10 bitb_62_10 bitb_62_11 R_bl
Cb_62_10 bit_62_10 gnd C_bl
Cbb_62_10 bitb_62_10 gnd C_bl
Rb_62_11 bit_62_11 bit_62_12 R_bl
Rbb_62_11 bitb_62_11 bitb_62_12 R_bl
Cb_62_11 bit_62_11 gnd C_bl
Cbb_62_11 bitb_62_11 gnd C_bl
Rb_62_12 bit_62_12 bit_62_13 R_bl
Rbb_62_12 bitb_62_12 bitb_62_13 R_bl
Cb_62_12 bit_62_12 gnd C_bl
Cbb_62_12 bitb_62_12 gnd C_bl
Rb_62_13 bit_62_13 bit_62_14 R_bl
Rbb_62_13 bitb_62_13 bitb_62_14 R_bl
Cb_62_13 bit_62_13 gnd C_bl
Cbb_62_13 bitb_62_13 gnd C_bl
Rb_62_14 bit_62_14 bit_62_15 R_bl
Rbb_62_14 bitb_62_14 bitb_62_15 R_bl
Cb_62_14 bit_62_14 gnd C_bl
Cbb_62_14 bitb_62_14 gnd C_bl
Rb_62_15 bit_62_15 bit_62_16 R_bl
Rbb_62_15 bitb_62_15 bitb_62_16 R_bl
Cb_62_15 bit_62_15 gnd C_bl
Cbb_62_15 bitb_62_15 gnd C_bl
Rb_62_16 bit_62_16 bit_62_17 R_bl
Rbb_62_16 bitb_62_16 bitb_62_17 R_bl
Cb_62_16 bit_62_16 gnd C_bl
Cbb_62_16 bitb_62_16 gnd C_bl
Rb_62_17 bit_62_17 bit_62_18 R_bl
Rbb_62_17 bitb_62_17 bitb_62_18 R_bl
Cb_62_17 bit_62_17 gnd C_bl
Cbb_62_17 bitb_62_17 gnd C_bl
Rb_62_18 bit_62_18 bit_62_19 R_bl
Rbb_62_18 bitb_62_18 bitb_62_19 R_bl
Cb_62_18 bit_62_18 gnd C_bl
Cbb_62_18 bitb_62_18 gnd C_bl
Rb_62_19 bit_62_19 bit_62_20 R_bl
Rbb_62_19 bitb_62_19 bitb_62_20 R_bl
Cb_62_19 bit_62_19 gnd C_bl
Cbb_62_19 bitb_62_19 gnd C_bl
Rb_62_20 bit_62_20 bit_62_21 R_bl
Rbb_62_20 bitb_62_20 bitb_62_21 R_bl
Cb_62_20 bit_62_20 gnd C_bl
Cbb_62_20 bitb_62_20 gnd C_bl
Rb_62_21 bit_62_21 bit_62_22 R_bl
Rbb_62_21 bitb_62_21 bitb_62_22 R_bl
Cb_62_21 bit_62_21 gnd C_bl
Cbb_62_21 bitb_62_21 gnd C_bl
Rb_62_22 bit_62_22 bit_62_23 R_bl
Rbb_62_22 bitb_62_22 bitb_62_23 R_bl
Cb_62_22 bit_62_22 gnd C_bl
Cbb_62_22 bitb_62_22 gnd C_bl
Rb_62_23 bit_62_23 bit_62_24 R_bl
Rbb_62_23 bitb_62_23 bitb_62_24 R_bl
Cb_62_23 bit_62_23 gnd C_bl
Cbb_62_23 bitb_62_23 gnd C_bl
Rb_62_24 bit_62_24 bit_62_25 R_bl
Rbb_62_24 bitb_62_24 bitb_62_25 R_bl
Cb_62_24 bit_62_24 gnd C_bl
Cbb_62_24 bitb_62_24 gnd C_bl
Rb_62_25 bit_62_25 bit_62_26 R_bl
Rbb_62_25 bitb_62_25 bitb_62_26 R_bl
Cb_62_25 bit_62_25 gnd C_bl
Cbb_62_25 bitb_62_25 gnd C_bl
Rb_62_26 bit_62_26 bit_62_27 R_bl
Rbb_62_26 bitb_62_26 bitb_62_27 R_bl
Cb_62_26 bit_62_26 gnd C_bl
Cbb_62_26 bitb_62_26 gnd C_bl
Rb_62_27 bit_62_27 bit_62_28 R_bl
Rbb_62_27 bitb_62_27 bitb_62_28 R_bl
Cb_62_27 bit_62_27 gnd C_bl
Cbb_62_27 bitb_62_27 gnd C_bl
Rb_62_28 bit_62_28 bit_62_29 R_bl
Rbb_62_28 bitb_62_28 bitb_62_29 R_bl
Cb_62_28 bit_62_28 gnd C_bl
Cbb_62_28 bitb_62_28 gnd C_bl
Rb_62_29 bit_62_29 bit_62_30 R_bl
Rbb_62_29 bitb_62_29 bitb_62_30 R_bl
Cb_62_29 bit_62_29 gnd C_bl
Cbb_62_29 bitb_62_29 gnd C_bl
Rb_62_30 bit_62_30 bit_62_31 R_bl
Rbb_62_30 bitb_62_30 bitb_62_31 R_bl
Cb_62_30 bit_62_30 gnd C_bl
Cbb_62_30 bitb_62_30 gnd C_bl
Rb_62_31 bit_62_31 bit_62_32 R_bl
Rbb_62_31 bitb_62_31 bitb_62_32 R_bl
Cb_62_31 bit_62_31 gnd C_bl
Cbb_62_31 bitb_62_31 gnd C_bl
Rb_62_32 bit_62_32 bit_62_33 R_bl
Rbb_62_32 bitb_62_32 bitb_62_33 R_bl
Cb_62_32 bit_62_32 gnd C_bl
Cbb_62_32 bitb_62_32 gnd C_bl
Rb_62_33 bit_62_33 bit_62_34 R_bl
Rbb_62_33 bitb_62_33 bitb_62_34 R_bl
Cb_62_33 bit_62_33 gnd C_bl
Cbb_62_33 bitb_62_33 gnd C_bl
Rb_62_34 bit_62_34 bit_62_35 R_bl
Rbb_62_34 bitb_62_34 bitb_62_35 R_bl
Cb_62_34 bit_62_34 gnd C_bl
Cbb_62_34 bitb_62_34 gnd C_bl
Rb_62_35 bit_62_35 bit_62_36 R_bl
Rbb_62_35 bitb_62_35 bitb_62_36 R_bl
Cb_62_35 bit_62_35 gnd C_bl
Cbb_62_35 bitb_62_35 gnd C_bl
Rb_62_36 bit_62_36 bit_62_37 R_bl
Rbb_62_36 bitb_62_36 bitb_62_37 R_bl
Cb_62_36 bit_62_36 gnd C_bl
Cbb_62_36 bitb_62_36 gnd C_bl
Rb_62_37 bit_62_37 bit_62_38 R_bl
Rbb_62_37 bitb_62_37 bitb_62_38 R_bl
Cb_62_37 bit_62_37 gnd C_bl
Cbb_62_37 bitb_62_37 gnd C_bl
Rb_62_38 bit_62_38 bit_62_39 R_bl
Rbb_62_38 bitb_62_38 bitb_62_39 R_bl
Cb_62_38 bit_62_38 gnd C_bl
Cbb_62_38 bitb_62_38 gnd C_bl
Rb_62_39 bit_62_39 bit_62_40 R_bl
Rbb_62_39 bitb_62_39 bitb_62_40 R_bl
Cb_62_39 bit_62_39 gnd C_bl
Cbb_62_39 bitb_62_39 gnd C_bl
Rb_62_40 bit_62_40 bit_62_41 R_bl
Rbb_62_40 bitb_62_40 bitb_62_41 R_bl
Cb_62_40 bit_62_40 gnd C_bl
Cbb_62_40 bitb_62_40 gnd C_bl
Rb_62_41 bit_62_41 bit_62_42 R_bl
Rbb_62_41 bitb_62_41 bitb_62_42 R_bl
Cb_62_41 bit_62_41 gnd C_bl
Cbb_62_41 bitb_62_41 gnd C_bl
Rb_62_42 bit_62_42 bit_62_43 R_bl
Rbb_62_42 bitb_62_42 bitb_62_43 R_bl
Cb_62_42 bit_62_42 gnd C_bl
Cbb_62_42 bitb_62_42 gnd C_bl
Rb_62_43 bit_62_43 bit_62_44 R_bl
Rbb_62_43 bitb_62_43 bitb_62_44 R_bl
Cb_62_43 bit_62_43 gnd C_bl
Cbb_62_43 bitb_62_43 gnd C_bl
Rb_62_44 bit_62_44 bit_62_45 R_bl
Rbb_62_44 bitb_62_44 bitb_62_45 R_bl
Cb_62_44 bit_62_44 gnd C_bl
Cbb_62_44 bitb_62_44 gnd C_bl
Rb_62_45 bit_62_45 bit_62_46 R_bl
Rbb_62_45 bitb_62_45 bitb_62_46 R_bl
Cb_62_45 bit_62_45 gnd C_bl
Cbb_62_45 bitb_62_45 gnd C_bl
Rb_62_46 bit_62_46 bit_62_47 R_bl
Rbb_62_46 bitb_62_46 bitb_62_47 R_bl
Cb_62_46 bit_62_46 gnd C_bl
Cbb_62_46 bitb_62_46 gnd C_bl
Rb_62_47 bit_62_47 bit_62_48 R_bl
Rbb_62_47 bitb_62_47 bitb_62_48 R_bl
Cb_62_47 bit_62_47 gnd C_bl
Cbb_62_47 bitb_62_47 gnd C_bl
Rb_62_48 bit_62_48 bit_62_49 R_bl
Rbb_62_48 bitb_62_48 bitb_62_49 R_bl
Cb_62_48 bit_62_48 gnd C_bl
Cbb_62_48 bitb_62_48 gnd C_bl
Rb_62_49 bit_62_49 bit_62_50 R_bl
Rbb_62_49 bitb_62_49 bitb_62_50 R_bl
Cb_62_49 bit_62_49 gnd C_bl
Cbb_62_49 bitb_62_49 gnd C_bl
Rb_62_50 bit_62_50 bit_62_51 R_bl
Rbb_62_50 bitb_62_50 bitb_62_51 R_bl
Cb_62_50 bit_62_50 gnd C_bl
Cbb_62_50 bitb_62_50 gnd C_bl
Rb_62_51 bit_62_51 bit_62_52 R_bl
Rbb_62_51 bitb_62_51 bitb_62_52 R_bl
Cb_62_51 bit_62_51 gnd C_bl
Cbb_62_51 bitb_62_51 gnd C_bl
Rb_62_52 bit_62_52 bit_62_53 R_bl
Rbb_62_52 bitb_62_52 bitb_62_53 R_bl
Cb_62_52 bit_62_52 gnd C_bl
Cbb_62_52 bitb_62_52 gnd C_bl
Rb_62_53 bit_62_53 bit_62_54 R_bl
Rbb_62_53 bitb_62_53 bitb_62_54 R_bl
Cb_62_53 bit_62_53 gnd C_bl
Cbb_62_53 bitb_62_53 gnd C_bl
Rb_62_54 bit_62_54 bit_62_55 R_bl
Rbb_62_54 bitb_62_54 bitb_62_55 R_bl
Cb_62_54 bit_62_54 gnd C_bl
Cbb_62_54 bitb_62_54 gnd C_bl
Rb_62_55 bit_62_55 bit_62_56 R_bl
Rbb_62_55 bitb_62_55 bitb_62_56 R_bl
Cb_62_55 bit_62_55 gnd C_bl
Cbb_62_55 bitb_62_55 gnd C_bl
Rb_62_56 bit_62_56 bit_62_57 R_bl
Rbb_62_56 bitb_62_56 bitb_62_57 R_bl
Cb_62_56 bit_62_56 gnd C_bl
Cbb_62_56 bitb_62_56 gnd C_bl
Rb_62_57 bit_62_57 bit_62_58 R_bl
Rbb_62_57 bitb_62_57 bitb_62_58 R_bl
Cb_62_57 bit_62_57 gnd C_bl
Cbb_62_57 bitb_62_57 gnd C_bl
Rb_62_58 bit_62_58 bit_62_59 R_bl
Rbb_62_58 bitb_62_58 bitb_62_59 R_bl
Cb_62_58 bit_62_58 gnd C_bl
Cbb_62_58 bitb_62_58 gnd C_bl
Rb_62_59 bit_62_59 bit_62_60 R_bl
Rbb_62_59 bitb_62_59 bitb_62_60 R_bl
Cb_62_59 bit_62_59 gnd C_bl
Cbb_62_59 bitb_62_59 gnd C_bl
Rb_62_60 bit_62_60 bit_62_61 R_bl
Rbb_62_60 bitb_62_60 bitb_62_61 R_bl
Cb_62_60 bit_62_60 gnd C_bl
Cbb_62_60 bitb_62_60 gnd C_bl
Rb_62_61 bit_62_61 bit_62_62 R_bl
Rbb_62_61 bitb_62_61 bitb_62_62 R_bl
Cb_62_61 bit_62_61 gnd C_bl
Cbb_62_61 bitb_62_61 gnd C_bl
Rb_62_62 bit_62_62 bit_62_63 R_bl
Rbb_62_62 bitb_62_62 bitb_62_63 R_bl
Cb_62_62 bit_62_62 gnd C_bl
Cbb_62_62 bitb_62_62 gnd C_bl
Rb_62_63 bit_62_63 bit_62_64 R_bl
Rbb_62_63 bitb_62_63 bitb_62_64 R_bl
Cb_62_63 bit_62_63 gnd C_bl
Cbb_62_63 bitb_62_63 gnd C_bl
Rb_62_64 bit_62_64 bit_62_65 R_bl
Rbb_62_64 bitb_62_64 bitb_62_65 R_bl
Cb_62_64 bit_62_64 gnd C_bl
Cbb_62_64 bitb_62_64 gnd C_bl
Rb_62_65 bit_62_65 bit_62_66 R_bl
Rbb_62_65 bitb_62_65 bitb_62_66 R_bl
Cb_62_65 bit_62_65 gnd C_bl
Cbb_62_65 bitb_62_65 gnd C_bl
Rb_62_66 bit_62_66 bit_62_67 R_bl
Rbb_62_66 bitb_62_66 bitb_62_67 R_bl
Cb_62_66 bit_62_66 gnd C_bl
Cbb_62_66 bitb_62_66 gnd C_bl
Rb_62_67 bit_62_67 bit_62_68 R_bl
Rbb_62_67 bitb_62_67 bitb_62_68 R_bl
Cb_62_67 bit_62_67 gnd C_bl
Cbb_62_67 bitb_62_67 gnd C_bl
Rb_62_68 bit_62_68 bit_62_69 R_bl
Rbb_62_68 bitb_62_68 bitb_62_69 R_bl
Cb_62_68 bit_62_68 gnd C_bl
Cbb_62_68 bitb_62_68 gnd C_bl
Rb_62_69 bit_62_69 bit_62_70 R_bl
Rbb_62_69 bitb_62_69 bitb_62_70 R_bl
Cb_62_69 bit_62_69 gnd C_bl
Cbb_62_69 bitb_62_69 gnd C_bl
Rb_62_70 bit_62_70 bit_62_71 R_bl
Rbb_62_70 bitb_62_70 bitb_62_71 R_bl
Cb_62_70 bit_62_70 gnd C_bl
Cbb_62_70 bitb_62_70 gnd C_bl
Rb_62_71 bit_62_71 bit_62_72 R_bl
Rbb_62_71 bitb_62_71 bitb_62_72 R_bl
Cb_62_71 bit_62_71 gnd C_bl
Cbb_62_71 bitb_62_71 gnd C_bl
Rb_62_72 bit_62_72 bit_62_73 R_bl
Rbb_62_72 bitb_62_72 bitb_62_73 R_bl
Cb_62_72 bit_62_72 gnd C_bl
Cbb_62_72 bitb_62_72 gnd C_bl
Rb_62_73 bit_62_73 bit_62_74 R_bl
Rbb_62_73 bitb_62_73 bitb_62_74 R_bl
Cb_62_73 bit_62_73 gnd C_bl
Cbb_62_73 bitb_62_73 gnd C_bl
Rb_62_74 bit_62_74 bit_62_75 R_bl
Rbb_62_74 bitb_62_74 bitb_62_75 R_bl
Cb_62_74 bit_62_74 gnd C_bl
Cbb_62_74 bitb_62_74 gnd C_bl
Rb_62_75 bit_62_75 bit_62_76 R_bl
Rbb_62_75 bitb_62_75 bitb_62_76 R_bl
Cb_62_75 bit_62_75 gnd C_bl
Cbb_62_75 bitb_62_75 gnd C_bl
Rb_62_76 bit_62_76 bit_62_77 R_bl
Rbb_62_76 bitb_62_76 bitb_62_77 R_bl
Cb_62_76 bit_62_76 gnd C_bl
Cbb_62_76 bitb_62_76 gnd C_bl
Rb_62_77 bit_62_77 bit_62_78 R_bl
Rbb_62_77 bitb_62_77 bitb_62_78 R_bl
Cb_62_77 bit_62_77 gnd C_bl
Cbb_62_77 bitb_62_77 gnd C_bl
Rb_62_78 bit_62_78 bit_62_79 R_bl
Rbb_62_78 bitb_62_78 bitb_62_79 R_bl
Cb_62_78 bit_62_78 gnd C_bl
Cbb_62_78 bitb_62_78 gnd C_bl
Rb_62_79 bit_62_79 bit_62_80 R_bl
Rbb_62_79 bitb_62_79 bitb_62_80 R_bl
Cb_62_79 bit_62_79 gnd C_bl
Cbb_62_79 bitb_62_79 gnd C_bl
Rb_62_80 bit_62_80 bit_62_81 R_bl
Rbb_62_80 bitb_62_80 bitb_62_81 R_bl
Cb_62_80 bit_62_80 gnd C_bl
Cbb_62_80 bitb_62_80 gnd C_bl
Rb_62_81 bit_62_81 bit_62_82 R_bl
Rbb_62_81 bitb_62_81 bitb_62_82 R_bl
Cb_62_81 bit_62_81 gnd C_bl
Cbb_62_81 bitb_62_81 gnd C_bl
Rb_62_82 bit_62_82 bit_62_83 R_bl
Rbb_62_82 bitb_62_82 bitb_62_83 R_bl
Cb_62_82 bit_62_82 gnd C_bl
Cbb_62_82 bitb_62_82 gnd C_bl
Rb_62_83 bit_62_83 bit_62_84 R_bl
Rbb_62_83 bitb_62_83 bitb_62_84 R_bl
Cb_62_83 bit_62_83 gnd C_bl
Cbb_62_83 bitb_62_83 gnd C_bl
Rb_62_84 bit_62_84 bit_62_85 R_bl
Rbb_62_84 bitb_62_84 bitb_62_85 R_bl
Cb_62_84 bit_62_84 gnd C_bl
Cbb_62_84 bitb_62_84 gnd C_bl
Rb_62_85 bit_62_85 bit_62_86 R_bl
Rbb_62_85 bitb_62_85 bitb_62_86 R_bl
Cb_62_85 bit_62_85 gnd C_bl
Cbb_62_85 bitb_62_85 gnd C_bl
Rb_62_86 bit_62_86 bit_62_87 R_bl
Rbb_62_86 bitb_62_86 bitb_62_87 R_bl
Cb_62_86 bit_62_86 gnd C_bl
Cbb_62_86 bitb_62_86 gnd C_bl
Rb_62_87 bit_62_87 bit_62_88 R_bl
Rbb_62_87 bitb_62_87 bitb_62_88 R_bl
Cb_62_87 bit_62_87 gnd C_bl
Cbb_62_87 bitb_62_87 gnd C_bl
Rb_62_88 bit_62_88 bit_62_89 R_bl
Rbb_62_88 bitb_62_88 bitb_62_89 R_bl
Cb_62_88 bit_62_88 gnd C_bl
Cbb_62_88 bitb_62_88 gnd C_bl
Rb_62_89 bit_62_89 bit_62_90 R_bl
Rbb_62_89 bitb_62_89 bitb_62_90 R_bl
Cb_62_89 bit_62_89 gnd C_bl
Cbb_62_89 bitb_62_89 gnd C_bl
Rb_62_90 bit_62_90 bit_62_91 R_bl
Rbb_62_90 bitb_62_90 bitb_62_91 R_bl
Cb_62_90 bit_62_90 gnd C_bl
Cbb_62_90 bitb_62_90 gnd C_bl
Rb_62_91 bit_62_91 bit_62_92 R_bl
Rbb_62_91 bitb_62_91 bitb_62_92 R_bl
Cb_62_91 bit_62_91 gnd C_bl
Cbb_62_91 bitb_62_91 gnd C_bl
Rb_62_92 bit_62_92 bit_62_93 R_bl
Rbb_62_92 bitb_62_92 bitb_62_93 R_bl
Cb_62_92 bit_62_92 gnd C_bl
Cbb_62_92 bitb_62_92 gnd C_bl
Rb_62_93 bit_62_93 bit_62_94 R_bl
Rbb_62_93 bitb_62_93 bitb_62_94 R_bl
Cb_62_93 bit_62_93 gnd C_bl
Cbb_62_93 bitb_62_93 gnd C_bl
Rb_62_94 bit_62_94 bit_62_95 R_bl
Rbb_62_94 bitb_62_94 bitb_62_95 R_bl
Cb_62_94 bit_62_94 gnd C_bl
Cbb_62_94 bitb_62_94 gnd C_bl
Rb_62_95 bit_62_95 bit_62_96 R_bl
Rbb_62_95 bitb_62_95 bitb_62_96 R_bl
Cb_62_95 bit_62_95 gnd C_bl
Cbb_62_95 bitb_62_95 gnd C_bl
Rb_62_96 bit_62_96 bit_62_97 R_bl
Rbb_62_96 bitb_62_96 bitb_62_97 R_bl
Cb_62_96 bit_62_96 gnd C_bl
Cbb_62_96 bitb_62_96 gnd C_bl
Rb_62_97 bit_62_97 bit_62_98 R_bl
Rbb_62_97 bitb_62_97 bitb_62_98 R_bl
Cb_62_97 bit_62_97 gnd C_bl
Cbb_62_97 bitb_62_97 gnd C_bl
Rb_62_98 bit_62_98 bit_62_99 R_bl
Rbb_62_98 bitb_62_98 bitb_62_99 R_bl
Cb_62_98 bit_62_98 gnd C_bl
Cbb_62_98 bitb_62_98 gnd C_bl
Rb_62_99 bit_62_99 bit_62_100 R_bl
Rbb_62_99 bitb_62_99 bitb_62_100 R_bl
Cb_62_99 bit_62_99 gnd C_bl
Cbb_62_99 bitb_62_99 gnd C_bl
Rb_63_0 bit_63_0 bit_63_1 R_bl
Rbb_63_0 bitb_63_0 bitb_63_1 R_bl
Cb_63_0 bit_63_0 gnd C_bl
Cbb_63_0 bitb_63_0 gnd C_bl
Rb_63_1 bit_63_1 bit_63_2 R_bl
Rbb_63_1 bitb_63_1 bitb_63_2 R_bl
Cb_63_1 bit_63_1 gnd C_bl
Cbb_63_1 bitb_63_1 gnd C_bl
Rb_63_2 bit_63_2 bit_63_3 R_bl
Rbb_63_2 bitb_63_2 bitb_63_3 R_bl
Cb_63_2 bit_63_2 gnd C_bl
Cbb_63_2 bitb_63_2 gnd C_bl
Rb_63_3 bit_63_3 bit_63_4 R_bl
Rbb_63_3 bitb_63_3 bitb_63_4 R_bl
Cb_63_3 bit_63_3 gnd C_bl
Cbb_63_3 bitb_63_3 gnd C_bl
Rb_63_4 bit_63_4 bit_63_5 R_bl
Rbb_63_4 bitb_63_4 bitb_63_5 R_bl
Cb_63_4 bit_63_4 gnd C_bl
Cbb_63_4 bitb_63_4 gnd C_bl
Rb_63_5 bit_63_5 bit_63_6 R_bl
Rbb_63_5 bitb_63_5 bitb_63_6 R_bl
Cb_63_5 bit_63_5 gnd C_bl
Cbb_63_5 bitb_63_5 gnd C_bl
Rb_63_6 bit_63_6 bit_63_7 R_bl
Rbb_63_6 bitb_63_6 bitb_63_7 R_bl
Cb_63_6 bit_63_6 gnd C_bl
Cbb_63_6 bitb_63_6 gnd C_bl
Rb_63_7 bit_63_7 bit_63_8 R_bl
Rbb_63_7 bitb_63_7 bitb_63_8 R_bl
Cb_63_7 bit_63_7 gnd C_bl
Cbb_63_7 bitb_63_7 gnd C_bl
Rb_63_8 bit_63_8 bit_63_9 R_bl
Rbb_63_8 bitb_63_8 bitb_63_9 R_bl
Cb_63_8 bit_63_8 gnd C_bl
Cbb_63_8 bitb_63_8 gnd C_bl
Rb_63_9 bit_63_9 bit_63_10 R_bl
Rbb_63_9 bitb_63_9 bitb_63_10 R_bl
Cb_63_9 bit_63_9 gnd C_bl
Cbb_63_9 bitb_63_9 gnd C_bl
Rb_63_10 bit_63_10 bit_63_11 R_bl
Rbb_63_10 bitb_63_10 bitb_63_11 R_bl
Cb_63_10 bit_63_10 gnd C_bl
Cbb_63_10 bitb_63_10 gnd C_bl
Rb_63_11 bit_63_11 bit_63_12 R_bl
Rbb_63_11 bitb_63_11 bitb_63_12 R_bl
Cb_63_11 bit_63_11 gnd C_bl
Cbb_63_11 bitb_63_11 gnd C_bl
Rb_63_12 bit_63_12 bit_63_13 R_bl
Rbb_63_12 bitb_63_12 bitb_63_13 R_bl
Cb_63_12 bit_63_12 gnd C_bl
Cbb_63_12 bitb_63_12 gnd C_bl
Rb_63_13 bit_63_13 bit_63_14 R_bl
Rbb_63_13 bitb_63_13 bitb_63_14 R_bl
Cb_63_13 bit_63_13 gnd C_bl
Cbb_63_13 bitb_63_13 gnd C_bl
Rb_63_14 bit_63_14 bit_63_15 R_bl
Rbb_63_14 bitb_63_14 bitb_63_15 R_bl
Cb_63_14 bit_63_14 gnd C_bl
Cbb_63_14 bitb_63_14 gnd C_bl
Rb_63_15 bit_63_15 bit_63_16 R_bl
Rbb_63_15 bitb_63_15 bitb_63_16 R_bl
Cb_63_15 bit_63_15 gnd C_bl
Cbb_63_15 bitb_63_15 gnd C_bl
Rb_63_16 bit_63_16 bit_63_17 R_bl
Rbb_63_16 bitb_63_16 bitb_63_17 R_bl
Cb_63_16 bit_63_16 gnd C_bl
Cbb_63_16 bitb_63_16 gnd C_bl
Rb_63_17 bit_63_17 bit_63_18 R_bl
Rbb_63_17 bitb_63_17 bitb_63_18 R_bl
Cb_63_17 bit_63_17 gnd C_bl
Cbb_63_17 bitb_63_17 gnd C_bl
Rb_63_18 bit_63_18 bit_63_19 R_bl
Rbb_63_18 bitb_63_18 bitb_63_19 R_bl
Cb_63_18 bit_63_18 gnd C_bl
Cbb_63_18 bitb_63_18 gnd C_bl
Rb_63_19 bit_63_19 bit_63_20 R_bl
Rbb_63_19 bitb_63_19 bitb_63_20 R_bl
Cb_63_19 bit_63_19 gnd C_bl
Cbb_63_19 bitb_63_19 gnd C_bl
Rb_63_20 bit_63_20 bit_63_21 R_bl
Rbb_63_20 bitb_63_20 bitb_63_21 R_bl
Cb_63_20 bit_63_20 gnd C_bl
Cbb_63_20 bitb_63_20 gnd C_bl
Rb_63_21 bit_63_21 bit_63_22 R_bl
Rbb_63_21 bitb_63_21 bitb_63_22 R_bl
Cb_63_21 bit_63_21 gnd C_bl
Cbb_63_21 bitb_63_21 gnd C_bl
Rb_63_22 bit_63_22 bit_63_23 R_bl
Rbb_63_22 bitb_63_22 bitb_63_23 R_bl
Cb_63_22 bit_63_22 gnd C_bl
Cbb_63_22 bitb_63_22 gnd C_bl
Rb_63_23 bit_63_23 bit_63_24 R_bl
Rbb_63_23 bitb_63_23 bitb_63_24 R_bl
Cb_63_23 bit_63_23 gnd C_bl
Cbb_63_23 bitb_63_23 gnd C_bl
Rb_63_24 bit_63_24 bit_63_25 R_bl
Rbb_63_24 bitb_63_24 bitb_63_25 R_bl
Cb_63_24 bit_63_24 gnd C_bl
Cbb_63_24 bitb_63_24 gnd C_bl
Rb_63_25 bit_63_25 bit_63_26 R_bl
Rbb_63_25 bitb_63_25 bitb_63_26 R_bl
Cb_63_25 bit_63_25 gnd C_bl
Cbb_63_25 bitb_63_25 gnd C_bl
Rb_63_26 bit_63_26 bit_63_27 R_bl
Rbb_63_26 bitb_63_26 bitb_63_27 R_bl
Cb_63_26 bit_63_26 gnd C_bl
Cbb_63_26 bitb_63_26 gnd C_bl
Rb_63_27 bit_63_27 bit_63_28 R_bl
Rbb_63_27 bitb_63_27 bitb_63_28 R_bl
Cb_63_27 bit_63_27 gnd C_bl
Cbb_63_27 bitb_63_27 gnd C_bl
Rb_63_28 bit_63_28 bit_63_29 R_bl
Rbb_63_28 bitb_63_28 bitb_63_29 R_bl
Cb_63_28 bit_63_28 gnd C_bl
Cbb_63_28 bitb_63_28 gnd C_bl
Rb_63_29 bit_63_29 bit_63_30 R_bl
Rbb_63_29 bitb_63_29 bitb_63_30 R_bl
Cb_63_29 bit_63_29 gnd C_bl
Cbb_63_29 bitb_63_29 gnd C_bl
Rb_63_30 bit_63_30 bit_63_31 R_bl
Rbb_63_30 bitb_63_30 bitb_63_31 R_bl
Cb_63_30 bit_63_30 gnd C_bl
Cbb_63_30 bitb_63_30 gnd C_bl
Rb_63_31 bit_63_31 bit_63_32 R_bl
Rbb_63_31 bitb_63_31 bitb_63_32 R_bl
Cb_63_31 bit_63_31 gnd C_bl
Cbb_63_31 bitb_63_31 gnd C_bl
Rb_63_32 bit_63_32 bit_63_33 R_bl
Rbb_63_32 bitb_63_32 bitb_63_33 R_bl
Cb_63_32 bit_63_32 gnd C_bl
Cbb_63_32 bitb_63_32 gnd C_bl
Rb_63_33 bit_63_33 bit_63_34 R_bl
Rbb_63_33 bitb_63_33 bitb_63_34 R_bl
Cb_63_33 bit_63_33 gnd C_bl
Cbb_63_33 bitb_63_33 gnd C_bl
Rb_63_34 bit_63_34 bit_63_35 R_bl
Rbb_63_34 bitb_63_34 bitb_63_35 R_bl
Cb_63_34 bit_63_34 gnd C_bl
Cbb_63_34 bitb_63_34 gnd C_bl
Rb_63_35 bit_63_35 bit_63_36 R_bl
Rbb_63_35 bitb_63_35 bitb_63_36 R_bl
Cb_63_35 bit_63_35 gnd C_bl
Cbb_63_35 bitb_63_35 gnd C_bl
Rb_63_36 bit_63_36 bit_63_37 R_bl
Rbb_63_36 bitb_63_36 bitb_63_37 R_bl
Cb_63_36 bit_63_36 gnd C_bl
Cbb_63_36 bitb_63_36 gnd C_bl
Rb_63_37 bit_63_37 bit_63_38 R_bl
Rbb_63_37 bitb_63_37 bitb_63_38 R_bl
Cb_63_37 bit_63_37 gnd C_bl
Cbb_63_37 bitb_63_37 gnd C_bl
Rb_63_38 bit_63_38 bit_63_39 R_bl
Rbb_63_38 bitb_63_38 bitb_63_39 R_bl
Cb_63_38 bit_63_38 gnd C_bl
Cbb_63_38 bitb_63_38 gnd C_bl
Rb_63_39 bit_63_39 bit_63_40 R_bl
Rbb_63_39 bitb_63_39 bitb_63_40 R_bl
Cb_63_39 bit_63_39 gnd C_bl
Cbb_63_39 bitb_63_39 gnd C_bl
Rb_63_40 bit_63_40 bit_63_41 R_bl
Rbb_63_40 bitb_63_40 bitb_63_41 R_bl
Cb_63_40 bit_63_40 gnd C_bl
Cbb_63_40 bitb_63_40 gnd C_bl
Rb_63_41 bit_63_41 bit_63_42 R_bl
Rbb_63_41 bitb_63_41 bitb_63_42 R_bl
Cb_63_41 bit_63_41 gnd C_bl
Cbb_63_41 bitb_63_41 gnd C_bl
Rb_63_42 bit_63_42 bit_63_43 R_bl
Rbb_63_42 bitb_63_42 bitb_63_43 R_bl
Cb_63_42 bit_63_42 gnd C_bl
Cbb_63_42 bitb_63_42 gnd C_bl
Rb_63_43 bit_63_43 bit_63_44 R_bl
Rbb_63_43 bitb_63_43 bitb_63_44 R_bl
Cb_63_43 bit_63_43 gnd C_bl
Cbb_63_43 bitb_63_43 gnd C_bl
Rb_63_44 bit_63_44 bit_63_45 R_bl
Rbb_63_44 bitb_63_44 bitb_63_45 R_bl
Cb_63_44 bit_63_44 gnd C_bl
Cbb_63_44 bitb_63_44 gnd C_bl
Rb_63_45 bit_63_45 bit_63_46 R_bl
Rbb_63_45 bitb_63_45 bitb_63_46 R_bl
Cb_63_45 bit_63_45 gnd C_bl
Cbb_63_45 bitb_63_45 gnd C_bl
Rb_63_46 bit_63_46 bit_63_47 R_bl
Rbb_63_46 bitb_63_46 bitb_63_47 R_bl
Cb_63_46 bit_63_46 gnd C_bl
Cbb_63_46 bitb_63_46 gnd C_bl
Rb_63_47 bit_63_47 bit_63_48 R_bl
Rbb_63_47 bitb_63_47 bitb_63_48 R_bl
Cb_63_47 bit_63_47 gnd C_bl
Cbb_63_47 bitb_63_47 gnd C_bl
Rb_63_48 bit_63_48 bit_63_49 R_bl
Rbb_63_48 bitb_63_48 bitb_63_49 R_bl
Cb_63_48 bit_63_48 gnd C_bl
Cbb_63_48 bitb_63_48 gnd C_bl
Rb_63_49 bit_63_49 bit_63_50 R_bl
Rbb_63_49 bitb_63_49 bitb_63_50 R_bl
Cb_63_49 bit_63_49 gnd C_bl
Cbb_63_49 bitb_63_49 gnd C_bl
Rb_63_50 bit_63_50 bit_63_51 R_bl
Rbb_63_50 bitb_63_50 bitb_63_51 R_bl
Cb_63_50 bit_63_50 gnd C_bl
Cbb_63_50 bitb_63_50 gnd C_bl
Rb_63_51 bit_63_51 bit_63_52 R_bl
Rbb_63_51 bitb_63_51 bitb_63_52 R_bl
Cb_63_51 bit_63_51 gnd C_bl
Cbb_63_51 bitb_63_51 gnd C_bl
Rb_63_52 bit_63_52 bit_63_53 R_bl
Rbb_63_52 bitb_63_52 bitb_63_53 R_bl
Cb_63_52 bit_63_52 gnd C_bl
Cbb_63_52 bitb_63_52 gnd C_bl
Rb_63_53 bit_63_53 bit_63_54 R_bl
Rbb_63_53 bitb_63_53 bitb_63_54 R_bl
Cb_63_53 bit_63_53 gnd C_bl
Cbb_63_53 bitb_63_53 gnd C_bl
Rb_63_54 bit_63_54 bit_63_55 R_bl
Rbb_63_54 bitb_63_54 bitb_63_55 R_bl
Cb_63_54 bit_63_54 gnd C_bl
Cbb_63_54 bitb_63_54 gnd C_bl
Rb_63_55 bit_63_55 bit_63_56 R_bl
Rbb_63_55 bitb_63_55 bitb_63_56 R_bl
Cb_63_55 bit_63_55 gnd C_bl
Cbb_63_55 bitb_63_55 gnd C_bl
Rb_63_56 bit_63_56 bit_63_57 R_bl
Rbb_63_56 bitb_63_56 bitb_63_57 R_bl
Cb_63_56 bit_63_56 gnd C_bl
Cbb_63_56 bitb_63_56 gnd C_bl
Rb_63_57 bit_63_57 bit_63_58 R_bl
Rbb_63_57 bitb_63_57 bitb_63_58 R_bl
Cb_63_57 bit_63_57 gnd C_bl
Cbb_63_57 bitb_63_57 gnd C_bl
Rb_63_58 bit_63_58 bit_63_59 R_bl
Rbb_63_58 bitb_63_58 bitb_63_59 R_bl
Cb_63_58 bit_63_58 gnd C_bl
Cbb_63_58 bitb_63_58 gnd C_bl
Rb_63_59 bit_63_59 bit_63_60 R_bl
Rbb_63_59 bitb_63_59 bitb_63_60 R_bl
Cb_63_59 bit_63_59 gnd C_bl
Cbb_63_59 bitb_63_59 gnd C_bl
Rb_63_60 bit_63_60 bit_63_61 R_bl
Rbb_63_60 bitb_63_60 bitb_63_61 R_bl
Cb_63_60 bit_63_60 gnd C_bl
Cbb_63_60 bitb_63_60 gnd C_bl
Rb_63_61 bit_63_61 bit_63_62 R_bl
Rbb_63_61 bitb_63_61 bitb_63_62 R_bl
Cb_63_61 bit_63_61 gnd C_bl
Cbb_63_61 bitb_63_61 gnd C_bl
Rb_63_62 bit_63_62 bit_63_63 R_bl
Rbb_63_62 bitb_63_62 bitb_63_63 R_bl
Cb_63_62 bit_63_62 gnd C_bl
Cbb_63_62 bitb_63_62 gnd C_bl
Rb_63_63 bit_63_63 bit_63_64 R_bl
Rbb_63_63 bitb_63_63 bitb_63_64 R_bl
Cb_63_63 bit_63_63 gnd C_bl
Cbb_63_63 bitb_63_63 gnd C_bl
Rb_63_64 bit_63_64 bit_63_65 R_bl
Rbb_63_64 bitb_63_64 bitb_63_65 R_bl
Cb_63_64 bit_63_64 gnd C_bl
Cbb_63_64 bitb_63_64 gnd C_bl
Rb_63_65 bit_63_65 bit_63_66 R_bl
Rbb_63_65 bitb_63_65 bitb_63_66 R_bl
Cb_63_65 bit_63_65 gnd C_bl
Cbb_63_65 bitb_63_65 gnd C_bl
Rb_63_66 bit_63_66 bit_63_67 R_bl
Rbb_63_66 bitb_63_66 bitb_63_67 R_bl
Cb_63_66 bit_63_66 gnd C_bl
Cbb_63_66 bitb_63_66 gnd C_bl
Rb_63_67 bit_63_67 bit_63_68 R_bl
Rbb_63_67 bitb_63_67 bitb_63_68 R_bl
Cb_63_67 bit_63_67 gnd C_bl
Cbb_63_67 bitb_63_67 gnd C_bl
Rb_63_68 bit_63_68 bit_63_69 R_bl
Rbb_63_68 bitb_63_68 bitb_63_69 R_bl
Cb_63_68 bit_63_68 gnd C_bl
Cbb_63_68 bitb_63_68 gnd C_bl
Rb_63_69 bit_63_69 bit_63_70 R_bl
Rbb_63_69 bitb_63_69 bitb_63_70 R_bl
Cb_63_69 bit_63_69 gnd C_bl
Cbb_63_69 bitb_63_69 gnd C_bl
Rb_63_70 bit_63_70 bit_63_71 R_bl
Rbb_63_70 bitb_63_70 bitb_63_71 R_bl
Cb_63_70 bit_63_70 gnd C_bl
Cbb_63_70 bitb_63_70 gnd C_bl
Rb_63_71 bit_63_71 bit_63_72 R_bl
Rbb_63_71 bitb_63_71 bitb_63_72 R_bl
Cb_63_71 bit_63_71 gnd C_bl
Cbb_63_71 bitb_63_71 gnd C_bl
Rb_63_72 bit_63_72 bit_63_73 R_bl
Rbb_63_72 bitb_63_72 bitb_63_73 R_bl
Cb_63_72 bit_63_72 gnd C_bl
Cbb_63_72 bitb_63_72 gnd C_bl
Rb_63_73 bit_63_73 bit_63_74 R_bl
Rbb_63_73 bitb_63_73 bitb_63_74 R_bl
Cb_63_73 bit_63_73 gnd C_bl
Cbb_63_73 bitb_63_73 gnd C_bl
Rb_63_74 bit_63_74 bit_63_75 R_bl
Rbb_63_74 bitb_63_74 bitb_63_75 R_bl
Cb_63_74 bit_63_74 gnd C_bl
Cbb_63_74 bitb_63_74 gnd C_bl
Rb_63_75 bit_63_75 bit_63_76 R_bl
Rbb_63_75 bitb_63_75 bitb_63_76 R_bl
Cb_63_75 bit_63_75 gnd C_bl
Cbb_63_75 bitb_63_75 gnd C_bl
Rb_63_76 bit_63_76 bit_63_77 R_bl
Rbb_63_76 bitb_63_76 bitb_63_77 R_bl
Cb_63_76 bit_63_76 gnd C_bl
Cbb_63_76 bitb_63_76 gnd C_bl
Rb_63_77 bit_63_77 bit_63_78 R_bl
Rbb_63_77 bitb_63_77 bitb_63_78 R_bl
Cb_63_77 bit_63_77 gnd C_bl
Cbb_63_77 bitb_63_77 gnd C_bl
Rb_63_78 bit_63_78 bit_63_79 R_bl
Rbb_63_78 bitb_63_78 bitb_63_79 R_bl
Cb_63_78 bit_63_78 gnd C_bl
Cbb_63_78 bitb_63_78 gnd C_bl
Rb_63_79 bit_63_79 bit_63_80 R_bl
Rbb_63_79 bitb_63_79 bitb_63_80 R_bl
Cb_63_79 bit_63_79 gnd C_bl
Cbb_63_79 bitb_63_79 gnd C_bl
Rb_63_80 bit_63_80 bit_63_81 R_bl
Rbb_63_80 bitb_63_80 bitb_63_81 R_bl
Cb_63_80 bit_63_80 gnd C_bl
Cbb_63_80 bitb_63_80 gnd C_bl
Rb_63_81 bit_63_81 bit_63_82 R_bl
Rbb_63_81 bitb_63_81 bitb_63_82 R_bl
Cb_63_81 bit_63_81 gnd C_bl
Cbb_63_81 bitb_63_81 gnd C_bl
Rb_63_82 bit_63_82 bit_63_83 R_bl
Rbb_63_82 bitb_63_82 bitb_63_83 R_bl
Cb_63_82 bit_63_82 gnd C_bl
Cbb_63_82 bitb_63_82 gnd C_bl
Rb_63_83 bit_63_83 bit_63_84 R_bl
Rbb_63_83 bitb_63_83 bitb_63_84 R_bl
Cb_63_83 bit_63_83 gnd C_bl
Cbb_63_83 bitb_63_83 gnd C_bl
Rb_63_84 bit_63_84 bit_63_85 R_bl
Rbb_63_84 bitb_63_84 bitb_63_85 R_bl
Cb_63_84 bit_63_84 gnd C_bl
Cbb_63_84 bitb_63_84 gnd C_bl
Rb_63_85 bit_63_85 bit_63_86 R_bl
Rbb_63_85 bitb_63_85 bitb_63_86 R_bl
Cb_63_85 bit_63_85 gnd C_bl
Cbb_63_85 bitb_63_85 gnd C_bl
Rb_63_86 bit_63_86 bit_63_87 R_bl
Rbb_63_86 bitb_63_86 bitb_63_87 R_bl
Cb_63_86 bit_63_86 gnd C_bl
Cbb_63_86 bitb_63_86 gnd C_bl
Rb_63_87 bit_63_87 bit_63_88 R_bl
Rbb_63_87 bitb_63_87 bitb_63_88 R_bl
Cb_63_87 bit_63_87 gnd C_bl
Cbb_63_87 bitb_63_87 gnd C_bl
Rb_63_88 bit_63_88 bit_63_89 R_bl
Rbb_63_88 bitb_63_88 bitb_63_89 R_bl
Cb_63_88 bit_63_88 gnd C_bl
Cbb_63_88 bitb_63_88 gnd C_bl
Rb_63_89 bit_63_89 bit_63_90 R_bl
Rbb_63_89 bitb_63_89 bitb_63_90 R_bl
Cb_63_89 bit_63_89 gnd C_bl
Cbb_63_89 bitb_63_89 gnd C_bl
Rb_63_90 bit_63_90 bit_63_91 R_bl
Rbb_63_90 bitb_63_90 bitb_63_91 R_bl
Cb_63_90 bit_63_90 gnd C_bl
Cbb_63_90 bitb_63_90 gnd C_bl
Rb_63_91 bit_63_91 bit_63_92 R_bl
Rbb_63_91 bitb_63_91 bitb_63_92 R_bl
Cb_63_91 bit_63_91 gnd C_bl
Cbb_63_91 bitb_63_91 gnd C_bl
Rb_63_92 bit_63_92 bit_63_93 R_bl
Rbb_63_92 bitb_63_92 bitb_63_93 R_bl
Cb_63_92 bit_63_92 gnd C_bl
Cbb_63_92 bitb_63_92 gnd C_bl
Rb_63_93 bit_63_93 bit_63_94 R_bl
Rbb_63_93 bitb_63_93 bitb_63_94 R_bl
Cb_63_93 bit_63_93 gnd C_bl
Cbb_63_93 bitb_63_93 gnd C_bl
Rb_63_94 bit_63_94 bit_63_95 R_bl
Rbb_63_94 bitb_63_94 bitb_63_95 R_bl
Cb_63_94 bit_63_94 gnd C_bl
Cbb_63_94 bitb_63_94 gnd C_bl
Rb_63_95 bit_63_95 bit_63_96 R_bl
Rbb_63_95 bitb_63_95 bitb_63_96 R_bl
Cb_63_95 bit_63_95 gnd C_bl
Cbb_63_95 bitb_63_95 gnd C_bl
Rb_63_96 bit_63_96 bit_63_97 R_bl
Rbb_63_96 bitb_63_96 bitb_63_97 R_bl
Cb_63_96 bit_63_96 gnd C_bl
Cbb_63_96 bitb_63_96 gnd C_bl
Rb_63_97 bit_63_97 bit_63_98 R_bl
Rbb_63_97 bitb_63_97 bitb_63_98 R_bl
Cb_63_97 bit_63_97 gnd C_bl
Cbb_63_97 bitb_63_97 gnd C_bl
Rb_63_98 bit_63_98 bit_63_99 R_bl
Rbb_63_98 bitb_63_98 bitb_63_99 R_bl
Cb_63_98 bit_63_98 gnd C_bl
Cbb_63_98 bitb_63_98 gnd C_bl
Rb_63_99 bit_63_99 bit_63_100 R_bl
Rbb_63_99 bitb_63_99 bitb_63_100 R_bl
Cb_63_99 bit_63_99 gnd C_bl
Cbb_63_99 bitb_63_99 gnd C_bl
Rb_64_0 bit_64_0 bit_64_1 R_bl
Rbb_64_0 bitb_64_0 bitb_64_1 R_bl
Cb_64_0 bit_64_0 gnd C_bl
Cbb_64_0 bitb_64_0 gnd C_bl
Rb_64_1 bit_64_1 bit_64_2 R_bl
Rbb_64_1 bitb_64_1 bitb_64_2 R_bl
Cb_64_1 bit_64_1 gnd C_bl
Cbb_64_1 bitb_64_1 gnd C_bl
Rb_64_2 bit_64_2 bit_64_3 R_bl
Rbb_64_2 bitb_64_2 bitb_64_3 R_bl
Cb_64_2 bit_64_2 gnd C_bl
Cbb_64_2 bitb_64_2 gnd C_bl
Rb_64_3 bit_64_3 bit_64_4 R_bl
Rbb_64_3 bitb_64_3 bitb_64_4 R_bl
Cb_64_3 bit_64_3 gnd C_bl
Cbb_64_3 bitb_64_3 gnd C_bl
Rb_64_4 bit_64_4 bit_64_5 R_bl
Rbb_64_4 bitb_64_4 bitb_64_5 R_bl
Cb_64_4 bit_64_4 gnd C_bl
Cbb_64_4 bitb_64_4 gnd C_bl
Rb_64_5 bit_64_5 bit_64_6 R_bl
Rbb_64_5 bitb_64_5 bitb_64_6 R_bl
Cb_64_5 bit_64_5 gnd C_bl
Cbb_64_5 bitb_64_5 gnd C_bl
Rb_64_6 bit_64_6 bit_64_7 R_bl
Rbb_64_6 bitb_64_6 bitb_64_7 R_bl
Cb_64_6 bit_64_6 gnd C_bl
Cbb_64_6 bitb_64_6 gnd C_bl
Rb_64_7 bit_64_7 bit_64_8 R_bl
Rbb_64_7 bitb_64_7 bitb_64_8 R_bl
Cb_64_7 bit_64_7 gnd C_bl
Cbb_64_7 bitb_64_7 gnd C_bl
Rb_64_8 bit_64_8 bit_64_9 R_bl
Rbb_64_8 bitb_64_8 bitb_64_9 R_bl
Cb_64_8 bit_64_8 gnd C_bl
Cbb_64_8 bitb_64_8 gnd C_bl
Rb_64_9 bit_64_9 bit_64_10 R_bl
Rbb_64_9 bitb_64_9 bitb_64_10 R_bl
Cb_64_9 bit_64_9 gnd C_bl
Cbb_64_9 bitb_64_9 gnd C_bl
Rb_64_10 bit_64_10 bit_64_11 R_bl
Rbb_64_10 bitb_64_10 bitb_64_11 R_bl
Cb_64_10 bit_64_10 gnd C_bl
Cbb_64_10 bitb_64_10 gnd C_bl
Rb_64_11 bit_64_11 bit_64_12 R_bl
Rbb_64_11 bitb_64_11 bitb_64_12 R_bl
Cb_64_11 bit_64_11 gnd C_bl
Cbb_64_11 bitb_64_11 gnd C_bl
Rb_64_12 bit_64_12 bit_64_13 R_bl
Rbb_64_12 bitb_64_12 bitb_64_13 R_bl
Cb_64_12 bit_64_12 gnd C_bl
Cbb_64_12 bitb_64_12 gnd C_bl
Rb_64_13 bit_64_13 bit_64_14 R_bl
Rbb_64_13 bitb_64_13 bitb_64_14 R_bl
Cb_64_13 bit_64_13 gnd C_bl
Cbb_64_13 bitb_64_13 gnd C_bl
Rb_64_14 bit_64_14 bit_64_15 R_bl
Rbb_64_14 bitb_64_14 bitb_64_15 R_bl
Cb_64_14 bit_64_14 gnd C_bl
Cbb_64_14 bitb_64_14 gnd C_bl
Rb_64_15 bit_64_15 bit_64_16 R_bl
Rbb_64_15 bitb_64_15 bitb_64_16 R_bl
Cb_64_15 bit_64_15 gnd C_bl
Cbb_64_15 bitb_64_15 gnd C_bl
Rb_64_16 bit_64_16 bit_64_17 R_bl
Rbb_64_16 bitb_64_16 bitb_64_17 R_bl
Cb_64_16 bit_64_16 gnd C_bl
Cbb_64_16 bitb_64_16 gnd C_bl
Rb_64_17 bit_64_17 bit_64_18 R_bl
Rbb_64_17 bitb_64_17 bitb_64_18 R_bl
Cb_64_17 bit_64_17 gnd C_bl
Cbb_64_17 bitb_64_17 gnd C_bl
Rb_64_18 bit_64_18 bit_64_19 R_bl
Rbb_64_18 bitb_64_18 bitb_64_19 R_bl
Cb_64_18 bit_64_18 gnd C_bl
Cbb_64_18 bitb_64_18 gnd C_bl
Rb_64_19 bit_64_19 bit_64_20 R_bl
Rbb_64_19 bitb_64_19 bitb_64_20 R_bl
Cb_64_19 bit_64_19 gnd C_bl
Cbb_64_19 bitb_64_19 gnd C_bl
Rb_64_20 bit_64_20 bit_64_21 R_bl
Rbb_64_20 bitb_64_20 bitb_64_21 R_bl
Cb_64_20 bit_64_20 gnd C_bl
Cbb_64_20 bitb_64_20 gnd C_bl
Rb_64_21 bit_64_21 bit_64_22 R_bl
Rbb_64_21 bitb_64_21 bitb_64_22 R_bl
Cb_64_21 bit_64_21 gnd C_bl
Cbb_64_21 bitb_64_21 gnd C_bl
Rb_64_22 bit_64_22 bit_64_23 R_bl
Rbb_64_22 bitb_64_22 bitb_64_23 R_bl
Cb_64_22 bit_64_22 gnd C_bl
Cbb_64_22 bitb_64_22 gnd C_bl
Rb_64_23 bit_64_23 bit_64_24 R_bl
Rbb_64_23 bitb_64_23 bitb_64_24 R_bl
Cb_64_23 bit_64_23 gnd C_bl
Cbb_64_23 bitb_64_23 gnd C_bl
Rb_64_24 bit_64_24 bit_64_25 R_bl
Rbb_64_24 bitb_64_24 bitb_64_25 R_bl
Cb_64_24 bit_64_24 gnd C_bl
Cbb_64_24 bitb_64_24 gnd C_bl
Rb_64_25 bit_64_25 bit_64_26 R_bl
Rbb_64_25 bitb_64_25 bitb_64_26 R_bl
Cb_64_25 bit_64_25 gnd C_bl
Cbb_64_25 bitb_64_25 gnd C_bl
Rb_64_26 bit_64_26 bit_64_27 R_bl
Rbb_64_26 bitb_64_26 bitb_64_27 R_bl
Cb_64_26 bit_64_26 gnd C_bl
Cbb_64_26 bitb_64_26 gnd C_bl
Rb_64_27 bit_64_27 bit_64_28 R_bl
Rbb_64_27 bitb_64_27 bitb_64_28 R_bl
Cb_64_27 bit_64_27 gnd C_bl
Cbb_64_27 bitb_64_27 gnd C_bl
Rb_64_28 bit_64_28 bit_64_29 R_bl
Rbb_64_28 bitb_64_28 bitb_64_29 R_bl
Cb_64_28 bit_64_28 gnd C_bl
Cbb_64_28 bitb_64_28 gnd C_bl
Rb_64_29 bit_64_29 bit_64_30 R_bl
Rbb_64_29 bitb_64_29 bitb_64_30 R_bl
Cb_64_29 bit_64_29 gnd C_bl
Cbb_64_29 bitb_64_29 gnd C_bl
Rb_64_30 bit_64_30 bit_64_31 R_bl
Rbb_64_30 bitb_64_30 bitb_64_31 R_bl
Cb_64_30 bit_64_30 gnd C_bl
Cbb_64_30 bitb_64_30 gnd C_bl
Rb_64_31 bit_64_31 bit_64_32 R_bl
Rbb_64_31 bitb_64_31 bitb_64_32 R_bl
Cb_64_31 bit_64_31 gnd C_bl
Cbb_64_31 bitb_64_31 gnd C_bl
Rb_64_32 bit_64_32 bit_64_33 R_bl
Rbb_64_32 bitb_64_32 bitb_64_33 R_bl
Cb_64_32 bit_64_32 gnd C_bl
Cbb_64_32 bitb_64_32 gnd C_bl
Rb_64_33 bit_64_33 bit_64_34 R_bl
Rbb_64_33 bitb_64_33 bitb_64_34 R_bl
Cb_64_33 bit_64_33 gnd C_bl
Cbb_64_33 bitb_64_33 gnd C_bl
Rb_64_34 bit_64_34 bit_64_35 R_bl
Rbb_64_34 bitb_64_34 bitb_64_35 R_bl
Cb_64_34 bit_64_34 gnd C_bl
Cbb_64_34 bitb_64_34 gnd C_bl
Rb_64_35 bit_64_35 bit_64_36 R_bl
Rbb_64_35 bitb_64_35 bitb_64_36 R_bl
Cb_64_35 bit_64_35 gnd C_bl
Cbb_64_35 bitb_64_35 gnd C_bl
Rb_64_36 bit_64_36 bit_64_37 R_bl
Rbb_64_36 bitb_64_36 bitb_64_37 R_bl
Cb_64_36 bit_64_36 gnd C_bl
Cbb_64_36 bitb_64_36 gnd C_bl
Rb_64_37 bit_64_37 bit_64_38 R_bl
Rbb_64_37 bitb_64_37 bitb_64_38 R_bl
Cb_64_37 bit_64_37 gnd C_bl
Cbb_64_37 bitb_64_37 gnd C_bl
Rb_64_38 bit_64_38 bit_64_39 R_bl
Rbb_64_38 bitb_64_38 bitb_64_39 R_bl
Cb_64_38 bit_64_38 gnd C_bl
Cbb_64_38 bitb_64_38 gnd C_bl
Rb_64_39 bit_64_39 bit_64_40 R_bl
Rbb_64_39 bitb_64_39 bitb_64_40 R_bl
Cb_64_39 bit_64_39 gnd C_bl
Cbb_64_39 bitb_64_39 gnd C_bl
Rb_64_40 bit_64_40 bit_64_41 R_bl
Rbb_64_40 bitb_64_40 bitb_64_41 R_bl
Cb_64_40 bit_64_40 gnd C_bl
Cbb_64_40 bitb_64_40 gnd C_bl
Rb_64_41 bit_64_41 bit_64_42 R_bl
Rbb_64_41 bitb_64_41 bitb_64_42 R_bl
Cb_64_41 bit_64_41 gnd C_bl
Cbb_64_41 bitb_64_41 gnd C_bl
Rb_64_42 bit_64_42 bit_64_43 R_bl
Rbb_64_42 bitb_64_42 bitb_64_43 R_bl
Cb_64_42 bit_64_42 gnd C_bl
Cbb_64_42 bitb_64_42 gnd C_bl
Rb_64_43 bit_64_43 bit_64_44 R_bl
Rbb_64_43 bitb_64_43 bitb_64_44 R_bl
Cb_64_43 bit_64_43 gnd C_bl
Cbb_64_43 bitb_64_43 gnd C_bl
Rb_64_44 bit_64_44 bit_64_45 R_bl
Rbb_64_44 bitb_64_44 bitb_64_45 R_bl
Cb_64_44 bit_64_44 gnd C_bl
Cbb_64_44 bitb_64_44 gnd C_bl
Rb_64_45 bit_64_45 bit_64_46 R_bl
Rbb_64_45 bitb_64_45 bitb_64_46 R_bl
Cb_64_45 bit_64_45 gnd C_bl
Cbb_64_45 bitb_64_45 gnd C_bl
Rb_64_46 bit_64_46 bit_64_47 R_bl
Rbb_64_46 bitb_64_46 bitb_64_47 R_bl
Cb_64_46 bit_64_46 gnd C_bl
Cbb_64_46 bitb_64_46 gnd C_bl
Rb_64_47 bit_64_47 bit_64_48 R_bl
Rbb_64_47 bitb_64_47 bitb_64_48 R_bl
Cb_64_47 bit_64_47 gnd C_bl
Cbb_64_47 bitb_64_47 gnd C_bl
Rb_64_48 bit_64_48 bit_64_49 R_bl
Rbb_64_48 bitb_64_48 bitb_64_49 R_bl
Cb_64_48 bit_64_48 gnd C_bl
Cbb_64_48 bitb_64_48 gnd C_bl
Rb_64_49 bit_64_49 bit_64_50 R_bl
Rbb_64_49 bitb_64_49 bitb_64_50 R_bl
Cb_64_49 bit_64_49 gnd C_bl
Cbb_64_49 bitb_64_49 gnd C_bl
Rb_64_50 bit_64_50 bit_64_51 R_bl
Rbb_64_50 bitb_64_50 bitb_64_51 R_bl
Cb_64_50 bit_64_50 gnd C_bl
Cbb_64_50 bitb_64_50 gnd C_bl
Rb_64_51 bit_64_51 bit_64_52 R_bl
Rbb_64_51 bitb_64_51 bitb_64_52 R_bl
Cb_64_51 bit_64_51 gnd C_bl
Cbb_64_51 bitb_64_51 gnd C_bl
Rb_64_52 bit_64_52 bit_64_53 R_bl
Rbb_64_52 bitb_64_52 bitb_64_53 R_bl
Cb_64_52 bit_64_52 gnd C_bl
Cbb_64_52 bitb_64_52 gnd C_bl
Rb_64_53 bit_64_53 bit_64_54 R_bl
Rbb_64_53 bitb_64_53 bitb_64_54 R_bl
Cb_64_53 bit_64_53 gnd C_bl
Cbb_64_53 bitb_64_53 gnd C_bl
Rb_64_54 bit_64_54 bit_64_55 R_bl
Rbb_64_54 bitb_64_54 bitb_64_55 R_bl
Cb_64_54 bit_64_54 gnd C_bl
Cbb_64_54 bitb_64_54 gnd C_bl
Rb_64_55 bit_64_55 bit_64_56 R_bl
Rbb_64_55 bitb_64_55 bitb_64_56 R_bl
Cb_64_55 bit_64_55 gnd C_bl
Cbb_64_55 bitb_64_55 gnd C_bl
Rb_64_56 bit_64_56 bit_64_57 R_bl
Rbb_64_56 bitb_64_56 bitb_64_57 R_bl
Cb_64_56 bit_64_56 gnd C_bl
Cbb_64_56 bitb_64_56 gnd C_bl
Rb_64_57 bit_64_57 bit_64_58 R_bl
Rbb_64_57 bitb_64_57 bitb_64_58 R_bl
Cb_64_57 bit_64_57 gnd C_bl
Cbb_64_57 bitb_64_57 gnd C_bl
Rb_64_58 bit_64_58 bit_64_59 R_bl
Rbb_64_58 bitb_64_58 bitb_64_59 R_bl
Cb_64_58 bit_64_58 gnd C_bl
Cbb_64_58 bitb_64_58 gnd C_bl
Rb_64_59 bit_64_59 bit_64_60 R_bl
Rbb_64_59 bitb_64_59 bitb_64_60 R_bl
Cb_64_59 bit_64_59 gnd C_bl
Cbb_64_59 bitb_64_59 gnd C_bl
Rb_64_60 bit_64_60 bit_64_61 R_bl
Rbb_64_60 bitb_64_60 bitb_64_61 R_bl
Cb_64_60 bit_64_60 gnd C_bl
Cbb_64_60 bitb_64_60 gnd C_bl
Rb_64_61 bit_64_61 bit_64_62 R_bl
Rbb_64_61 bitb_64_61 bitb_64_62 R_bl
Cb_64_61 bit_64_61 gnd C_bl
Cbb_64_61 bitb_64_61 gnd C_bl
Rb_64_62 bit_64_62 bit_64_63 R_bl
Rbb_64_62 bitb_64_62 bitb_64_63 R_bl
Cb_64_62 bit_64_62 gnd C_bl
Cbb_64_62 bitb_64_62 gnd C_bl
Rb_64_63 bit_64_63 bit_64_64 R_bl
Rbb_64_63 bitb_64_63 bitb_64_64 R_bl
Cb_64_63 bit_64_63 gnd C_bl
Cbb_64_63 bitb_64_63 gnd C_bl
Rb_64_64 bit_64_64 bit_64_65 R_bl
Rbb_64_64 bitb_64_64 bitb_64_65 R_bl
Cb_64_64 bit_64_64 gnd C_bl
Cbb_64_64 bitb_64_64 gnd C_bl
Rb_64_65 bit_64_65 bit_64_66 R_bl
Rbb_64_65 bitb_64_65 bitb_64_66 R_bl
Cb_64_65 bit_64_65 gnd C_bl
Cbb_64_65 bitb_64_65 gnd C_bl
Rb_64_66 bit_64_66 bit_64_67 R_bl
Rbb_64_66 bitb_64_66 bitb_64_67 R_bl
Cb_64_66 bit_64_66 gnd C_bl
Cbb_64_66 bitb_64_66 gnd C_bl
Rb_64_67 bit_64_67 bit_64_68 R_bl
Rbb_64_67 bitb_64_67 bitb_64_68 R_bl
Cb_64_67 bit_64_67 gnd C_bl
Cbb_64_67 bitb_64_67 gnd C_bl
Rb_64_68 bit_64_68 bit_64_69 R_bl
Rbb_64_68 bitb_64_68 bitb_64_69 R_bl
Cb_64_68 bit_64_68 gnd C_bl
Cbb_64_68 bitb_64_68 gnd C_bl
Rb_64_69 bit_64_69 bit_64_70 R_bl
Rbb_64_69 bitb_64_69 bitb_64_70 R_bl
Cb_64_69 bit_64_69 gnd C_bl
Cbb_64_69 bitb_64_69 gnd C_bl
Rb_64_70 bit_64_70 bit_64_71 R_bl
Rbb_64_70 bitb_64_70 bitb_64_71 R_bl
Cb_64_70 bit_64_70 gnd C_bl
Cbb_64_70 bitb_64_70 gnd C_bl
Rb_64_71 bit_64_71 bit_64_72 R_bl
Rbb_64_71 bitb_64_71 bitb_64_72 R_bl
Cb_64_71 bit_64_71 gnd C_bl
Cbb_64_71 bitb_64_71 gnd C_bl
Rb_64_72 bit_64_72 bit_64_73 R_bl
Rbb_64_72 bitb_64_72 bitb_64_73 R_bl
Cb_64_72 bit_64_72 gnd C_bl
Cbb_64_72 bitb_64_72 gnd C_bl
Rb_64_73 bit_64_73 bit_64_74 R_bl
Rbb_64_73 bitb_64_73 bitb_64_74 R_bl
Cb_64_73 bit_64_73 gnd C_bl
Cbb_64_73 bitb_64_73 gnd C_bl
Rb_64_74 bit_64_74 bit_64_75 R_bl
Rbb_64_74 bitb_64_74 bitb_64_75 R_bl
Cb_64_74 bit_64_74 gnd C_bl
Cbb_64_74 bitb_64_74 gnd C_bl
Rb_64_75 bit_64_75 bit_64_76 R_bl
Rbb_64_75 bitb_64_75 bitb_64_76 R_bl
Cb_64_75 bit_64_75 gnd C_bl
Cbb_64_75 bitb_64_75 gnd C_bl
Rb_64_76 bit_64_76 bit_64_77 R_bl
Rbb_64_76 bitb_64_76 bitb_64_77 R_bl
Cb_64_76 bit_64_76 gnd C_bl
Cbb_64_76 bitb_64_76 gnd C_bl
Rb_64_77 bit_64_77 bit_64_78 R_bl
Rbb_64_77 bitb_64_77 bitb_64_78 R_bl
Cb_64_77 bit_64_77 gnd C_bl
Cbb_64_77 bitb_64_77 gnd C_bl
Rb_64_78 bit_64_78 bit_64_79 R_bl
Rbb_64_78 bitb_64_78 bitb_64_79 R_bl
Cb_64_78 bit_64_78 gnd C_bl
Cbb_64_78 bitb_64_78 gnd C_bl
Rb_64_79 bit_64_79 bit_64_80 R_bl
Rbb_64_79 bitb_64_79 bitb_64_80 R_bl
Cb_64_79 bit_64_79 gnd C_bl
Cbb_64_79 bitb_64_79 gnd C_bl
Rb_64_80 bit_64_80 bit_64_81 R_bl
Rbb_64_80 bitb_64_80 bitb_64_81 R_bl
Cb_64_80 bit_64_80 gnd C_bl
Cbb_64_80 bitb_64_80 gnd C_bl
Rb_64_81 bit_64_81 bit_64_82 R_bl
Rbb_64_81 bitb_64_81 bitb_64_82 R_bl
Cb_64_81 bit_64_81 gnd C_bl
Cbb_64_81 bitb_64_81 gnd C_bl
Rb_64_82 bit_64_82 bit_64_83 R_bl
Rbb_64_82 bitb_64_82 bitb_64_83 R_bl
Cb_64_82 bit_64_82 gnd C_bl
Cbb_64_82 bitb_64_82 gnd C_bl
Rb_64_83 bit_64_83 bit_64_84 R_bl
Rbb_64_83 bitb_64_83 bitb_64_84 R_bl
Cb_64_83 bit_64_83 gnd C_bl
Cbb_64_83 bitb_64_83 gnd C_bl
Rb_64_84 bit_64_84 bit_64_85 R_bl
Rbb_64_84 bitb_64_84 bitb_64_85 R_bl
Cb_64_84 bit_64_84 gnd C_bl
Cbb_64_84 bitb_64_84 gnd C_bl
Rb_64_85 bit_64_85 bit_64_86 R_bl
Rbb_64_85 bitb_64_85 bitb_64_86 R_bl
Cb_64_85 bit_64_85 gnd C_bl
Cbb_64_85 bitb_64_85 gnd C_bl
Rb_64_86 bit_64_86 bit_64_87 R_bl
Rbb_64_86 bitb_64_86 bitb_64_87 R_bl
Cb_64_86 bit_64_86 gnd C_bl
Cbb_64_86 bitb_64_86 gnd C_bl
Rb_64_87 bit_64_87 bit_64_88 R_bl
Rbb_64_87 bitb_64_87 bitb_64_88 R_bl
Cb_64_87 bit_64_87 gnd C_bl
Cbb_64_87 bitb_64_87 gnd C_bl
Rb_64_88 bit_64_88 bit_64_89 R_bl
Rbb_64_88 bitb_64_88 bitb_64_89 R_bl
Cb_64_88 bit_64_88 gnd C_bl
Cbb_64_88 bitb_64_88 gnd C_bl
Rb_64_89 bit_64_89 bit_64_90 R_bl
Rbb_64_89 bitb_64_89 bitb_64_90 R_bl
Cb_64_89 bit_64_89 gnd C_bl
Cbb_64_89 bitb_64_89 gnd C_bl
Rb_64_90 bit_64_90 bit_64_91 R_bl
Rbb_64_90 bitb_64_90 bitb_64_91 R_bl
Cb_64_90 bit_64_90 gnd C_bl
Cbb_64_90 bitb_64_90 gnd C_bl
Rb_64_91 bit_64_91 bit_64_92 R_bl
Rbb_64_91 bitb_64_91 bitb_64_92 R_bl
Cb_64_91 bit_64_91 gnd C_bl
Cbb_64_91 bitb_64_91 gnd C_bl
Rb_64_92 bit_64_92 bit_64_93 R_bl
Rbb_64_92 bitb_64_92 bitb_64_93 R_bl
Cb_64_92 bit_64_92 gnd C_bl
Cbb_64_92 bitb_64_92 gnd C_bl
Rb_64_93 bit_64_93 bit_64_94 R_bl
Rbb_64_93 bitb_64_93 bitb_64_94 R_bl
Cb_64_93 bit_64_93 gnd C_bl
Cbb_64_93 bitb_64_93 gnd C_bl
Rb_64_94 bit_64_94 bit_64_95 R_bl
Rbb_64_94 bitb_64_94 bitb_64_95 R_bl
Cb_64_94 bit_64_94 gnd C_bl
Cbb_64_94 bitb_64_94 gnd C_bl
Rb_64_95 bit_64_95 bit_64_96 R_bl
Rbb_64_95 bitb_64_95 bitb_64_96 R_bl
Cb_64_95 bit_64_95 gnd C_bl
Cbb_64_95 bitb_64_95 gnd C_bl
Rb_64_96 bit_64_96 bit_64_97 R_bl
Rbb_64_96 bitb_64_96 bitb_64_97 R_bl
Cb_64_96 bit_64_96 gnd C_bl
Cbb_64_96 bitb_64_96 gnd C_bl
Rb_64_97 bit_64_97 bit_64_98 R_bl
Rbb_64_97 bitb_64_97 bitb_64_98 R_bl
Cb_64_97 bit_64_97 gnd C_bl
Cbb_64_97 bitb_64_97 gnd C_bl
Rb_64_98 bit_64_98 bit_64_99 R_bl
Rbb_64_98 bitb_64_98 bitb_64_99 R_bl
Cb_64_98 bit_64_98 gnd C_bl
Cbb_64_98 bitb_64_98 gnd C_bl
Rb_64_99 bit_64_99 bit_64_100 R_bl
Rbb_64_99 bitb_64_99 bitb_64_100 R_bl
Cb_64_99 bit_64_99 gnd C_bl
Cbb_64_99 bitb_64_99 gnd C_bl
Rb_65_0 bit_65_0 bit_65_1 R_bl
Rbb_65_0 bitb_65_0 bitb_65_1 R_bl
Cb_65_0 bit_65_0 gnd C_bl
Cbb_65_0 bitb_65_0 gnd C_bl
Rb_65_1 bit_65_1 bit_65_2 R_bl
Rbb_65_1 bitb_65_1 bitb_65_2 R_bl
Cb_65_1 bit_65_1 gnd C_bl
Cbb_65_1 bitb_65_1 gnd C_bl
Rb_65_2 bit_65_2 bit_65_3 R_bl
Rbb_65_2 bitb_65_2 bitb_65_3 R_bl
Cb_65_2 bit_65_2 gnd C_bl
Cbb_65_2 bitb_65_2 gnd C_bl
Rb_65_3 bit_65_3 bit_65_4 R_bl
Rbb_65_3 bitb_65_3 bitb_65_4 R_bl
Cb_65_3 bit_65_3 gnd C_bl
Cbb_65_3 bitb_65_3 gnd C_bl
Rb_65_4 bit_65_4 bit_65_5 R_bl
Rbb_65_4 bitb_65_4 bitb_65_5 R_bl
Cb_65_4 bit_65_4 gnd C_bl
Cbb_65_4 bitb_65_4 gnd C_bl
Rb_65_5 bit_65_5 bit_65_6 R_bl
Rbb_65_5 bitb_65_5 bitb_65_6 R_bl
Cb_65_5 bit_65_5 gnd C_bl
Cbb_65_5 bitb_65_5 gnd C_bl
Rb_65_6 bit_65_6 bit_65_7 R_bl
Rbb_65_6 bitb_65_6 bitb_65_7 R_bl
Cb_65_6 bit_65_6 gnd C_bl
Cbb_65_6 bitb_65_6 gnd C_bl
Rb_65_7 bit_65_7 bit_65_8 R_bl
Rbb_65_7 bitb_65_7 bitb_65_8 R_bl
Cb_65_7 bit_65_7 gnd C_bl
Cbb_65_7 bitb_65_7 gnd C_bl
Rb_65_8 bit_65_8 bit_65_9 R_bl
Rbb_65_8 bitb_65_8 bitb_65_9 R_bl
Cb_65_8 bit_65_8 gnd C_bl
Cbb_65_8 bitb_65_8 gnd C_bl
Rb_65_9 bit_65_9 bit_65_10 R_bl
Rbb_65_9 bitb_65_9 bitb_65_10 R_bl
Cb_65_9 bit_65_9 gnd C_bl
Cbb_65_9 bitb_65_9 gnd C_bl
Rb_65_10 bit_65_10 bit_65_11 R_bl
Rbb_65_10 bitb_65_10 bitb_65_11 R_bl
Cb_65_10 bit_65_10 gnd C_bl
Cbb_65_10 bitb_65_10 gnd C_bl
Rb_65_11 bit_65_11 bit_65_12 R_bl
Rbb_65_11 bitb_65_11 bitb_65_12 R_bl
Cb_65_11 bit_65_11 gnd C_bl
Cbb_65_11 bitb_65_11 gnd C_bl
Rb_65_12 bit_65_12 bit_65_13 R_bl
Rbb_65_12 bitb_65_12 bitb_65_13 R_bl
Cb_65_12 bit_65_12 gnd C_bl
Cbb_65_12 bitb_65_12 gnd C_bl
Rb_65_13 bit_65_13 bit_65_14 R_bl
Rbb_65_13 bitb_65_13 bitb_65_14 R_bl
Cb_65_13 bit_65_13 gnd C_bl
Cbb_65_13 bitb_65_13 gnd C_bl
Rb_65_14 bit_65_14 bit_65_15 R_bl
Rbb_65_14 bitb_65_14 bitb_65_15 R_bl
Cb_65_14 bit_65_14 gnd C_bl
Cbb_65_14 bitb_65_14 gnd C_bl
Rb_65_15 bit_65_15 bit_65_16 R_bl
Rbb_65_15 bitb_65_15 bitb_65_16 R_bl
Cb_65_15 bit_65_15 gnd C_bl
Cbb_65_15 bitb_65_15 gnd C_bl
Rb_65_16 bit_65_16 bit_65_17 R_bl
Rbb_65_16 bitb_65_16 bitb_65_17 R_bl
Cb_65_16 bit_65_16 gnd C_bl
Cbb_65_16 bitb_65_16 gnd C_bl
Rb_65_17 bit_65_17 bit_65_18 R_bl
Rbb_65_17 bitb_65_17 bitb_65_18 R_bl
Cb_65_17 bit_65_17 gnd C_bl
Cbb_65_17 bitb_65_17 gnd C_bl
Rb_65_18 bit_65_18 bit_65_19 R_bl
Rbb_65_18 bitb_65_18 bitb_65_19 R_bl
Cb_65_18 bit_65_18 gnd C_bl
Cbb_65_18 bitb_65_18 gnd C_bl
Rb_65_19 bit_65_19 bit_65_20 R_bl
Rbb_65_19 bitb_65_19 bitb_65_20 R_bl
Cb_65_19 bit_65_19 gnd C_bl
Cbb_65_19 bitb_65_19 gnd C_bl
Rb_65_20 bit_65_20 bit_65_21 R_bl
Rbb_65_20 bitb_65_20 bitb_65_21 R_bl
Cb_65_20 bit_65_20 gnd C_bl
Cbb_65_20 bitb_65_20 gnd C_bl
Rb_65_21 bit_65_21 bit_65_22 R_bl
Rbb_65_21 bitb_65_21 bitb_65_22 R_bl
Cb_65_21 bit_65_21 gnd C_bl
Cbb_65_21 bitb_65_21 gnd C_bl
Rb_65_22 bit_65_22 bit_65_23 R_bl
Rbb_65_22 bitb_65_22 bitb_65_23 R_bl
Cb_65_22 bit_65_22 gnd C_bl
Cbb_65_22 bitb_65_22 gnd C_bl
Rb_65_23 bit_65_23 bit_65_24 R_bl
Rbb_65_23 bitb_65_23 bitb_65_24 R_bl
Cb_65_23 bit_65_23 gnd C_bl
Cbb_65_23 bitb_65_23 gnd C_bl
Rb_65_24 bit_65_24 bit_65_25 R_bl
Rbb_65_24 bitb_65_24 bitb_65_25 R_bl
Cb_65_24 bit_65_24 gnd C_bl
Cbb_65_24 bitb_65_24 gnd C_bl
Rb_65_25 bit_65_25 bit_65_26 R_bl
Rbb_65_25 bitb_65_25 bitb_65_26 R_bl
Cb_65_25 bit_65_25 gnd C_bl
Cbb_65_25 bitb_65_25 gnd C_bl
Rb_65_26 bit_65_26 bit_65_27 R_bl
Rbb_65_26 bitb_65_26 bitb_65_27 R_bl
Cb_65_26 bit_65_26 gnd C_bl
Cbb_65_26 bitb_65_26 gnd C_bl
Rb_65_27 bit_65_27 bit_65_28 R_bl
Rbb_65_27 bitb_65_27 bitb_65_28 R_bl
Cb_65_27 bit_65_27 gnd C_bl
Cbb_65_27 bitb_65_27 gnd C_bl
Rb_65_28 bit_65_28 bit_65_29 R_bl
Rbb_65_28 bitb_65_28 bitb_65_29 R_bl
Cb_65_28 bit_65_28 gnd C_bl
Cbb_65_28 bitb_65_28 gnd C_bl
Rb_65_29 bit_65_29 bit_65_30 R_bl
Rbb_65_29 bitb_65_29 bitb_65_30 R_bl
Cb_65_29 bit_65_29 gnd C_bl
Cbb_65_29 bitb_65_29 gnd C_bl
Rb_65_30 bit_65_30 bit_65_31 R_bl
Rbb_65_30 bitb_65_30 bitb_65_31 R_bl
Cb_65_30 bit_65_30 gnd C_bl
Cbb_65_30 bitb_65_30 gnd C_bl
Rb_65_31 bit_65_31 bit_65_32 R_bl
Rbb_65_31 bitb_65_31 bitb_65_32 R_bl
Cb_65_31 bit_65_31 gnd C_bl
Cbb_65_31 bitb_65_31 gnd C_bl
Rb_65_32 bit_65_32 bit_65_33 R_bl
Rbb_65_32 bitb_65_32 bitb_65_33 R_bl
Cb_65_32 bit_65_32 gnd C_bl
Cbb_65_32 bitb_65_32 gnd C_bl
Rb_65_33 bit_65_33 bit_65_34 R_bl
Rbb_65_33 bitb_65_33 bitb_65_34 R_bl
Cb_65_33 bit_65_33 gnd C_bl
Cbb_65_33 bitb_65_33 gnd C_bl
Rb_65_34 bit_65_34 bit_65_35 R_bl
Rbb_65_34 bitb_65_34 bitb_65_35 R_bl
Cb_65_34 bit_65_34 gnd C_bl
Cbb_65_34 bitb_65_34 gnd C_bl
Rb_65_35 bit_65_35 bit_65_36 R_bl
Rbb_65_35 bitb_65_35 bitb_65_36 R_bl
Cb_65_35 bit_65_35 gnd C_bl
Cbb_65_35 bitb_65_35 gnd C_bl
Rb_65_36 bit_65_36 bit_65_37 R_bl
Rbb_65_36 bitb_65_36 bitb_65_37 R_bl
Cb_65_36 bit_65_36 gnd C_bl
Cbb_65_36 bitb_65_36 gnd C_bl
Rb_65_37 bit_65_37 bit_65_38 R_bl
Rbb_65_37 bitb_65_37 bitb_65_38 R_bl
Cb_65_37 bit_65_37 gnd C_bl
Cbb_65_37 bitb_65_37 gnd C_bl
Rb_65_38 bit_65_38 bit_65_39 R_bl
Rbb_65_38 bitb_65_38 bitb_65_39 R_bl
Cb_65_38 bit_65_38 gnd C_bl
Cbb_65_38 bitb_65_38 gnd C_bl
Rb_65_39 bit_65_39 bit_65_40 R_bl
Rbb_65_39 bitb_65_39 bitb_65_40 R_bl
Cb_65_39 bit_65_39 gnd C_bl
Cbb_65_39 bitb_65_39 gnd C_bl
Rb_65_40 bit_65_40 bit_65_41 R_bl
Rbb_65_40 bitb_65_40 bitb_65_41 R_bl
Cb_65_40 bit_65_40 gnd C_bl
Cbb_65_40 bitb_65_40 gnd C_bl
Rb_65_41 bit_65_41 bit_65_42 R_bl
Rbb_65_41 bitb_65_41 bitb_65_42 R_bl
Cb_65_41 bit_65_41 gnd C_bl
Cbb_65_41 bitb_65_41 gnd C_bl
Rb_65_42 bit_65_42 bit_65_43 R_bl
Rbb_65_42 bitb_65_42 bitb_65_43 R_bl
Cb_65_42 bit_65_42 gnd C_bl
Cbb_65_42 bitb_65_42 gnd C_bl
Rb_65_43 bit_65_43 bit_65_44 R_bl
Rbb_65_43 bitb_65_43 bitb_65_44 R_bl
Cb_65_43 bit_65_43 gnd C_bl
Cbb_65_43 bitb_65_43 gnd C_bl
Rb_65_44 bit_65_44 bit_65_45 R_bl
Rbb_65_44 bitb_65_44 bitb_65_45 R_bl
Cb_65_44 bit_65_44 gnd C_bl
Cbb_65_44 bitb_65_44 gnd C_bl
Rb_65_45 bit_65_45 bit_65_46 R_bl
Rbb_65_45 bitb_65_45 bitb_65_46 R_bl
Cb_65_45 bit_65_45 gnd C_bl
Cbb_65_45 bitb_65_45 gnd C_bl
Rb_65_46 bit_65_46 bit_65_47 R_bl
Rbb_65_46 bitb_65_46 bitb_65_47 R_bl
Cb_65_46 bit_65_46 gnd C_bl
Cbb_65_46 bitb_65_46 gnd C_bl
Rb_65_47 bit_65_47 bit_65_48 R_bl
Rbb_65_47 bitb_65_47 bitb_65_48 R_bl
Cb_65_47 bit_65_47 gnd C_bl
Cbb_65_47 bitb_65_47 gnd C_bl
Rb_65_48 bit_65_48 bit_65_49 R_bl
Rbb_65_48 bitb_65_48 bitb_65_49 R_bl
Cb_65_48 bit_65_48 gnd C_bl
Cbb_65_48 bitb_65_48 gnd C_bl
Rb_65_49 bit_65_49 bit_65_50 R_bl
Rbb_65_49 bitb_65_49 bitb_65_50 R_bl
Cb_65_49 bit_65_49 gnd C_bl
Cbb_65_49 bitb_65_49 gnd C_bl
Rb_65_50 bit_65_50 bit_65_51 R_bl
Rbb_65_50 bitb_65_50 bitb_65_51 R_bl
Cb_65_50 bit_65_50 gnd C_bl
Cbb_65_50 bitb_65_50 gnd C_bl
Rb_65_51 bit_65_51 bit_65_52 R_bl
Rbb_65_51 bitb_65_51 bitb_65_52 R_bl
Cb_65_51 bit_65_51 gnd C_bl
Cbb_65_51 bitb_65_51 gnd C_bl
Rb_65_52 bit_65_52 bit_65_53 R_bl
Rbb_65_52 bitb_65_52 bitb_65_53 R_bl
Cb_65_52 bit_65_52 gnd C_bl
Cbb_65_52 bitb_65_52 gnd C_bl
Rb_65_53 bit_65_53 bit_65_54 R_bl
Rbb_65_53 bitb_65_53 bitb_65_54 R_bl
Cb_65_53 bit_65_53 gnd C_bl
Cbb_65_53 bitb_65_53 gnd C_bl
Rb_65_54 bit_65_54 bit_65_55 R_bl
Rbb_65_54 bitb_65_54 bitb_65_55 R_bl
Cb_65_54 bit_65_54 gnd C_bl
Cbb_65_54 bitb_65_54 gnd C_bl
Rb_65_55 bit_65_55 bit_65_56 R_bl
Rbb_65_55 bitb_65_55 bitb_65_56 R_bl
Cb_65_55 bit_65_55 gnd C_bl
Cbb_65_55 bitb_65_55 gnd C_bl
Rb_65_56 bit_65_56 bit_65_57 R_bl
Rbb_65_56 bitb_65_56 bitb_65_57 R_bl
Cb_65_56 bit_65_56 gnd C_bl
Cbb_65_56 bitb_65_56 gnd C_bl
Rb_65_57 bit_65_57 bit_65_58 R_bl
Rbb_65_57 bitb_65_57 bitb_65_58 R_bl
Cb_65_57 bit_65_57 gnd C_bl
Cbb_65_57 bitb_65_57 gnd C_bl
Rb_65_58 bit_65_58 bit_65_59 R_bl
Rbb_65_58 bitb_65_58 bitb_65_59 R_bl
Cb_65_58 bit_65_58 gnd C_bl
Cbb_65_58 bitb_65_58 gnd C_bl
Rb_65_59 bit_65_59 bit_65_60 R_bl
Rbb_65_59 bitb_65_59 bitb_65_60 R_bl
Cb_65_59 bit_65_59 gnd C_bl
Cbb_65_59 bitb_65_59 gnd C_bl
Rb_65_60 bit_65_60 bit_65_61 R_bl
Rbb_65_60 bitb_65_60 bitb_65_61 R_bl
Cb_65_60 bit_65_60 gnd C_bl
Cbb_65_60 bitb_65_60 gnd C_bl
Rb_65_61 bit_65_61 bit_65_62 R_bl
Rbb_65_61 bitb_65_61 bitb_65_62 R_bl
Cb_65_61 bit_65_61 gnd C_bl
Cbb_65_61 bitb_65_61 gnd C_bl
Rb_65_62 bit_65_62 bit_65_63 R_bl
Rbb_65_62 bitb_65_62 bitb_65_63 R_bl
Cb_65_62 bit_65_62 gnd C_bl
Cbb_65_62 bitb_65_62 gnd C_bl
Rb_65_63 bit_65_63 bit_65_64 R_bl
Rbb_65_63 bitb_65_63 bitb_65_64 R_bl
Cb_65_63 bit_65_63 gnd C_bl
Cbb_65_63 bitb_65_63 gnd C_bl
Rb_65_64 bit_65_64 bit_65_65 R_bl
Rbb_65_64 bitb_65_64 bitb_65_65 R_bl
Cb_65_64 bit_65_64 gnd C_bl
Cbb_65_64 bitb_65_64 gnd C_bl
Rb_65_65 bit_65_65 bit_65_66 R_bl
Rbb_65_65 bitb_65_65 bitb_65_66 R_bl
Cb_65_65 bit_65_65 gnd C_bl
Cbb_65_65 bitb_65_65 gnd C_bl
Rb_65_66 bit_65_66 bit_65_67 R_bl
Rbb_65_66 bitb_65_66 bitb_65_67 R_bl
Cb_65_66 bit_65_66 gnd C_bl
Cbb_65_66 bitb_65_66 gnd C_bl
Rb_65_67 bit_65_67 bit_65_68 R_bl
Rbb_65_67 bitb_65_67 bitb_65_68 R_bl
Cb_65_67 bit_65_67 gnd C_bl
Cbb_65_67 bitb_65_67 gnd C_bl
Rb_65_68 bit_65_68 bit_65_69 R_bl
Rbb_65_68 bitb_65_68 bitb_65_69 R_bl
Cb_65_68 bit_65_68 gnd C_bl
Cbb_65_68 bitb_65_68 gnd C_bl
Rb_65_69 bit_65_69 bit_65_70 R_bl
Rbb_65_69 bitb_65_69 bitb_65_70 R_bl
Cb_65_69 bit_65_69 gnd C_bl
Cbb_65_69 bitb_65_69 gnd C_bl
Rb_65_70 bit_65_70 bit_65_71 R_bl
Rbb_65_70 bitb_65_70 bitb_65_71 R_bl
Cb_65_70 bit_65_70 gnd C_bl
Cbb_65_70 bitb_65_70 gnd C_bl
Rb_65_71 bit_65_71 bit_65_72 R_bl
Rbb_65_71 bitb_65_71 bitb_65_72 R_bl
Cb_65_71 bit_65_71 gnd C_bl
Cbb_65_71 bitb_65_71 gnd C_bl
Rb_65_72 bit_65_72 bit_65_73 R_bl
Rbb_65_72 bitb_65_72 bitb_65_73 R_bl
Cb_65_72 bit_65_72 gnd C_bl
Cbb_65_72 bitb_65_72 gnd C_bl
Rb_65_73 bit_65_73 bit_65_74 R_bl
Rbb_65_73 bitb_65_73 bitb_65_74 R_bl
Cb_65_73 bit_65_73 gnd C_bl
Cbb_65_73 bitb_65_73 gnd C_bl
Rb_65_74 bit_65_74 bit_65_75 R_bl
Rbb_65_74 bitb_65_74 bitb_65_75 R_bl
Cb_65_74 bit_65_74 gnd C_bl
Cbb_65_74 bitb_65_74 gnd C_bl
Rb_65_75 bit_65_75 bit_65_76 R_bl
Rbb_65_75 bitb_65_75 bitb_65_76 R_bl
Cb_65_75 bit_65_75 gnd C_bl
Cbb_65_75 bitb_65_75 gnd C_bl
Rb_65_76 bit_65_76 bit_65_77 R_bl
Rbb_65_76 bitb_65_76 bitb_65_77 R_bl
Cb_65_76 bit_65_76 gnd C_bl
Cbb_65_76 bitb_65_76 gnd C_bl
Rb_65_77 bit_65_77 bit_65_78 R_bl
Rbb_65_77 bitb_65_77 bitb_65_78 R_bl
Cb_65_77 bit_65_77 gnd C_bl
Cbb_65_77 bitb_65_77 gnd C_bl
Rb_65_78 bit_65_78 bit_65_79 R_bl
Rbb_65_78 bitb_65_78 bitb_65_79 R_bl
Cb_65_78 bit_65_78 gnd C_bl
Cbb_65_78 bitb_65_78 gnd C_bl
Rb_65_79 bit_65_79 bit_65_80 R_bl
Rbb_65_79 bitb_65_79 bitb_65_80 R_bl
Cb_65_79 bit_65_79 gnd C_bl
Cbb_65_79 bitb_65_79 gnd C_bl
Rb_65_80 bit_65_80 bit_65_81 R_bl
Rbb_65_80 bitb_65_80 bitb_65_81 R_bl
Cb_65_80 bit_65_80 gnd C_bl
Cbb_65_80 bitb_65_80 gnd C_bl
Rb_65_81 bit_65_81 bit_65_82 R_bl
Rbb_65_81 bitb_65_81 bitb_65_82 R_bl
Cb_65_81 bit_65_81 gnd C_bl
Cbb_65_81 bitb_65_81 gnd C_bl
Rb_65_82 bit_65_82 bit_65_83 R_bl
Rbb_65_82 bitb_65_82 bitb_65_83 R_bl
Cb_65_82 bit_65_82 gnd C_bl
Cbb_65_82 bitb_65_82 gnd C_bl
Rb_65_83 bit_65_83 bit_65_84 R_bl
Rbb_65_83 bitb_65_83 bitb_65_84 R_bl
Cb_65_83 bit_65_83 gnd C_bl
Cbb_65_83 bitb_65_83 gnd C_bl
Rb_65_84 bit_65_84 bit_65_85 R_bl
Rbb_65_84 bitb_65_84 bitb_65_85 R_bl
Cb_65_84 bit_65_84 gnd C_bl
Cbb_65_84 bitb_65_84 gnd C_bl
Rb_65_85 bit_65_85 bit_65_86 R_bl
Rbb_65_85 bitb_65_85 bitb_65_86 R_bl
Cb_65_85 bit_65_85 gnd C_bl
Cbb_65_85 bitb_65_85 gnd C_bl
Rb_65_86 bit_65_86 bit_65_87 R_bl
Rbb_65_86 bitb_65_86 bitb_65_87 R_bl
Cb_65_86 bit_65_86 gnd C_bl
Cbb_65_86 bitb_65_86 gnd C_bl
Rb_65_87 bit_65_87 bit_65_88 R_bl
Rbb_65_87 bitb_65_87 bitb_65_88 R_bl
Cb_65_87 bit_65_87 gnd C_bl
Cbb_65_87 bitb_65_87 gnd C_bl
Rb_65_88 bit_65_88 bit_65_89 R_bl
Rbb_65_88 bitb_65_88 bitb_65_89 R_bl
Cb_65_88 bit_65_88 gnd C_bl
Cbb_65_88 bitb_65_88 gnd C_bl
Rb_65_89 bit_65_89 bit_65_90 R_bl
Rbb_65_89 bitb_65_89 bitb_65_90 R_bl
Cb_65_89 bit_65_89 gnd C_bl
Cbb_65_89 bitb_65_89 gnd C_bl
Rb_65_90 bit_65_90 bit_65_91 R_bl
Rbb_65_90 bitb_65_90 bitb_65_91 R_bl
Cb_65_90 bit_65_90 gnd C_bl
Cbb_65_90 bitb_65_90 gnd C_bl
Rb_65_91 bit_65_91 bit_65_92 R_bl
Rbb_65_91 bitb_65_91 bitb_65_92 R_bl
Cb_65_91 bit_65_91 gnd C_bl
Cbb_65_91 bitb_65_91 gnd C_bl
Rb_65_92 bit_65_92 bit_65_93 R_bl
Rbb_65_92 bitb_65_92 bitb_65_93 R_bl
Cb_65_92 bit_65_92 gnd C_bl
Cbb_65_92 bitb_65_92 gnd C_bl
Rb_65_93 bit_65_93 bit_65_94 R_bl
Rbb_65_93 bitb_65_93 bitb_65_94 R_bl
Cb_65_93 bit_65_93 gnd C_bl
Cbb_65_93 bitb_65_93 gnd C_bl
Rb_65_94 bit_65_94 bit_65_95 R_bl
Rbb_65_94 bitb_65_94 bitb_65_95 R_bl
Cb_65_94 bit_65_94 gnd C_bl
Cbb_65_94 bitb_65_94 gnd C_bl
Rb_65_95 bit_65_95 bit_65_96 R_bl
Rbb_65_95 bitb_65_95 bitb_65_96 R_bl
Cb_65_95 bit_65_95 gnd C_bl
Cbb_65_95 bitb_65_95 gnd C_bl
Rb_65_96 bit_65_96 bit_65_97 R_bl
Rbb_65_96 bitb_65_96 bitb_65_97 R_bl
Cb_65_96 bit_65_96 gnd C_bl
Cbb_65_96 bitb_65_96 gnd C_bl
Rb_65_97 bit_65_97 bit_65_98 R_bl
Rbb_65_97 bitb_65_97 bitb_65_98 R_bl
Cb_65_97 bit_65_97 gnd C_bl
Cbb_65_97 bitb_65_97 gnd C_bl
Rb_65_98 bit_65_98 bit_65_99 R_bl
Rbb_65_98 bitb_65_98 bitb_65_99 R_bl
Cb_65_98 bit_65_98 gnd C_bl
Cbb_65_98 bitb_65_98 gnd C_bl
Rb_65_99 bit_65_99 bit_65_100 R_bl
Rbb_65_99 bitb_65_99 bitb_65_100 R_bl
Cb_65_99 bit_65_99 gnd C_bl
Cbb_65_99 bitb_65_99 gnd C_bl
Rb_66_0 bit_66_0 bit_66_1 R_bl
Rbb_66_0 bitb_66_0 bitb_66_1 R_bl
Cb_66_0 bit_66_0 gnd C_bl
Cbb_66_0 bitb_66_0 gnd C_bl
Rb_66_1 bit_66_1 bit_66_2 R_bl
Rbb_66_1 bitb_66_1 bitb_66_2 R_bl
Cb_66_1 bit_66_1 gnd C_bl
Cbb_66_1 bitb_66_1 gnd C_bl
Rb_66_2 bit_66_2 bit_66_3 R_bl
Rbb_66_2 bitb_66_2 bitb_66_3 R_bl
Cb_66_2 bit_66_2 gnd C_bl
Cbb_66_2 bitb_66_2 gnd C_bl
Rb_66_3 bit_66_3 bit_66_4 R_bl
Rbb_66_3 bitb_66_3 bitb_66_4 R_bl
Cb_66_3 bit_66_3 gnd C_bl
Cbb_66_3 bitb_66_3 gnd C_bl
Rb_66_4 bit_66_4 bit_66_5 R_bl
Rbb_66_4 bitb_66_4 bitb_66_5 R_bl
Cb_66_4 bit_66_4 gnd C_bl
Cbb_66_4 bitb_66_4 gnd C_bl
Rb_66_5 bit_66_5 bit_66_6 R_bl
Rbb_66_5 bitb_66_5 bitb_66_6 R_bl
Cb_66_5 bit_66_5 gnd C_bl
Cbb_66_5 bitb_66_5 gnd C_bl
Rb_66_6 bit_66_6 bit_66_7 R_bl
Rbb_66_6 bitb_66_6 bitb_66_7 R_bl
Cb_66_6 bit_66_6 gnd C_bl
Cbb_66_6 bitb_66_6 gnd C_bl
Rb_66_7 bit_66_7 bit_66_8 R_bl
Rbb_66_7 bitb_66_7 bitb_66_8 R_bl
Cb_66_7 bit_66_7 gnd C_bl
Cbb_66_7 bitb_66_7 gnd C_bl
Rb_66_8 bit_66_8 bit_66_9 R_bl
Rbb_66_8 bitb_66_8 bitb_66_9 R_bl
Cb_66_8 bit_66_8 gnd C_bl
Cbb_66_8 bitb_66_8 gnd C_bl
Rb_66_9 bit_66_9 bit_66_10 R_bl
Rbb_66_9 bitb_66_9 bitb_66_10 R_bl
Cb_66_9 bit_66_9 gnd C_bl
Cbb_66_9 bitb_66_9 gnd C_bl
Rb_66_10 bit_66_10 bit_66_11 R_bl
Rbb_66_10 bitb_66_10 bitb_66_11 R_bl
Cb_66_10 bit_66_10 gnd C_bl
Cbb_66_10 bitb_66_10 gnd C_bl
Rb_66_11 bit_66_11 bit_66_12 R_bl
Rbb_66_11 bitb_66_11 bitb_66_12 R_bl
Cb_66_11 bit_66_11 gnd C_bl
Cbb_66_11 bitb_66_11 gnd C_bl
Rb_66_12 bit_66_12 bit_66_13 R_bl
Rbb_66_12 bitb_66_12 bitb_66_13 R_bl
Cb_66_12 bit_66_12 gnd C_bl
Cbb_66_12 bitb_66_12 gnd C_bl
Rb_66_13 bit_66_13 bit_66_14 R_bl
Rbb_66_13 bitb_66_13 bitb_66_14 R_bl
Cb_66_13 bit_66_13 gnd C_bl
Cbb_66_13 bitb_66_13 gnd C_bl
Rb_66_14 bit_66_14 bit_66_15 R_bl
Rbb_66_14 bitb_66_14 bitb_66_15 R_bl
Cb_66_14 bit_66_14 gnd C_bl
Cbb_66_14 bitb_66_14 gnd C_bl
Rb_66_15 bit_66_15 bit_66_16 R_bl
Rbb_66_15 bitb_66_15 bitb_66_16 R_bl
Cb_66_15 bit_66_15 gnd C_bl
Cbb_66_15 bitb_66_15 gnd C_bl
Rb_66_16 bit_66_16 bit_66_17 R_bl
Rbb_66_16 bitb_66_16 bitb_66_17 R_bl
Cb_66_16 bit_66_16 gnd C_bl
Cbb_66_16 bitb_66_16 gnd C_bl
Rb_66_17 bit_66_17 bit_66_18 R_bl
Rbb_66_17 bitb_66_17 bitb_66_18 R_bl
Cb_66_17 bit_66_17 gnd C_bl
Cbb_66_17 bitb_66_17 gnd C_bl
Rb_66_18 bit_66_18 bit_66_19 R_bl
Rbb_66_18 bitb_66_18 bitb_66_19 R_bl
Cb_66_18 bit_66_18 gnd C_bl
Cbb_66_18 bitb_66_18 gnd C_bl
Rb_66_19 bit_66_19 bit_66_20 R_bl
Rbb_66_19 bitb_66_19 bitb_66_20 R_bl
Cb_66_19 bit_66_19 gnd C_bl
Cbb_66_19 bitb_66_19 gnd C_bl
Rb_66_20 bit_66_20 bit_66_21 R_bl
Rbb_66_20 bitb_66_20 bitb_66_21 R_bl
Cb_66_20 bit_66_20 gnd C_bl
Cbb_66_20 bitb_66_20 gnd C_bl
Rb_66_21 bit_66_21 bit_66_22 R_bl
Rbb_66_21 bitb_66_21 bitb_66_22 R_bl
Cb_66_21 bit_66_21 gnd C_bl
Cbb_66_21 bitb_66_21 gnd C_bl
Rb_66_22 bit_66_22 bit_66_23 R_bl
Rbb_66_22 bitb_66_22 bitb_66_23 R_bl
Cb_66_22 bit_66_22 gnd C_bl
Cbb_66_22 bitb_66_22 gnd C_bl
Rb_66_23 bit_66_23 bit_66_24 R_bl
Rbb_66_23 bitb_66_23 bitb_66_24 R_bl
Cb_66_23 bit_66_23 gnd C_bl
Cbb_66_23 bitb_66_23 gnd C_bl
Rb_66_24 bit_66_24 bit_66_25 R_bl
Rbb_66_24 bitb_66_24 bitb_66_25 R_bl
Cb_66_24 bit_66_24 gnd C_bl
Cbb_66_24 bitb_66_24 gnd C_bl
Rb_66_25 bit_66_25 bit_66_26 R_bl
Rbb_66_25 bitb_66_25 bitb_66_26 R_bl
Cb_66_25 bit_66_25 gnd C_bl
Cbb_66_25 bitb_66_25 gnd C_bl
Rb_66_26 bit_66_26 bit_66_27 R_bl
Rbb_66_26 bitb_66_26 bitb_66_27 R_bl
Cb_66_26 bit_66_26 gnd C_bl
Cbb_66_26 bitb_66_26 gnd C_bl
Rb_66_27 bit_66_27 bit_66_28 R_bl
Rbb_66_27 bitb_66_27 bitb_66_28 R_bl
Cb_66_27 bit_66_27 gnd C_bl
Cbb_66_27 bitb_66_27 gnd C_bl
Rb_66_28 bit_66_28 bit_66_29 R_bl
Rbb_66_28 bitb_66_28 bitb_66_29 R_bl
Cb_66_28 bit_66_28 gnd C_bl
Cbb_66_28 bitb_66_28 gnd C_bl
Rb_66_29 bit_66_29 bit_66_30 R_bl
Rbb_66_29 bitb_66_29 bitb_66_30 R_bl
Cb_66_29 bit_66_29 gnd C_bl
Cbb_66_29 bitb_66_29 gnd C_bl
Rb_66_30 bit_66_30 bit_66_31 R_bl
Rbb_66_30 bitb_66_30 bitb_66_31 R_bl
Cb_66_30 bit_66_30 gnd C_bl
Cbb_66_30 bitb_66_30 gnd C_bl
Rb_66_31 bit_66_31 bit_66_32 R_bl
Rbb_66_31 bitb_66_31 bitb_66_32 R_bl
Cb_66_31 bit_66_31 gnd C_bl
Cbb_66_31 bitb_66_31 gnd C_bl
Rb_66_32 bit_66_32 bit_66_33 R_bl
Rbb_66_32 bitb_66_32 bitb_66_33 R_bl
Cb_66_32 bit_66_32 gnd C_bl
Cbb_66_32 bitb_66_32 gnd C_bl
Rb_66_33 bit_66_33 bit_66_34 R_bl
Rbb_66_33 bitb_66_33 bitb_66_34 R_bl
Cb_66_33 bit_66_33 gnd C_bl
Cbb_66_33 bitb_66_33 gnd C_bl
Rb_66_34 bit_66_34 bit_66_35 R_bl
Rbb_66_34 bitb_66_34 bitb_66_35 R_bl
Cb_66_34 bit_66_34 gnd C_bl
Cbb_66_34 bitb_66_34 gnd C_bl
Rb_66_35 bit_66_35 bit_66_36 R_bl
Rbb_66_35 bitb_66_35 bitb_66_36 R_bl
Cb_66_35 bit_66_35 gnd C_bl
Cbb_66_35 bitb_66_35 gnd C_bl
Rb_66_36 bit_66_36 bit_66_37 R_bl
Rbb_66_36 bitb_66_36 bitb_66_37 R_bl
Cb_66_36 bit_66_36 gnd C_bl
Cbb_66_36 bitb_66_36 gnd C_bl
Rb_66_37 bit_66_37 bit_66_38 R_bl
Rbb_66_37 bitb_66_37 bitb_66_38 R_bl
Cb_66_37 bit_66_37 gnd C_bl
Cbb_66_37 bitb_66_37 gnd C_bl
Rb_66_38 bit_66_38 bit_66_39 R_bl
Rbb_66_38 bitb_66_38 bitb_66_39 R_bl
Cb_66_38 bit_66_38 gnd C_bl
Cbb_66_38 bitb_66_38 gnd C_bl
Rb_66_39 bit_66_39 bit_66_40 R_bl
Rbb_66_39 bitb_66_39 bitb_66_40 R_bl
Cb_66_39 bit_66_39 gnd C_bl
Cbb_66_39 bitb_66_39 gnd C_bl
Rb_66_40 bit_66_40 bit_66_41 R_bl
Rbb_66_40 bitb_66_40 bitb_66_41 R_bl
Cb_66_40 bit_66_40 gnd C_bl
Cbb_66_40 bitb_66_40 gnd C_bl
Rb_66_41 bit_66_41 bit_66_42 R_bl
Rbb_66_41 bitb_66_41 bitb_66_42 R_bl
Cb_66_41 bit_66_41 gnd C_bl
Cbb_66_41 bitb_66_41 gnd C_bl
Rb_66_42 bit_66_42 bit_66_43 R_bl
Rbb_66_42 bitb_66_42 bitb_66_43 R_bl
Cb_66_42 bit_66_42 gnd C_bl
Cbb_66_42 bitb_66_42 gnd C_bl
Rb_66_43 bit_66_43 bit_66_44 R_bl
Rbb_66_43 bitb_66_43 bitb_66_44 R_bl
Cb_66_43 bit_66_43 gnd C_bl
Cbb_66_43 bitb_66_43 gnd C_bl
Rb_66_44 bit_66_44 bit_66_45 R_bl
Rbb_66_44 bitb_66_44 bitb_66_45 R_bl
Cb_66_44 bit_66_44 gnd C_bl
Cbb_66_44 bitb_66_44 gnd C_bl
Rb_66_45 bit_66_45 bit_66_46 R_bl
Rbb_66_45 bitb_66_45 bitb_66_46 R_bl
Cb_66_45 bit_66_45 gnd C_bl
Cbb_66_45 bitb_66_45 gnd C_bl
Rb_66_46 bit_66_46 bit_66_47 R_bl
Rbb_66_46 bitb_66_46 bitb_66_47 R_bl
Cb_66_46 bit_66_46 gnd C_bl
Cbb_66_46 bitb_66_46 gnd C_bl
Rb_66_47 bit_66_47 bit_66_48 R_bl
Rbb_66_47 bitb_66_47 bitb_66_48 R_bl
Cb_66_47 bit_66_47 gnd C_bl
Cbb_66_47 bitb_66_47 gnd C_bl
Rb_66_48 bit_66_48 bit_66_49 R_bl
Rbb_66_48 bitb_66_48 bitb_66_49 R_bl
Cb_66_48 bit_66_48 gnd C_bl
Cbb_66_48 bitb_66_48 gnd C_bl
Rb_66_49 bit_66_49 bit_66_50 R_bl
Rbb_66_49 bitb_66_49 bitb_66_50 R_bl
Cb_66_49 bit_66_49 gnd C_bl
Cbb_66_49 bitb_66_49 gnd C_bl
Rb_66_50 bit_66_50 bit_66_51 R_bl
Rbb_66_50 bitb_66_50 bitb_66_51 R_bl
Cb_66_50 bit_66_50 gnd C_bl
Cbb_66_50 bitb_66_50 gnd C_bl
Rb_66_51 bit_66_51 bit_66_52 R_bl
Rbb_66_51 bitb_66_51 bitb_66_52 R_bl
Cb_66_51 bit_66_51 gnd C_bl
Cbb_66_51 bitb_66_51 gnd C_bl
Rb_66_52 bit_66_52 bit_66_53 R_bl
Rbb_66_52 bitb_66_52 bitb_66_53 R_bl
Cb_66_52 bit_66_52 gnd C_bl
Cbb_66_52 bitb_66_52 gnd C_bl
Rb_66_53 bit_66_53 bit_66_54 R_bl
Rbb_66_53 bitb_66_53 bitb_66_54 R_bl
Cb_66_53 bit_66_53 gnd C_bl
Cbb_66_53 bitb_66_53 gnd C_bl
Rb_66_54 bit_66_54 bit_66_55 R_bl
Rbb_66_54 bitb_66_54 bitb_66_55 R_bl
Cb_66_54 bit_66_54 gnd C_bl
Cbb_66_54 bitb_66_54 gnd C_bl
Rb_66_55 bit_66_55 bit_66_56 R_bl
Rbb_66_55 bitb_66_55 bitb_66_56 R_bl
Cb_66_55 bit_66_55 gnd C_bl
Cbb_66_55 bitb_66_55 gnd C_bl
Rb_66_56 bit_66_56 bit_66_57 R_bl
Rbb_66_56 bitb_66_56 bitb_66_57 R_bl
Cb_66_56 bit_66_56 gnd C_bl
Cbb_66_56 bitb_66_56 gnd C_bl
Rb_66_57 bit_66_57 bit_66_58 R_bl
Rbb_66_57 bitb_66_57 bitb_66_58 R_bl
Cb_66_57 bit_66_57 gnd C_bl
Cbb_66_57 bitb_66_57 gnd C_bl
Rb_66_58 bit_66_58 bit_66_59 R_bl
Rbb_66_58 bitb_66_58 bitb_66_59 R_bl
Cb_66_58 bit_66_58 gnd C_bl
Cbb_66_58 bitb_66_58 gnd C_bl
Rb_66_59 bit_66_59 bit_66_60 R_bl
Rbb_66_59 bitb_66_59 bitb_66_60 R_bl
Cb_66_59 bit_66_59 gnd C_bl
Cbb_66_59 bitb_66_59 gnd C_bl
Rb_66_60 bit_66_60 bit_66_61 R_bl
Rbb_66_60 bitb_66_60 bitb_66_61 R_bl
Cb_66_60 bit_66_60 gnd C_bl
Cbb_66_60 bitb_66_60 gnd C_bl
Rb_66_61 bit_66_61 bit_66_62 R_bl
Rbb_66_61 bitb_66_61 bitb_66_62 R_bl
Cb_66_61 bit_66_61 gnd C_bl
Cbb_66_61 bitb_66_61 gnd C_bl
Rb_66_62 bit_66_62 bit_66_63 R_bl
Rbb_66_62 bitb_66_62 bitb_66_63 R_bl
Cb_66_62 bit_66_62 gnd C_bl
Cbb_66_62 bitb_66_62 gnd C_bl
Rb_66_63 bit_66_63 bit_66_64 R_bl
Rbb_66_63 bitb_66_63 bitb_66_64 R_bl
Cb_66_63 bit_66_63 gnd C_bl
Cbb_66_63 bitb_66_63 gnd C_bl
Rb_66_64 bit_66_64 bit_66_65 R_bl
Rbb_66_64 bitb_66_64 bitb_66_65 R_bl
Cb_66_64 bit_66_64 gnd C_bl
Cbb_66_64 bitb_66_64 gnd C_bl
Rb_66_65 bit_66_65 bit_66_66 R_bl
Rbb_66_65 bitb_66_65 bitb_66_66 R_bl
Cb_66_65 bit_66_65 gnd C_bl
Cbb_66_65 bitb_66_65 gnd C_bl
Rb_66_66 bit_66_66 bit_66_67 R_bl
Rbb_66_66 bitb_66_66 bitb_66_67 R_bl
Cb_66_66 bit_66_66 gnd C_bl
Cbb_66_66 bitb_66_66 gnd C_bl
Rb_66_67 bit_66_67 bit_66_68 R_bl
Rbb_66_67 bitb_66_67 bitb_66_68 R_bl
Cb_66_67 bit_66_67 gnd C_bl
Cbb_66_67 bitb_66_67 gnd C_bl
Rb_66_68 bit_66_68 bit_66_69 R_bl
Rbb_66_68 bitb_66_68 bitb_66_69 R_bl
Cb_66_68 bit_66_68 gnd C_bl
Cbb_66_68 bitb_66_68 gnd C_bl
Rb_66_69 bit_66_69 bit_66_70 R_bl
Rbb_66_69 bitb_66_69 bitb_66_70 R_bl
Cb_66_69 bit_66_69 gnd C_bl
Cbb_66_69 bitb_66_69 gnd C_bl
Rb_66_70 bit_66_70 bit_66_71 R_bl
Rbb_66_70 bitb_66_70 bitb_66_71 R_bl
Cb_66_70 bit_66_70 gnd C_bl
Cbb_66_70 bitb_66_70 gnd C_bl
Rb_66_71 bit_66_71 bit_66_72 R_bl
Rbb_66_71 bitb_66_71 bitb_66_72 R_bl
Cb_66_71 bit_66_71 gnd C_bl
Cbb_66_71 bitb_66_71 gnd C_bl
Rb_66_72 bit_66_72 bit_66_73 R_bl
Rbb_66_72 bitb_66_72 bitb_66_73 R_bl
Cb_66_72 bit_66_72 gnd C_bl
Cbb_66_72 bitb_66_72 gnd C_bl
Rb_66_73 bit_66_73 bit_66_74 R_bl
Rbb_66_73 bitb_66_73 bitb_66_74 R_bl
Cb_66_73 bit_66_73 gnd C_bl
Cbb_66_73 bitb_66_73 gnd C_bl
Rb_66_74 bit_66_74 bit_66_75 R_bl
Rbb_66_74 bitb_66_74 bitb_66_75 R_bl
Cb_66_74 bit_66_74 gnd C_bl
Cbb_66_74 bitb_66_74 gnd C_bl
Rb_66_75 bit_66_75 bit_66_76 R_bl
Rbb_66_75 bitb_66_75 bitb_66_76 R_bl
Cb_66_75 bit_66_75 gnd C_bl
Cbb_66_75 bitb_66_75 gnd C_bl
Rb_66_76 bit_66_76 bit_66_77 R_bl
Rbb_66_76 bitb_66_76 bitb_66_77 R_bl
Cb_66_76 bit_66_76 gnd C_bl
Cbb_66_76 bitb_66_76 gnd C_bl
Rb_66_77 bit_66_77 bit_66_78 R_bl
Rbb_66_77 bitb_66_77 bitb_66_78 R_bl
Cb_66_77 bit_66_77 gnd C_bl
Cbb_66_77 bitb_66_77 gnd C_bl
Rb_66_78 bit_66_78 bit_66_79 R_bl
Rbb_66_78 bitb_66_78 bitb_66_79 R_bl
Cb_66_78 bit_66_78 gnd C_bl
Cbb_66_78 bitb_66_78 gnd C_bl
Rb_66_79 bit_66_79 bit_66_80 R_bl
Rbb_66_79 bitb_66_79 bitb_66_80 R_bl
Cb_66_79 bit_66_79 gnd C_bl
Cbb_66_79 bitb_66_79 gnd C_bl
Rb_66_80 bit_66_80 bit_66_81 R_bl
Rbb_66_80 bitb_66_80 bitb_66_81 R_bl
Cb_66_80 bit_66_80 gnd C_bl
Cbb_66_80 bitb_66_80 gnd C_bl
Rb_66_81 bit_66_81 bit_66_82 R_bl
Rbb_66_81 bitb_66_81 bitb_66_82 R_bl
Cb_66_81 bit_66_81 gnd C_bl
Cbb_66_81 bitb_66_81 gnd C_bl
Rb_66_82 bit_66_82 bit_66_83 R_bl
Rbb_66_82 bitb_66_82 bitb_66_83 R_bl
Cb_66_82 bit_66_82 gnd C_bl
Cbb_66_82 bitb_66_82 gnd C_bl
Rb_66_83 bit_66_83 bit_66_84 R_bl
Rbb_66_83 bitb_66_83 bitb_66_84 R_bl
Cb_66_83 bit_66_83 gnd C_bl
Cbb_66_83 bitb_66_83 gnd C_bl
Rb_66_84 bit_66_84 bit_66_85 R_bl
Rbb_66_84 bitb_66_84 bitb_66_85 R_bl
Cb_66_84 bit_66_84 gnd C_bl
Cbb_66_84 bitb_66_84 gnd C_bl
Rb_66_85 bit_66_85 bit_66_86 R_bl
Rbb_66_85 bitb_66_85 bitb_66_86 R_bl
Cb_66_85 bit_66_85 gnd C_bl
Cbb_66_85 bitb_66_85 gnd C_bl
Rb_66_86 bit_66_86 bit_66_87 R_bl
Rbb_66_86 bitb_66_86 bitb_66_87 R_bl
Cb_66_86 bit_66_86 gnd C_bl
Cbb_66_86 bitb_66_86 gnd C_bl
Rb_66_87 bit_66_87 bit_66_88 R_bl
Rbb_66_87 bitb_66_87 bitb_66_88 R_bl
Cb_66_87 bit_66_87 gnd C_bl
Cbb_66_87 bitb_66_87 gnd C_bl
Rb_66_88 bit_66_88 bit_66_89 R_bl
Rbb_66_88 bitb_66_88 bitb_66_89 R_bl
Cb_66_88 bit_66_88 gnd C_bl
Cbb_66_88 bitb_66_88 gnd C_bl
Rb_66_89 bit_66_89 bit_66_90 R_bl
Rbb_66_89 bitb_66_89 bitb_66_90 R_bl
Cb_66_89 bit_66_89 gnd C_bl
Cbb_66_89 bitb_66_89 gnd C_bl
Rb_66_90 bit_66_90 bit_66_91 R_bl
Rbb_66_90 bitb_66_90 bitb_66_91 R_bl
Cb_66_90 bit_66_90 gnd C_bl
Cbb_66_90 bitb_66_90 gnd C_bl
Rb_66_91 bit_66_91 bit_66_92 R_bl
Rbb_66_91 bitb_66_91 bitb_66_92 R_bl
Cb_66_91 bit_66_91 gnd C_bl
Cbb_66_91 bitb_66_91 gnd C_bl
Rb_66_92 bit_66_92 bit_66_93 R_bl
Rbb_66_92 bitb_66_92 bitb_66_93 R_bl
Cb_66_92 bit_66_92 gnd C_bl
Cbb_66_92 bitb_66_92 gnd C_bl
Rb_66_93 bit_66_93 bit_66_94 R_bl
Rbb_66_93 bitb_66_93 bitb_66_94 R_bl
Cb_66_93 bit_66_93 gnd C_bl
Cbb_66_93 bitb_66_93 gnd C_bl
Rb_66_94 bit_66_94 bit_66_95 R_bl
Rbb_66_94 bitb_66_94 bitb_66_95 R_bl
Cb_66_94 bit_66_94 gnd C_bl
Cbb_66_94 bitb_66_94 gnd C_bl
Rb_66_95 bit_66_95 bit_66_96 R_bl
Rbb_66_95 bitb_66_95 bitb_66_96 R_bl
Cb_66_95 bit_66_95 gnd C_bl
Cbb_66_95 bitb_66_95 gnd C_bl
Rb_66_96 bit_66_96 bit_66_97 R_bl
Rbb_66_96 bitb_66_96 bitb_66_97 R_bl
Cb_66_96 bit_66_96 gnd C_bl
Cbb_66_96 bitb_66_96 gnd C_bl
Rb_66_97 bit_66_97 bit_66_98 R_bl
Rbb_66_97 bitb_66_97 bitb_66_98 R_bl
Cb_66_97 bit_66_97 gnd C_bl
Cbb_66_97 bitb_66_97 gnd C_bl
Rb_66_98 bit_66_98 bit_66_99 R_bl
Rbb_66_98 bitb_66_98 bitb_66_99 R_bl
Cb_66_98 bit_66_98 gnd C_bl
Cbb_66_98 bitb_66_98 gnd C_bl
Rb_66_99 bit_66_99 bit_66_100 R_bl
Rbb_66_99 bitb_66_99 bitb_66_100 R_bl
Cb_66_99 bit_66_99 gnd C_bl
Cbb_66_99 bitb_66_99 gnd C_bl
Rb_67_0 bit_67_0 bit_67_1 R_bl
Rbb_67_0 bitb_67_0 bitb_67_1 R_bl
Cb_67_0 bit_67_0 gnd C_bl
Cbb_67_0 bitb_67_0 gnd C_bl
Rb_67_1 bit_67_1 bit_67_2 R_bl
Rbb_67_1 bitb_67_1 bitb_67_2 R_bl
Cb_67_1 bit_67_1 gnd C_bl
Cbb_67_1 bitb_67_1 gnd C_bl
Rb_67_2 bit_67_2 bit_67_3 R_bl
Rbb_67_2 bitb_67_2 bitb_67_3 R_bl
Cb_67_2 bit_67_2 gnd C_bl
Cbb_67_2 bitb_67_2 gnd C_bl
Rb_67_3 bit_67_3 bit_67_4 R_bl
Rbb_67_3 bitb_67_3 bitb_67_4 R_bl
Cb_67_3 bit_67_3 gnd C_bl
Cbb_67_3 bitb_67_3 gnd C_bl
Rb_67_4 bit_67_4 bit_67_5 R_bl
Rbb_67_4 bitb_67_4 bitb_67_5 R_bl
Cb_67_4 bit_67_4 gnd C_bl
Cbb_67_4 bitb_67_4 gnd C_bl
Rb_67_5 bit_67_5 bit_67_6 R_bl
Rbb_67_5 bitb_67_5 bitb_67_6 R_bl
Cb_67_5 bit_67_5 gnd C_bl
Cbb_67_5 bitb_67_5 gnd C_bl
Rb_67_6 bit_67_6 bit_67_7 R_bl
Rbb_67_6 bitb_67_6 bitb_67_7 R_bl
Cb_67_6 bit_67_6 gnd C_bl
Cbb_67_6 bitb_67_6 gnd C_bl
Rb_67_7 bit_67_7 bit_67_8 R_bl
Rbb_67_7 bitb_67_7 bitb_67_8 R_bl
Cb_67_7 bit_67_7 gnd C_bl
Cbb_67_7 bitb_67_7 gnd C_bl
Rb_67_8 bit_67_8 bit_67_9 R_bl
Rbb_67_8 bitb_67_8 bitb_67_9 R_bl
Cb_67_8 bit_67_8 gnd C_bl
Cbb_67_8 bitb_67_8 gnd C_bl
Rb_67_9 bit_67_9 bit_67_10 R_bl
Rbb_67_9 bitb_67_9 bitb_67_10 R_bl
Cb_67_9 bit_67_9 gnd C_bl
Cbb_67_9 bitb_67_9 gnd C_bl
Rb_67_10 bit_67_10 bit_67_11 R_bl
Rbb_67_10 bitb_67_10 bitb_67_11 R_bl
Cb_67_10 bit_67_10 gnd C_bl
Cbb_67_10 bitb_67_10 gnd C_bl
Rb_67_11 bit_67_11 bit_67_12 R_bl
Rbb_67_11 bitb_67_11 bitb_67_12 R_bl
Cb_67_11 bit_67_11 gnd C_bl
Cbb_67_11 bitb_67_11 gnd C_bl
Rb_67_12 bit_67_12 bit_67_13 R_bl
Rbb_67_12 bitb_67_12 bitb_67_13 R_bl
Cb_67_12 bit_67_12 gnd C_bl
Cbb_67_12 bitb_67_12 gnd C_bl
Rb_67_13 bit_67_13 bit_67_14 R_bl
Rbb_67_13 bitb_67_13 bitb_67_14 R_bl
Cb_67_13 bit_67_13 gnd C_bl
Cbb_67_13 bitb_67_13 gnd C_bl
Rb_67_14 bit_67_14 bit_67_15 R_bl
Rbb_67_14 bitb_67_14 bitb_67_15 R_bl
Cb_67_14 bit_67_14 gnd C_bl
Cbb_67_14 bitb_67_14 gnd C_bl
Rb_67_15 bit_67_15 bit_67_16 R_bl
Rbb_67_15 bitb_67_15 bitb_67_16 R_bl
Cb_67_15 bit_67_15 gnd C_bl
Cbb_67_15 bitb_67_15 gnd C_bl
Rb_67_16 bit_67_16 bit_67_17 R_bl
Rbb_67_16 bitb_67_16 bitb_67_17 R_bl
Cb_67_16 bit_67_16 gnd C_bl
Cbb_67_16 bitb_67_16 gnd C_bl
Rb_67_17 bit_67_17 bit_67_18 R_bl
Rbb_67_17 bitb_67_17 bitb_67_18 R_bl
Cb_67_17 bit_67_17 gnd C_bl
Cbb_67_17 bitb_67_17 gnd C_bl
Rb_67_18 bit_67_18 bit_67_19 R_bl
Rbb_67_18 bitb_67_18 bitb_67_19 R_bl
Cb_67_18 bit_67_18 gnd C_bl
Cbb_67_18 bitb_67_18 gnd C_bl
Rb_67_19 bit_67_19 bit_67_20 R_bl
Rbb_67_19 bitb_67_19 bitb_67_20 R_bl
Cb_67_19 bit_67_19 gnd C_bl
Cbb_67_19 bitb_67_19 gnd C_bl
Rb_67_20 bit_67_20 bit_67_21 R_bl
Rbb_67_20 bitb_67_20 bitb_67_21 R_bl
Cb_67_20 bit_67_20 gnd C_bl
Cbb_67_20 bitb_67_20 gnd C_bl
Rb_67_21 bit_67_21 bit_67_22 R_bl
Rbb_67_21 bitb_67_21 bitb_67_22 R_bl
Cb_67_21 bit_67_21 gnd C_bl
Cbb_67_21 bitb_67_21 gnd C_bl
Rb_67_22 bit_67_22 bit_67_23 R_bl
Rbb_67_22 bitb_67_22 bitb_67_23 R_bl
Cb_67_22 bit_67_22 gnd C_bl
Cbb_67_22 bitb_67_22 gnd C_bl
Rb_67_23 bit_67_23 bit_67_24 R_bl
Rbb_67_23 bitb_67_23 bitb_67_24 R_bl
Cb_67_23 bit_67_23 gnd C_bl
Cbb_67_23 bitb_67_23 gnd C_bl
Rb_67_24 bit_67_24 bit_67_25 R_bl
Rbb_67_24 bitb_67_24 bitb_67_25 R_bl
Cb_67_24 bit_67_24 gnd C_bl
Cbb_67_24 bitb_67_24 gnd C_bl
Rb_67_25 bit_67_25 bit_67_26 R_bl
Rbb_67_25 bitb_67_25 bitb_67_26 R_bl
Cb_67_25 bit_67_25 gnd C_bl
Cbb_67_25 bitb_67_25 gnd C_bl
Rb_67_26 bit_67_26 bit_67_27 R_bl
Rbb_67_26 bitb_67_26 bitb_67_27 R_bl
Cb_67_26 bit_67_26 gnd C_bl
Cbb_67_26 bitb_67_26 gnd C_bl
Rb_67_27 bit_67_27 bit_67_28 R_bl
Rbb_67_27 bitb_67_27 bitb_67_28 R_bl
Cb_67_27 bit_67_27 gnd C_bl
Cbb_67_27 bitb_67_27 gnd C_bl
Rb_67_28 bit_67_28 bit_67_29 R_bl
Rbb_67_28 bitb_67_28 bitb_67_29 R_bl
Cb_67_28 bit_67_28 gnd C_bl
Cbb_67_28 bitb_67_28 gnd C_bl
Rb_67_29 bit_67_29 bit_67_30 R_bl
Rbb_67_29 bitb_67_29 bitb_67_30 R_bl
Cb_67_29 bit_67_29 gnd C_bl
Cbb_67_29 bitb_67_29 gnd C_bl
Rb_67_30 bit_67_30 bit_67_31 R_bl
Rbb_67_30 bitb_67_30 bitb_67_31 R_bl
Cb_67_30 bit_67_30 gnd C_bl
Cbb_67_30 bitb_67_30 gnd C_bl
Rb_67_31 bit_67_31 bit_67_32 R_bl
Rbb_67_31 bitb_67_31 bitb_67_32 R_bl
Cb_67_31 bit_67_31 gnd C_bl
Cbb_67_31 bitb_67_31 gnd C_bl
Rb_67_32 bit_67_32 bit_67_33 R_bl
Rbb_67_32 bitb_67_32 bitb_67_33 R_bl
Cb_67_32 bit_67_32 gnd C_bl
Cbb_67_32 bitb_67_32 gnd C_bl
Rb_67_33 bit_67_33 bit_67_34 R_bl
Rbb_67_33 bitb_67_33 bitb_67_34 R_bl
Cb_67_33 bit_67_33 gnd C_bl
Cbb_67_33 bitb_67_33 gnd C_bl
Rb_67_34 bit_67_34 bit_67_35 R_bl
Rbb_67_34 bitb_67_34 bitb_67_35 R_bl
Cb_67_34 bit_67_34 gnd C_bl
Cbb_67_34 bitb_67_34 gnd C_bl
Rb_67_35 bit_67_35 bit_67_36 R_bl
Rbb_67_35 bitb_67_35 bitb_67_36 R_bl
Cb_67_35 bit_67_35 gnd C_bl
Cbb_67_35 bitb_67_35 gnd C_bl
Rb_67_36 bit_67_36 bit_67_37 R_bl
Rbb_67_36 bitb_67_36 bitb_67_37 R_bl
Cb_67_36 bit_67_36 gnd C_bl
Cbb_67_36 bitb_67_36 gnd C_bl
Rb_67_37 bit_67_37 bit_67_38 R_bl
Rbb_67_37 bitb_67_37 bitb_67_38 R_bl
Cb_67_37 bit_67_37 gnd C_bl
Cbb_67_37 bitb_67_37 gnd C_bl
Rb_67_38 bit_67_38 bit_67_39 R_bl
Rbb_67_38 bitb_67_38 bitb_67_39 R_bl
Cb_67_38 bit_67_38 gnd C_bl
Cbb_67_38 bitb_67_38 gnd C_bl
Rb_67_39 bit_67_39 bit_67_40 R_bl
Rbb_67_39 bitb_67_39 bitb_67_40 R_bl
Cb_67_39 bit_67_39 gnd C_bl
Cbb_67_39 bitb_67_39 gnd C_bl
Rb_67_40 bit_67_40 bit_67_41 R_bl
Rbb_67_40 bitb_67_40 bitb_67_41 R_bl
Cb_67_40 bit_67_40 gnd C_bl
Cbb_67_40 bitb_67_40 gnd C_bl
Rb_67_41 bit_67_41 bit_67_42 R_bl
Rbb_67_41 bitb_67_41 bitb_67_42 R_bl
Cb_67_41 bit_67_41 gnd C_bl
Cbb_67_41 bitb_67_41 gnd C_bl
Rb_67_42 bit_67_42 bit_67_43 R_bl
Rbb_67_42 bitb_67_42 bitb_67_43 R_bl
Cb_67_42 bit_67_42 gnd C_bl
Cbb_67_42 bitb_67_42 gnd C_bl
Rb_67_43 bit_67_43 bit_67_44 R_bl
Rbb_67_43 bitb_67_43 bitb_67_44 R_bl
Cb_67_43 bit_67_43 gnd C_bl
Cbb_67_43 bitb_67_43 gnd C_bl
Rb_67_44 bit_67_44 bit_67_45 R_bl
Rbb_67_44 bitb_67_44 bitb_67_45 R_bl
Cb_67_44 bit_67_44 gnd C_bl
Cbb_67_44 bitb_67_44 gnd C_bl
Rb_67_45 bit_67_45 bit_67_46 R_bl
Rbb_67_45 bitb_67_45 bitb_67_46 R_bl
Cb_67_45 bit_67_45 gnd C_bl
Cbb_67_45 bitb_67_45 gnd C_bl
Rb_67_46 bit_67_46 bit_67_47 R_bl
Rbb_67_46 bitb_67_46 bitb_67_47 R_bl
Cb_67_46 bit_67_46 gnd C_bl
Cbb_67_46 bitb_67_46 gnd C_bl
Rb_67_47 bit_67_47 bit_67_48 R_bl
Rbb_67_47 bitb_67_47 bitb_67_48 R_bl
Cb_67_47 bit_67_47 gnd C_bl
Cbb_67_47 bitb_67_47 gnd C_bl
Rb_67_48 bit_67_48 bit_67_49 R_bl
Rbb_67_48 bitb_67_48 bitb_67_49 R_bl
Cb_67_48 bit_67_48 gnd C_bl
Cbb_67_48 bitb_67_48 gnd C_bl
Rb_67_49 bit_67_49 bit_67_50 R_bl
Rbb_67_49 bitb_67_49 bitb_67_50 R_bl
Cb_67_49 bit_67_49 gnd C_bl
Cbb_67_49 bitb_67_49 gnd C_bl
Rb_67_50 bit_67_50 bit_67_51 R_bl
Rbb_67_50 bitb_67_50 bitb_67_51 R_bl
Cb_67_50 bit_67_50 gnd C_bl
Cbb_67_50 bitb_67_50 gnd C_bl
Rb_67_51 bit_67_51 bit_67_52 R_bl
Rbb_67_51 bitb_67_51 bitb_67_52 R_bl
Cb_67_51 bit_67_51 gnd C_bl
Cbb_67_51 bitb_67_51 gnd C_bl
Rb_67_52 bit_67_52 bit_67_53 R_bl
Rbb_67_52 bitb_67_52 bitb_67_53 R_bl
Cb_67_52 bit_67_52 gnd C_bl
Cbb_67_52 bitb_67_52 gnd C_bl
Rb_67_53 bit_67_53 bit_67_54 R_bl
Rbb_67_53 bitb_67_53 bitb_67_54 R_bl
Cb_67_53 bit_67_53 gnd C_bl
Cbb_67_53 bitb_67_53 gnd C_bl
Rb_67_54 bit_67_54 bit_67_55 R_bl
Rbb_67_54 bitb_67_54 bitb_67_55 R_bl
Cb_67_54 bit_67_54 gnd C_bl
Cbb_67_54 bitb_67_54 gnd C_bl
Rb_67_55 bit_67_55 bit_67_56 R_bl
Rbb_67_55 bitb_67_55 bitb_67_56 R_bl
Cb_67_55 bit_67_55 gnd C_bl
Cbb_67_55 bitb_67_55 gnd C_bl
Rb_67_56 bit_67_56 bit_67_57 R_bl
Rbb_67_56 bitb_67_56 bitb_67_57 R_bl
Cb_67_56 bit_67_56 gnd C_bl
Cbb_67_56 bitb_67_56 gnd C_bl
Rb_67_57 bit_67_57 bit_67_58 R_bl
Rbb_67_57 bitb_67_57 bitb_67_58 R_bl
Cb_67_57 bit_67_57 gnd C_bl
Cbb_67_57 bitb_67_57 gnd C_bl
Rb_67_58 bit_67_58 bit_67_59 R_bl
Rbb_67_58 bitb_67_58 bitb_67_59 R_bl
Cb_67_58 bit_67_58 gnd C_bl
Cbb_67_58 bitb_67_58 gnd C_bl
Rb_67_59 bit_67_59 bit_67_60 R_bl
Rbb_67_59 bitb_67_59 bitb_67_60 R_bl
Cb_67_59 bit_67_59 gnd C_bl
Cbb_67_59 bitb_67_59 gnd C_bl
Rb_67_60 bit_67_60 bit_67_61 R_bl
Rbb_67_60 bitb_67_60 bitb_67_61 R_bl
Cb_67_60 bit_67_60 gnd C_bl
Cbb_67_60 bitb_67_60 gnd C_bl
Rb_67_61 bit_67_61 bit_67_62 R_bl
Rbb_67_61 bitb_67_61 bitb_67_62 R_bl
Cb_67_61 bit_67_61 gnd C_bl
Cbb_67_61 bitb_67_61 gnd C_bl
Rb_67_62 bit_67_62 bit_67_63 R_bl
Rbb_67_62 bitb_67_62 bitb_67_63 R_bl
Cb_67_62 bit_67_62 gnd C_bl
Cbb_67_62 bitb_67_62 gnd C_bl
Rb_67_63 bit_67_63 bit_67_64 R_bl
Rbb_67_63 bitb_67_63 bitb_67_64 R_bl
Cb_67_63 bit_67_63 gnd C_bl
Cbb_67_63 bitb_67_63 gnd C_bl
Rb_67_64 bit_67_64 bit_67_65 R_bl
Rbb_67_64 bitb_67_64 bitb_67_65 R_bl
Cb_67_64 bit_67_64 gnd C_bl
Cbb_67_64 bitb_67_64 gnd C_bl
Rb_67_65 bit_67_65 bit_67_66 R_bl
Rbb_67_65 bitb_67_65 bitb_67_66 R_bl
Cb_67_65 bit_67_65 gnd C_bl
Cbb_67_65 bitb_67_65 gnd C_bl
Rb_67_66 bit_67_66 bit_67_67 R_bl
Rbb_67_66 bitb_67_66 bitb_67_67 R_bl
Cb_67_66 bit_67_66 gnd C_bl
Cbb_67_66 bitb_67_66 gnd C_bl
Rb_67_67 bit_67_67 bit_67_68 R_bl
Rbb_67_67 bitb_67_67 bitb_67_68 R_bl
Cb_67_67 bit_67_67 gnd C_bl
Cbb_67_67 bitb_67_67 gnd C_bl
Rb_67_68 bit_67_68 bit_67_69 R_bl
Rbb_67_68 bitb_67_68 bitb_67_69 R_bl
Cb_67_68 bit_67_68 gnd C_bl
Cbb_67_68 bitb_67_68 gnd C_bl
Rb_67_69 bit_67_69 bit_67_70 R_bl
Rbb_67_69 bitb_67_69 bitb_67_70 R_bl
Cb_67_69 bit_67_69 gnd C_bl
Cbb_67_69 bitb_67_69 gnd C_bl
Rb_67_70 bit_67_70 bit_67_71 R_bl
Rbb_67_70 bitb_67_70 bitb_67_71 R_bl
Cb_67_70 bit_67_70 gnd C_bl
Cbb_67_70 bitb_67_70 gnd C_bl
Rb_67_71 bit_67_71 bit_67_72 R_bl
Rbb_67_71 bitb_67_71 bitb_67_72 R_bl
Cb_67_71 bit_67_71 gnd C_bl
Cbb_67_71 bitb_67_71 gnd C_bl
Rb_67_72 bit_67_72 bit_67_73 R_bl
Rbb_67_72 bitb_67_72 bitb_67_73 R_bl
Cb_67_72 bit_67_72 gnd C_bl
Cbb_67_72 bitb_67_72 gnd C_bl
Rb_67_73 bit_67_73 bit_67_74 R_bl
Rbb_67_73 bitb_67_73 bitb_67_74 R_bl
Cb_67_73 bit_67_73 gnd C_bl
Cbb_67_73 bitb_67_73 gnd C_bl
Rb_67_74 bit_67_74 bit_67_75 R_bl
Rbb_67_74 bitb_67_74 bitb_67_75 R_bl
Cb_67_74 bit_67_74 gnd C_bl
Cbb_67_74 bitb_67_74 gnd C_bl
Rb_67_75 bit_67_75 bit_67_76 R_bl
Rbb_67_75 bitb_67_75 bitb_67_76 R_bl
Cb_67_75 bit_67_75 gnd C_bl
Cbb_67_75 bitb_67_75 gnd C_bl
Rb_67_76 bit_67_76 bit_67_77 R_bl
Rbb_67_76 bitb_67_76 bitb_67_77 R_bl
Cb_67_76 bit_67_76 gnd C_bl
Cbb_67_76 bitb_67_76 gnd C_bl
Rb_67_77 bit_67_77 bit_67_78 R_bl
Rbb_67_77 bitb_67_77 bitb_67_78 R_bl
Cb_67_77 bit_67_77 gnd C_bl
Cbb_67_77 bitb_67_77 gnd C_bl
Rb_67_78 bit_67_78 bit_67_79 R_bl
Rbb_67_78 bitb_67_78 bitb_67_79 R_bl
Cb_67_78 bit_67_78 gnd C_bl
Cbb_67_78 bitb_67_78 gnd C_bl
Rb_67_79 bit_67_79 bit_67_80 R_bl
Rbb_67_79 bitb_67_79 bitb_67_80 R_bl
Cb_67_79 bit_67_79 gnd C_bl
Cbb_67_79 bitb_67_79 gnd C_bl
Rb_67_80 bit_67_80 bit_67_81 R_bl
Rbb_67_80 bitb_67_80 bitb_67_81 R_bl
Cb_67_80 bit_67_80 gnd C_bl
Cbb_67_80 bitb_67_80 gnd C_bl
Rb_67_81 bit_67_81 bit_67_82 R_bl
Rbb_67_81 bitb_67_81 bitb_67_82 R_bl
Cb_67_81 bit_67_81 gnd C_bl
Cbb_67_81 bitb_67_81 gnd C_bl
Rb_67_82 bit_67_82 bit_67_83 R_bl
Rbb_67_82 bitb_67_82 bitb_67_83 R_bl
Cb_67_82 bit_67_82 gnd C_bl
Cbb_67_82 bitb_67_82 gnd C_bl
Rb_67_83 bit_67_83 bit_67_84 R_bl
Rbb_67_83 bitb_67_83 bitb_67_84 R_bl
Cb_67_83 bit_67_83 gnd C_bl
Cbb_67_83 bitb_67_83 gnd C_bl
Rb_67_84 bit_67_84 bit_67_85 R_bl
Rbb_67_84 bitb_67_84 bitb_67_85 R_bl
Cb_67_84 bit_67_84 gnd C_bl
Cbb_67_84 bitb_67_84 gnd C_bl
Rb_67_85 bit_67_85 bit_67_86 R_bl
Rbb_67_85 bitb_67_85 bitb_67_86 R_bl
Cb_67_85 bit_67_85 gnd C_bl
Cbb_67_85 bitb_67_85 gnd C_bl
Rb_67_86 bit_67_86 bit_67_87 R_bl
Rbb_67_86 bitb_67_86 bitb_67_87 R_bl
Cb_67_86 bit_67_86 gnd C_bl
Cbb_67_86 bitb_67_86 gnd C_bl
Rb_67_87 bit_67_87 bit_67_88 R_bl
Rbb_67_87 bitb_67_87 bitb_67_88 R_bl
Cb_67_87 bit_67_87 gnd C_bl
Cbb_67_87 bitb_67_87 gnd C_bl
Rb_67_88 bit_67_88 bit_67_89 R_bl
Rbb_67_88 bitb_67_88 bitb_67_89 R_bl
Cb_67_88 bit_67_88 gnd C_bl
Cbb_67_88 bitb_67_88 gnd C_bl
Rb_67_89 bit_67_89 bit_67_90 R_bl
Rbb_67_89 bitb_67_89 bitb_67_90 R_bl
Cb_67_89 bit_67_89 gnd C_bl
Cbb_67_89 bitb_67_89 gnd C_bl
Rb_67_90 bit_67_90 bit_67_91 R_bl
Rbb_67_90 bitb_67_90 bitb_67_91 R_bl
Cb_67_90 bit_67_90 gnd C_bl
Cbb_67_90 bitb_67_90 gnd C_bl
Rb_67_91 bit_67_91 bit_67_92 R_bl
Rbb_67_91 bitb_67_91 bitb_67_92 R_bl
Cb_67_91 bit_67_91 gnd C_bl
Cbb_67_91 bitb_67_91 gnd C_bl
Rb_67_92 bit_67_92 bit_67_93 R_bl
Rbb_67_92 bitb_67_92 bitb_67_93 R_bl
Cb_67_92 bit_67_92 gnd C_bl
Cbb_67_92 bitb_67_92 gnd C_bl
Rb_67_93 bit_67_93 bit_67_94 R_bl
Rbb_67_93 bitb_67_93 bitb_67_94 R_bl
Cb_67_93 bit_67_93 gnd C_bl
Cbb_67_93 bitb_67_93 gnd C_bl
Rb_67_94 bit_67_94 bit_67_95 R_bl
Rbb_67_94 bitb_67_94 bitb_67_95 R_bl
Cb_67_94 bit_67_94 gnd C_bl
Cbb_67_94 bitb_67_94 gnd C_bl
Rb_67_95 bit_67_95 bit_67_96 R_bl
Rbb_67_95 bitb_67_95 bitb_67_96 R_bl
Cb_67_95 bit_67_95 gnd C_bl
Cbb_67_95 bitb_67_95 gnd C_bl
Rb_67_96 bit_67_96 bit_67_97 R_bl
Rbb_67_96 bitb_67_96 bitb_67_97 R_bl
Cb_67_96 bit_67_96 gnd C_bl
Cbb_67_96 bitb_67_96 gnd C_bl
Rb_67_97 bit_67_97 bit_67_98 R_bl
Rbb_67_97 bitb_67_97 bitb_67_98 R_bl
Cb_67_97 bit_67_97 gnd C_bl
Cbb_67_97 bitb_67_97 gnd C_bl
Rb_67_98 bit_67_98 bit_67_99 R_bl
Rbb_67_98 bitb_67_98 bitb_67_99 R_bl
Cb_67_98 bit_67_98 gnd C_bl
Cbb_67_98 bitb_67_98 gnd C_bl
Rb_67_99 bit_67_99 bit_67_100 R_bl
Rbb_67_99 bitb_67_99 bitb_67_100 R_bl
Cb_67_99 bit_67_99 gnd C_bl
Cbb_67_99 bitb_67_99 gnd C_bl
Rb_68_0 bit_68_0 bit_68_1 R_bl
Rbb_68_0 bitb_68_0 bitb_68_1 R_bl
Cb_68_0 bit_68_0 gnd C_bl
Cbb_68_0 bitb_68_0 gnd C_bl
Rb_68_1 bit_68_1 bit_68_2 R_bl
Rbb_68_1 bitb_68_1 bitb_68_2 R_bl
Cb_68_1 bit_68_1 gnd C_bl
Cbb_68_1 bitb_68_1 gnd C_bl
Rb_68_2 bit_68_2 bit_68_3 R_bl
Rbb_68_2 bitb_68_2 bitb_68_3 R_bl
Cb_68_2 bit_68_2 gnd C_bl
Cbb_68_2 bitb_68_2 gnd C_bl
Rb_68_3 bit_68_3 bit_68_4 R_bl
Rbb_68_3 bitb_68_3 bitb_68_4 R_bl
Cb_68_3 bit_68_3 gnd C_bl
Cbb_68_3 bitb_68_3 gnd C_bl
Rb_68_4 bit_68_4 bit_68_5 R_bl
Rbb_68_4 bitb_68_4 bitb_68_5 R_bl
Cb_68_4 bit_68_4 gnd C_bl
Cbb_68_4 bitb_68_4 gnd C_bl
Rb_68_5 bit_68_5 bit_68_6 R_bl
Rbb_68_5 bitb_68_5 bitb_68_6 R_bl
Cb_68_5 bit_68_5 gnd C_bl
Cbb_68_5 bitb_68_5 gnd C_bl
Rb_68_6 bit_68_6 bit_68_7 R_bl
Rbb_68_6 bitb_68_6 bitb_68_7 R_bl
Cb_68_6 bit_68_6 gnd C_bl
Cbb_68_6 bitb_68_6 gnd C_bl
Rb_68_7 bit_68_7 bit_68_8 R_bl
Rbb_68_7 bitb_68_7 bitb_68_8 R_bl
Cb_68_7 bit_68_7 gnd C_bl
Cbb_68_7 bitb_68_7 gnd C_bl
Rb_68_8 bit_68_8 bit_68_9 R_bl
Rbb_68_8 bitb_68_8 bitb_68_9 R_bl
Cb_68_8 bit_68_8 gnd C_bl
Cbb_68_8 bitb_68_8 gnd C_bl
Rb_68_9 bit_68_9 bit_68_10 R_bl
Rbb_68_9 bitb_68_9 bitb_68_10 R_bl
Cb_68_9 bit_68_9 gnd C_bl
Cbb_68_9 bitb_68_9 gnd C_bl
Rb_68_10 bit_68_10 bit_68_11 R_bl
Rbb_68_10 bitb_68_10 bitb_68_11 R_bl
Cb_68_10 bit_68_10 gnd C_bl
Cbb_68_10 bitb_68_10 gnd C_bl
Rb_68_11 bit_68_11 bit_68_12 R_bl
Rbb_68_11 bitb_68_11 bitb_68_12 R_bl
Cb_68_11 bit_68_11 gnd C_bl
Cbb_68_11 bitb_68_11 gnd C_bl
Rb_68_12 bit_68_12 bit_68_13 R_bl
Rbb_68_12 bitb_68_12 bitb_68_13 R_bl
Cb_68_12 bit_68_12 gnd C_bl
Cbb_68_12 bitb_68_12 gnd C_bl
Rb_68_13 bit_68_13 bit_68_14 R_bl
Rbb_68_13 bitb_68_13 bitb_68_14 R_bl
Cb_68_13 bit_68_13 gnd C_bl
Cbb_68_13 bitb_68_13 gnd C_bl
Rb_68_14 bit_68_14 bit_68_15 R_bl
Rbb_68_14 bitb_68_14 bitb_68_15 R_bl
Cb_68_14 bit_68_14 gnd C_bl
Cbb_68_14 bitb_68_14 gnd C_bl
Rb_68_15 bit_68_15 bit_68_16 R_bl
Rbb_68_15 bitb_68_15 bitb_68_16 R_bl
Cb_68_15 bit_68_15 gnd C_bl
Cbb_68_15 bitb_68_15 gnd C_bl
Rb_68_16 bit_68_16 bit_68_17 R_bl
Rbb_68_16 bitb_68_16 bitb_68_17 R_bl
Cb_68_16 bit_68_16 gnd C_bl
Cbb_68_16 bitb_68_16 gnd C_bl
Rb_68_17 bit_68_17 bit_68_18 R_bl
Rbb_68_17 bitb_68_17 bitb_68_18 R_bl
Cb_68_17 bit_68_17 gnd C_bl
Cbb_68_17 bitb_68_17 gnd C_bl
Rb_68_18 bit_68_18 bit_68_19 R_bl
Rbb_68_18 bitb_68_18 bitb_68_19 R_bl
Cb_68_18 bit_68_18 gnd C_bl
Cbb_68_18 bitb_68_18 gnd C_bl
Rb_68_19 bit_68_19 bit_68_20 R_bl
Rbb_68_19 bitb_68_19 bitb_68_20 R_bl
Cb_68_19 bit_68_19 gnd C_bl
Cbb_68_19 bitb_68_19 gnd C_bl
Rb_68_20 bit_68_20 bit_68_21 R_bl
Rbb_68_20 bitb_68_20 bitb_68_21 R_bl
Cb_68_20 bit_68_20 gnd C_bl
Cbb_68_20 bitb_68_20 gnd C_bl
Rb_68_21 bit_68_21 bit_68_22 R_bl
Rbb_68_21 bitb_68_21 bitb_68_22 R_bl
Cb_68_21 bit_68_21 gnd C_bl
Cbb_68_21 bitb_68_21 gnd C_bl
Rb_68_22 bit_68_22 bit_68_23 R_bl
Rbb_68_22 bitb_68_22 bitb_68_23 R_bl
Cb_68_22 bit_68_22 gnd C_bl
Cbb_68_22 bitb_68_22 gnd C_bl
Rb_68_23 bit_68_23 bit_68_24 R_bl
Rbb_68_23 bitb_68_23 bitb_68_24 R_bl
Cb_68_23 bit_68_23 gnd C_bl
Cbb_68_23 bitb_68_23 gnd C_bl
Rb_68_24 bit_68_24 bit_68_25 R_bl
Rbb_68_24 bitb_68_24 bitb_68_25 R_bl
Cb_68_24 bit_68_24 gnd C_bl
Cbb_68_24 bitb_68_24 gnd C_bl
Rb_68_25 bit_68_25 bit_68_26 R_bl
Rbb_68_25 bitb_68_25 bitb_68_26 R_bl
Cb_68_25 bit_68_25 gnd C_bl
Cbb_68_25 bitb_68_25 gnd C_bl
Rb_68_26 bit_68_26 bit_68_27 R_bl
Rbb_68_26 bitb_68_26 bitb_68_27 R_bl
Cb_68_26 bit_68_26 gnd C_bl
Cbb_68_26 bitb_68_26 gnd C_bl
Rb_68_27 bit_68_27 bit_68_28 R_bl
Rbb_68_27 bitb_68_27 bitb_68_28 R_bl
Cb_68_27 bit_68_27 gnd C_bl
Cbb_68_27 bitb_68_27 gnd C_bl
Rb_68_28 bit_68_28 bit_68_29 R_bl
Rbb_68_28 bitb_68_28 bitb_68_29 R_bl
Cb_68_28 bit_68_28 gnd C_bl
Cbb_68_28 bitb_68_28 gnd C_bl
Rb_68_29 bit_68_29 bit_68_30 R_bl
Rbb_68_29 bitb_68_29 bitb_68_30 R_bl
Cb_68_29 bit_68_29 gnd C_bl
Cbb_68_29 bitb_68_29 gnd C_bl
Rb_68_30 bit_68_30 bit_68_31 R_bl
Rbb_68_30 bitb_68_30 bitb_68_31 R_bl
Cb_68_30 bit_68_30 gnd C_bl
Cbb_68_30 bitb_68_30 gnd C_bl
Rb_68_31 bit_68_31 bit_68_32 R_bl
Rbb_68_31 bitb_68_31 bitb_68_32 R_bl
Cb_68_31 bit_68_31 gnd C_bl
Cbb_68_31 bitb_68_31 gnd C_bl
Rb_68_32 bit_68_32 bit_68_33 R_bl
Rbb_68_32 bitb_68_32 bitb_68_33 R_bl
Cb_68_32 bit_68_32 gnd C_bl
Cbb_68_32 bitb_68_32 gnd C_bl
Rb_68_33 bit_68_33 bit_68_34 R_bl
Rbb_68_33 bitb_68_33 bitb_68_34 R_bl
Cb_68_33 bit_68_33 gnd C_bl
Cbb_68_33 bitb_68_33 gnd C_bl
Rb_68_34 bit_68_34 bit_68_35 R_bl
Rbb_68_34 bitb_68_34 bitb_68_35 R_bl
Cb_68_34 bit_68_34 gnd C_bl
Cbb_68_34 bitb_68_34 gnd C_bl
Rb_68_35 bit_68_35 bit_68_36 R_bl
Rbb_68_35 bitb_68_35 bitb_68_36 R_bl
Cb_68_35 bit_68_35 gnd C_bl
Cbb_68_35 bitb_68_35 gnd C_bl
Rb_68_36 bit_68_36 bit_68_37 R_bl
Rbb_68_36 bitb_68_36 bitb_68_37 R_bl
Cb_68_36 bit_68_36 gnd C_bl
Cbb_68_36 bitb_68_36 gnd C_bl
Rb_68_37 bit_68_37 bit_68_38 R_bl
Rbb_68_37 bitb_68_37 bitb_68_38 R_bl
Cb_68_37 bit_68_37 gnd C_bl
Cbb_68_37 bitb_68_37 gnd C_bl
Rb_68_38 bit_68_38 bit_68_39 R_bl
Rbb_68_38 bitb_68_38 bitb_68_39 R_bl
Cb_68_38 bit_68_38 gnd C_bl
Cbb_68_38 bitb_68_38 gnd C_bl
Rb_68_39 bit_68_39 bit_68_40 R_bl
Rbb_68_39 bitb_68_39 bitb_68_40 R_bl
Cb_68_39 bit_68_39 gnd C_bl
Cbb_68_39 bitb_68_39 gnd C_bl
Rb_68_40 bit_68_40 bit_68_41 R_bl
Rbb_68_40 bitb_68_40 bitb_68_41 R_bl
Cb_68_40 bit_68_40 gnd C_bl
Cbb_68_40 bitb_68_40 gnd C_bl
Rb_68_41 bit_68_41 bit_68_42 R_bl
Rbb_68_41 bitb_68_41 bitb_68_42 R_bl
Cb_68_41 bit_68_41 gnd C_bl
Cbb_68_41 bitb_68_41 gnd C_bl
Rb_68_42 bit_68_42 bit_68_43 R_bl
Rbb_68_42 bitb_68_42 bitb_68_43 R_bl
Cb_68_42 bit_68_42 gnd C_bl
Cbb_68_42 bitb_68_42 gnd C_bl
Rb_68_43 bit_68_43 bit_68_44 R_bl
Rbb_68_43 bitb_68_43 bitb_68_44 R_bl
Cb_68_43 bit_68_43 gnd C_bl
Cbb_68_43 bitb_68_43 gnd C_bl
Rb_68_44 bit_68_44 bit_68_45 R_bl
Rbb_68_44 bitb_68_44 bitb_68_45 R_bl
Cb_68_44 bit_68_44 gnd C_bl
Cbb_68_44 bitb_68_44 gnd C_bl
Rb_68_45 bit_68_45 bit_68_46 R_bl
Rbb_68_45 bitb_68_45 bitb_68_46 R_bl
Cb_68_45 bit_68_45 gnd C_bl
Cbb_68_45 bitb_68_45 gnd C_bl
Rb_68_46 bit_68_46 bit_68_47 R_bl
Rbb_68_46 bitb_68_46 bitb_68_47 R_bl
Cb_68_46 bit_68_46 gnd C_bl
Cbb_68_46 bitb_68_46 gnd C_bl
Rb_68_47 bit_68_47 bit_68_48 R_bl
Rbb_68_47 bitb_68_47 bitb_68_48 R_bl
Cb_68_47 bit_68_47 gnd C_bl
Cbb_68_47 bitb_68_47 gnd C_bl
Rb_68_48 bit_68_48 bit_68_49 R_bl
Rbb_68_48 bitb_68_48 bitb_68_49 R_bl
Cb_68_48 bit_68_48 gnd C_bl
Cbb_68_48 bitb_68_48 gnd C_bl
Rb_68_49 bit_68_49 bit_68_50 R_bl
Rbb_68_49 bitb_68_49 bitb_68_50 R_bl
Cb_68_49 bit_68_49 gnd C_bl
Cbb_68_49 bitb_68_49 gnd C_bl
Rb_68_50 bit_68_50 bit_68_51 R_bl
Rbb_68_50 bitb_68_50 bitb_68_51 R_bl
Cb_68_50 bit_68_50 gnd C_bl
Cbb_68_50 bitb_68_50 gnd C_bl
Rb_68_51 bit_68_51 bit_68_52 R_bl
Rbb_68_51 bitb_68_51 bitb_68_52 R_bl
Cb_68_51 bit_68_51 gnd C_bl
Cbb_68_51 bitb_68_51 gnd C_bl
Rb_68_52 bit_68_52 bit_68_53 R_bl
Rbb_68_52 bitb_68_52 bitb_68_53 R_bl
Cb_68_52 bit_68_52 gnd C_bl
Cbb_68_52 bitb_68_52 gnd C_bl
Rb_68_53 bit_68_53 bit_68_54 R_bl
Rbb_68_53 bitb_68_53 bitb_68_54 R_bl
Cb_68_53 bit_68_53 gnd C_bl
Cbb_68_53 bitb_68_53 gnd C_bl
Rb_68_54 bit_68_54 bit_68_55 R_bl
Rbb_68_54 bitb_68_54 bitb_68_55 R_bl
Cb_68_54 bit_68_54 gnd C_bl
Cbb_68_54 bitb_68_54 gnd C_bl
Rb_68_55 bit_68_55 bit_68_56 R_bl
Rbb_68_55 bitb_68_55 bitb_68_56 R_bl
Cb_68_55 bit_68_55 gnd C_bl
Cbb_68_55 bitb_68_55 gnd C_bl
Rb_68_56 bit_68_56 bit_68_57 R_bl
Rbb_68_56 bitb_68_56 bitb_68_57 R_bl
Cb_68_56 bit_68_56 gnd C_bl
Cbb_68_56 bitb_68_56 gnd C_bl
Rb_68_57 bit_68_57 bit_68_58 R_bl
Rbb_68_57 bitb_68_57 bitb_68_58 R_bl
Cb_68_57 bit_68_57 gnd C_bl
Cbb_68_57 bitb_68_57 gnd C_bl
Rb_68_58 bit_68_58 bit_68_59 R_bl
Rbb_68_58 bitb_68_58 bitb_68_59 R_bl
Cb_68_58 bit_68_58 gnd C_bl
Cbb_68_58 bitb_68_58 gnd C_bl
Rb_68_59 bit_68_59 bit_68_60 R_bl
Rbb_68_59 bitb_68_59 bitb_68_60 R_bl
Cb_68_59 bit_68_59 gnd C_bl
Cbb_68_59 bitb_68_59 gnd C_bl
Rb_68_60 bit_68_60 bit_68_61 R_bl
Rbb_68_60 bitb_68_60 bitb_68_61 R_bl
Cb_68_60 bit_68_60 gnd C_bl
Cbb_68_60 bitb_68_60 gnd C_bl
Rb_68_61 bit_68_61 bit_68_62 R_bl
Rbb_68_61 bitb_68_61 bitb_68_62 R_bl
Cb_68_61 bit_68_61 gnd C_bl
Cbb_68_61 bitb_68_61 gnd C_bl
Rb_68_62 bit_68_62 bit_68_63 R_bl
Rbb_68_62 bitb_68_62 bitb_68_63 R_bl
Cb_68_62 bit_68_62 gnd C_bl
Cbb_68_62 bitb_68_62 gnd C_bl
Rb_68_63 bit_68_63 bit_68_64 R_bl
Rbb_68_63 bitb_68_63 bitb_68_64 R_bl
Cb_68_63 bit_68_63 gnd C_bl
Cbb_68_63 bitb_68_63 gnd C_bl
Rb_68_64 bit_68_64 bit_68_65 R_bl
Rbb_68_64 bitb_68_64 bitb_68_65 R_bl
Cb_68_64 bit_68_64 gnd C_bl
Cbb_68_64 bitb_68_64 gnd C_bl
Rb_68_65 bit_68_65 bit_68_66 R_bl
Rbb_68_65 bitb_68_65 bitb_68_66 R_bl
Cb_68_65 bit_68_65 gnd C_bl
Cbb_68_65 bitb_68_65 gnd C_bl
Rb_68_66 bit_68_66 bit_68_67 R_bl
Rbb_68_66 bitb_68_66 bitb_68_67 R_bl
Cb_68_66 bit_68_66 gnd C_bl
Cbb_68_66 bitb_68_66 gnd C_bl
Rb_68_67 bit_68_67 bit_68_68 R_bl
Rbb_68_67 bitb_68_67 bitb_68_68 R_bl
Cb_68_67 bit_68_67 gnd C_bl
Cbb_68_67 bitb_68_67 gnd C_bl
Rb_68_68 bit_68_68 bit_68_69 R_bl
Rbb_68_68 bitb_68_68 bitb_68_69 R_bl
Cb_68_68 bit_68_68 gnd C_bl
Cbb_68_68 bitb_68_68 gnd C_bl
Rb_68_69 bit_68_69 bit_68_70 R_bl
Rbb_68_69 bitb_68_69 bitb_68_70 R_bl
Cb_68_69 bit_68_69 gnd C_bl
Cbb_68_69 bitb_68_69 gnd C_bl
Rb_68_70 bit_68_70 bit_68_71 R_bl
Rbb_68_70 bitb_68_70 bitb_68_71 R_bl
Cb_68_70 bit_68_70 gnd C_bl
Cbb_68_70 bitb_68_70 gnd C_bl
Rb_68_71 bit_68_71 bit_68_72 R_bl
Rbb_68_71 bitb_68_71 bitb_68_72 R_bl
Cb_68_71 bit_68_71 gnd C_bl
Cbb_68_71 bitb_68_71 gnd C_bl
Rb_68_72 bit_68_72 bit_68_73 R_bl
Rbb_68_72 bitb_68_72 bitb_68_73 R_bl
Cb_68_72 bit_68_72 gnd C_bl
Cbb_68_72 bitb_68_72 gnd C_bl
Rb_68_73 bit_68_73 bit_68_74 R_bl
Rbb_68_73 bitb_68_73 bitb_68_74 R_bl
Cb_68_73 bit_68_73 gnd C_bl
Cbb_68_73 bitb_68_73 gnd C_bl
Rb_68_74 bit_68_74 bit_68_75 R_bl
Rbb_68_74 bitb_68_74 bitb_68_75 R_bl
Cb_68_74 bit_68_74 gnd C_bl
Cbb_68_74 bitb_68_74 gnd C_bl
Rb_68_75 bit_68_75 bit_68_76 R_bl
Rbb_68_75 bitb_68_75 bitb_68_76 R_bl
Cb_68_75 bit_68_75 gnd C_bl
Cbb_68_75 bitb_68_75 gnd C_bl
Rb_68_76 bit_68_76 bit_68_77 R_bl
Rbb_68_76 bitb_68_76 bitb_68_77 R_bl
Cb_68_76 bit_68_76 gnd C_bl
Cbb_68_76 bitb_68_76 gnd C_bl
Rb_68_77 bit_68_77 bit_68_78 R_bl
Rbb_68_77 bitb_68_77 bitb_68_78 R_bl
Cb_68_77 bit_68_77 gnd C_bl
Cbb_68_77 bitb_68_77 gnd C_bl
Rb_68_78 bit_68_78 bit_68_79 R_bl
Rbb_68_78 bitb_68_78 bitb_68_79 R_bl
Cb_68_78 bit_68_78 gnd C_bl
Cbb_68_78 bitb_68_78 gnd C_bl
Rb_68_79 bit_68_79 bit_68_80 R_bl
Rbb_68_79 bitb_68_79 bitb_68_80 R_bl
Cb_68_79 bit_68_79 gnd C_bl
Cbb_68_79 bitb_68_79 gnd C_bl
Rb_68_80 bit_68_80 bit_68_81 R_bl
Rbb_68_80 bitb_68_80 bitb_68_81 R_bl
Cb_68_80 bit_68_80 gnd C_bl
Cbb_68_80 bitb_68_80 gnd C_bl
Rb_68_81 bit_68_81 bit_68_82 R_bl
Rbb_68_81 bitb_68_81 bitb_68_82 R_bl
Cb_68_81 bit_68_81 gnd C_bl
Cbb_68_81 bitb_68_81 gnd C_bl
Rb_68_82 bit_68_82 bit_68_83 R_bl
Rbb_68_82 bitb_68_82 bitb_68_83 R_bl
Cb_68_82 bit_68_82 gnd C_bl
Cbb_68_82 bitb_68_82 gnd C_bl
Rb_68_83 bit_68_83 bit_68_84 R_bl
Rbb_68_83 bitb_68_83 bitb_68_84 R_bl
Cb_68_83 bit_68_83 gnd C_bl
Cbb_68_83 bitb_68_83 gnd C_bl
Rb_68_84 bit_68_84 bit_68_85 R_bl
Rbb_68_84 bitb_68_84 bitb_68_85 R_bl
Cb_68_84 bit_68_84 gnd C_bl
Cbb_68_84 bitb_68_84 gnd C_bl
Rb_68_85 bit_68_85 bit_68_86 R_bl
Rbb_68_85 bitb_68_85 bitb_68_86 R_bl
Cb_68_85 bit_68_85 gnd C_bl
Cbb_68_85 bitb_68_85 gnd C_bl
Rb_68_86 bit_68_86 bit_68_87 R_bl
Rbb_68_86 bitb_68_86 bitb_68_87 R_bl
Cb_68_86 bit_68_86 gnd C_bl
Cbb_68_86 bitb_68_86 gnd C_bl
Rb_68_87 bit_68_87 bit_68_88 R_bl
Rbb_68_87 bitb_68_87 bitb_68_88 R_bl
Cb_68_87 bit_68_87 gnd C_bl
Cbb_68_87 bitb_68_87 gnd C_bl
Rb_68_88 bit_68_88 bit_68_89 R_bl
Rbb_68_88 bitb_68_88 bitb_68_89 R_bl
Cb_68_88 bit_68_88 gnd C_bl
Cbb_68_88 bitb_68_88 gnd C_bl
Rb_68_89 bit_68_89 bit_68_90 R_bl
Rbb_68_89 bitb_68_89 bitb_68_90 R_bl
Cb_68_89 bit_68_89 gnd C_bl
Cbb_68_89 bitb_68_89 gnd C_bl
Rb_68_90 bit_68_90 bit_68_91 R_bl
Rbb_68_90 bitb_68_90 bitb_68_91 R_bl
Cb_68_90 bit_68_90 gnd C_bl
Cbb_68_90 bitb_68_90 gnd C_bl
Rb_68_91 bit_68_91 bit_68_92 R_bl
Rbb_68_91 bitb_68_91 bitb_68_92 R_bl
Cb_68_91 bit_68_91 gnd C_bl
Cbb_68_91 bitb_68_91 gnd C_bl
Rb_68_92 bit_68_92 bit_68_93 R_bl
Rbb_68_92 bitb_68_92 bitb_68_93 R_bl
Cb_68_92 bit_68_92 gnd C_bl
Cbb_68_92 bitb_68_92 gnd C_bl
Rb_68_93 bit_68_93 bit_68_94 R_bl
Rbb_68_93 bitb_68_93 bitb_68_94 R_bl
Cb_68_93 bit_68_93 gnd C_bl
Cbb_68_93 bitb_68_93 gnd C_bl
Rb_68_94 bit_68_94 bit_68_95 R_bl
Rbb_68_94 bitb_68_94 bitb_68_95 R_bl
Cb_68_94 bit_68_94 gnd C_bl
Cbb_68_94 bitb_68_94 gnd C_bl
Rb_68_95 bit_68_95 bit_68_96 R_bl
Rbb_68_95 bitb_68_95 bitb_68_96 R_bl
Cb_68_95 bit_68_95 gnd C_bl
Cbb_68_95 bitb_68_95 gnd C_bl
Rb_68_96 bit_68_96 bit_68_97 R_bl
Rbb_68_96 bitb_68_96 bitb_68_97 R_bl
Cb_68_96 bit_68_96 gnd C_bl
Cbb_68_96 bitb_68_96 gnd C_bl
Rb_68_97 bit_68_97 bit_68_98 R_bl
Rbb_68_97 bitb_68_97 bitb_68_98 R_bl
Cb_68_97 bit_68_97 gnd C_bl
Cbb_68_97 bitb_68_97 gnd C_bl
Rb_68_98 bit_68_98 bit_68_99 R_bl
Rbb_68_98 bitb_68_98 bitb_68_99 R_bl
Cb_68_98 bit_68_98 gnd C_bl
Cbb_68_98 bitb_68_98 gnd C_bl
Rb_68_99 bit_68_99 bit_68_100 R_bl
Rbb_68_99 bitb_68_99 bitb_68_100 R_bl
Cb_68_99 bit_68_99 gnd C_bl
Cbb_68_99 bitb_68_99 gnd C_bl
Rb_69_0 bit_69_0 bit_69_1 R_bl
Rbb_69_0 bitb_69_0 bitb_69_1 R_bl
Cb_69_0 bit_69_0 gnd C_bl
Cbb_69_0 bitb_69_0 gnd C_bl
Rb_69_1 bit_69_1 bit_69_2 R_bl
Rbb_69_1 bitb_69_1 bitb_69_2 R_bl
Cb_69_1 bit_69_1 gnd C_bl
Cbb_69_1 bitb_69_1 gnd C_bl
Rb_69_2 bit_69_2 bit_69_3 R_bl
Rbb_69_2 bitb_69_2 bitb_69_3 R_bl
Cb_69_2 bit_69_2 gnd C_bl
Cbb_69_2 bitb_69_2 gnd C_bl
Rb_69_3 bit_69_3 bit_69_4 R_bl
Rbb_69_3 bitb_69_3 bitb_69_4 R_bl
Cb_69_3 bit_69_3 gnd C_bl
Cbb_69_3 bitb_69_3 gnd C_bl
Rb_69_4 bit_69_4 bit_69_5 R_bl
Rbb_69_4 bitb_69_4 bitb_69_5 R_bl
Cb_69_4 bit_69_4 gnd C_bl
Cbb_69_4 bitb_69_4 gnd C_bl
Rb_69_5 bit_69_5 bit_69_6 R_bl
Rbb_69_5 bitb_69_5 bitb_69_6 R_bl
Cb_69_5 bit_69_5 gnd C_bl
Cbb_69_5 bitb_69_5 gnd C_bl
Rb_69_6 bit_69_6 bit_69_7 R_bl
Rbb_69_6 bitb_69_6 bitb_69_7 R_bl
Cb_69_6 bit_69_6 gnd C_bl
Cbb_69_6 bitb_69_6 gnd C_bl
Rb_69_7 bit_69_7 bit_69_8 R_bl
Rbb_69_7 bitb_69_7 bitb_69_8 R_bl
Cb_69_7 bit_69_7 gnd C_bl
Cbb_69_7 bitb_69_7 gnd C_bl
Rb_69_8 bit_69_8 bit_69_9 R_bl
Rbb_69_8 bitb_69_8 bitb_69_9 R_bl
Cb_69_8 bit_69_8 gnd C_bl
Cbb_69_8 bitb_69_8 gnd C_bl
Rb_69_9 bit_69_9 bit_69_10 R_bl
Rbb_69_9 bitb_69_9 bitb_69_10 R_bl
Cb_69_9 bit_69_9 gnd C_bl
Cbb_69_9 bitb_69_9 gnd C_bl
Rb_69_10 bit_69_10 bit_69_11 R_bl
Rbb_69_10 bitb_69_10 bitb_69_11 R_bl
Cb_69_10 bit_69_10 gnd C_bl
Cbb_69_10 bitb_69_10 gnd C_bl
Rb_69_11 bit_69_11 bit_69_12 R_bl
Rbb_69_11 bitb_69_11 bitb_69_12 R_bl
Cb_69_11 bit_69_11 gnd C_bl
Cbb_69_11 bitb_69_11 gnd C_bl
Rb_69_12 bit_69_12 bit_69_13 R_bl
Rbb_69_12 bitb_69_12 bitb_69_13 R_bl
Cb_69_12 bit_69_12 gnd C_bl
Cbb_69_12 bitb_69_12 gnd C_bl
Rb_69_13 bit_69_13 bit_69_14 R_bl
Rbb_69_13 bitb_69_13 bitb_69_14 R_bl
Cb_69_13 bit_69_13 gnd C_bl
Cbb_69_13 bitb_69_13 gnd C_bl
Rb_69_14 bit_69_14 bit_69_15 R_bl
Rbb_69_14 bitb_69_14 bitb_69_15 R_bl
Cb_69_14 bit_69_14 gnd C_bl
Cbb_69_14 bitb_69_14 gnd C_bl
Rb_69_15 bit_69_15 bit_69_16 R_bl
Rbb_69_15 bitb_69_15 bitb_69_16 R_bl
Cb_69_15 bit_69_15 gnd C_bl
Cbb_69_15 bitb_69_15 gnd C_bl
Rb_69_16 bit_69_16 bit_69_17 R_bl
Rbb_69_16 bitb_69_16 bitb_69_17 R_bl
Cb_69_16 bit_69_16 gnd C_bl
Cbb_69_16 bitb_69_16 gnd C_bl
Rb_69_17 bit_69_17 bit_69_18 R_bl
Rbb_69_17 bitb_69_17 bitb_69_18 R_bl
Cb_69_17 bit_69_17 gnd C_bl
Cbb_69_17 bitb_69_17 gnd C_bl
Rb_69_18 bit_69_18 bit_69_19 R_bl
Rbb_69_18 bitb_69_18 bitb_69_19 R_bl
Cb_69_18 bit_69_18 gnd C_bl
Cbb_69_18 bitb_69_18 gnd C_bl
Rb_69_19 bit_69_19 bit_69_20 R_bl
Rbb_69_19 bitb_69_19 bitb_69_20 R_bl
Cb_69_19 bit_69_19 gnd C_bl
Cbb_69_19 bitb_69_19 gnd C_bl
Rb_69_20 bit_69_20 bit_69_21 R_bl
Rbb_69_20 bitb_69_20 bitb_69_21 R_bl
Cb_69_20 bit_69_20 gnd C_bl
Cbb_69_20 bitb_69_20 gnd C_bl
Rb_69_21 bit_69_21 bit_69_22 R_bl
Rbb_69_21 bitb_69_21 bitb_69_22 R_bl
Cb_69_21 bit_69_21 gnd C_bl
Cbb_69_21 bitb_69_21 gnd C_bl
Rb_69_22 bit_69_22 bit_69_23 R_bl
Rbb_69_22 bitb_69_22 bitb_69_23 R_bl
Cb_69_22 bit_69_22 gnd C_bl
Cbb_69_22 bitb_69_22 gnd C_bl
Rb_69_23 bit_69_23 bit_69_24 R_bl
Rbb_69_23 bitb_69_23 bitb_69_24 R_bl
Cb_69_23 bit_69_23 gnd C_bl
Cbb_69_23 bitb_69_23 gnd C_bl
Rb_69_24 bit_69_24 bit_69_25 R_bl
Rbb_69_24 bitb_69_24 bitb_69_25 R_bl
Cb_69_24 bit_69_24 gnd C_bl
Cbb_69_24 bitb_69_24 gnd C_bl
Rb_69_25 bit_69_25 bit_69_26 R_bl
Rbb_69_25 bitb_69_25 bitb_69_26 R_bl
Cb_69_25 bit_69_25 gnd C_bl
Cbb_69_25 bitb_69_25 gnd C_bl
Rb_69_26 bit_69_26 bit_69_27 R_bl
Rbb_69_26 bitb_69_26 bitb_69_27 R_bl
Cb_69_26 bit_69_26 gnd C_bl
Cbb_69_26 bitb_69_26 gnd C_bl
Rb_69_27 bit_69_27 bit_69_28 R_bl
Rbb_69_27 bitb_69_27 bitb_69_28 R_bl
Cb_69_27 bit_69_27 gnd C_bl
Cbb_69_27 bitb_69_27 gnd C_bl
Rb_69_28 bit_69_28 bit_69_29 R_bl
Rbb_69_28 bitb_69_28 bitb_69_29 R_bl
Cb_69_28 bit_69_28 gnd C_bl
Cbb_69_28 bitb_69_28 gnd C_bl
Rb_69_29 bit_69_29 bit_69_30 R_bl
Rbb_69_29 bitb_69_29 bitb_69_30 R_bl
Cb_69_29 bit_69_29 gnd C_bl
Cbb_69_29 bitb_69_29 gnd C_bl
Rb_69_30 bit_69_30 bit_69_31 R_bl
Rbb_69_30 bitb_69_30 bitb_69_31 R_bl
Cb_69_30 bit_69_30 gnd C_bl
Cbb_69_30 bitb_69_30 gnd C_bl
Rb_69_31 bit_69_31 bit_69_32 R_bl
Rbb_69_31 bitb_69_31 bitb_69_32 R_bl
Cb_69_31 bit_69_31 gnd C_bl
Cbb_69_31 bitb_69_31 gnd C_bl
Rb_69_32 bit_69_32 bit_69_33 R_bl
Rbb_69_32 bitb_69_32 bitb_69_33 R_bl
Cb_69_32 bit_69_32 gnd C_bl
Cbb_69_32 bitb_69_32 gnd C_bl
Rb_69_33 bit_69_33 bit_69_34 R_bl
Rbb_69_33 bitb_69_33 bitb_69_34 R_bl
Cb_69_33 bit_69_33 gnd C_bl
Cbb_69_33 bitb_69_33 gnd C_bl
Rb_69_34 bit_69_34 bit_69_35 R_bl
Rbb_69_34 bitb_69_34 bitb_69_35 R_bl
Cb_69_34 bit_69_34 gnd C_bl
Cbb_69_34 bitb_69_34 gnd C_bl
Rb_69_35 bit_69_35 bit_69_36 R_bl
Rbb_69_35 bitb_69_35 bitb_69_36 R_bl
Cb_69_35 bit_69_35 gnd C_bl
Cbb_69_35 bitb_69_35 gnd C_bl
Rb_69_36 bit_69_36 bit_69_37 R_bl
Rbb_69_36 bitb_69_36 bitb_69_37 R_bl
Cb_69_36 bit_69_36 gnd C_bl
Cbb_69_36 bitb_69_36 gnd C_bl
Rb_69_37 bit_69_37 bit_69_38 R_bl
Rbb_69_37 bitb_69_37 bitb_69_38 R_bl
Cb_69_37 bit_69_37 gnd C_bl
Cbb_69_37 bitb_69_37 gnd C_bl
Rb_69_38 bit_69_38 bit_69_39 R_bl
Rbb_69_38 bitb_69_38 bitb_69_39 R_bl
Cb_69_38 bit_69_38 gnd C_bl
Cbb_69_38 bitb_69_38 gnd C_bl
Rb_69_39 bit_69_39 bit_69_40 R_bl
Rbb_69_39 bitb_69_39 bitb_69_40 R_bl
Cb_69_39 bit_69_39 gnd C_bl
Cbb_69_39 bitb_69_39 gnd C_bl
Rb_69_40 bit_69_40 bit_69_41 R_bl
Rbb_69_40 bitb_69_40 bitb_69_41 R_bl
Cb_69_40 bit_69_40 gnd C_bl
Cbb_69_40 bitb_69_40 gnd C_bl
Rb_69_41 bit_69_41 bit_69_42 R_bl
Rbb_69_41 bitb_69_41 bitb_69_42 R_bl
Cb_69_41 bit_69_41 gnd C_bl
Cbb_69_41 bitb_69_41 gnd C_bl
Rb_69_42 bit_69_42 bit_69_43 R_bl
Rbb_69_42 bitb_69_42 bitb_69_43 R_bl
Cb_69_42 bit_69_42 gnd C_bl
Cbb_69_42 bitb_69_42 gnd C_bl
Rb_69_43 bit_69_43 bit_69_44 R_bl
Rbb_69_43 bitb_69_43 bitb_69_44 R_bl
Cb_69_43 bit_69_43 gnd C_bl
Cbb_69_43 bitb_69_43 gnd C_bl
Rb_69_44 bit_69_44 bit_69_45 R_bl
Rbb_69_44 bitb_69_44 bitb_69_45 R_bl
Cb_69_44 bit_69_44 gnd C_bl
Cbb_69_44 bitb_69_44 gnd C_bl
Rb_69_45 bit_69_45 bit_69_46 R_bl
Rbb_69_45 bitb_69_45 bitb_69_46 R_bl
Cb_69_45 bit_69_45 gnd C_bl
Cbb_69_45 bitb_69_45 gnd C_bl
Rb_69_46 bit_69_46 bit_69_47 R_bl
Rbb_69_46 bitb_69_46 bitb_69_47 R_bl
Cb_69_46 bit_69_46 gnd C_bl
Cbb_69_46 bitb_69_46 gnd C_bl
Rb_69_47 bit_69_47 bit_69_48 R_bl
Rbb_69_47 bitb_69_47 bitb_69_48 R_bl
Cb_69_47 bit_69_47 gnd C_bl
Cbb_69_47 bitb_69_47 gnd C_bl
Rb_69_48 bit_69_48 bit_69_49 R_bl
Rbb_69_48 bitb_69_48 bitb_69_49 R_bl
Cb_69_48 bit_69_48 gnd C_bl
Cbb_69_48 bitb_69_48 gnd C_bl
Rb_69_49 bit_69_49 bit_69_50 R_bl
Rbb_69_49 bitb_69_49 bitb_69_50 R_bl
Cb_69_49 bit_69_49 gnd C_bl
Cbb_69_49 bitb_69_49 gnd C_bl
Rb_69_50 bit_69_50 bit_69_51 R_bl
Rbb_69_50 bitb_69_50 bitb_69_51 R_bl
Cb_69_50 bit_69_50 gnd C_bl
Cbb_69_50 bitb_69_50 gnd C_bl
Rb_69_51 bit_69_51 bit_69_52 R_bl
Rbb_69_51 bitb_69_51 bitb_69_52 R_bl
Cb_69_51 bit_69_51 gnd C_bl
Cbb_69_51 bitb_69_51 gnd C_bl
Rb_69_52 bit_69_52 bit_69_53 R_bl
Rbb_69_52 bitb_69_52 bitb_69_53 R_bl
Cb_69_52 bit_69_52 gnd C_bl
Cbb_69_52 bitb_69_52 gnd C_bl
Rb_69_53 bit_69_53 bit_69_54 R_bl
Rbb_69_53 bitb_69_53 bitb_69_54 R_bl
Cb_69_53 bit_69_53 gnd C_bl
Cbb_69_53 bitb_69_53 gnd C_bl
Rb_69_54 bit_69_54 bit_69_55 R_bl
Rbb_69_54 bitb_69_54 bitb_69_55 R_bl
Cb_69_54 bit_69_54 gnd C_bl
Cbb_69_54 bitb_69_54 gnd C_bl
Rb_69_55 bit_69_55 bit_69_56 R_bl
Rbb_69_55 bitb_69_55 bitb_69_56 R_bl
Cb_69_55 bit_69_55 gnd C_bl
Cbb_69_55 bitb_69_55 gnd C_bl
Rb_69_56 bit_69_56 bit_69_57 R_bl
Rbb_69_56 bitb_69_56 bitb_69_57 R_bl
Cb_69_56 bit_69_56 gnd C_bl
Cbb_69_56 bitb_69_56 gnd C_bl
Rb_69_57 bit_69_57 bit_69_58 R_bl
Rbb_69_57 bitb_69_57 bitb_69_58 R_bl
Cb_69_57 bit_69_57 gnd C_bl
Cbb_69_57 bitb_69_57 gnd C_bl
Rb_69_58 bit_69_58 bit_69_59 R_bl
Rbb_69_58 bitb_69_58 bitb_69_59 R_bl
Cb_69_58 bit_69_58 gnd C_bl
Cbb_69_58 bitb_69_58 gnd C_bl
Rb_69_59 bit_69_59 bit_69_60 R_bl
Rbb_69_59 bitb_69_59 bitb_69_60 R_bl
Cb_69_59 bit_69_59 gnd C_bl
Cbb_69_59 bitb_69_59 gnd C_bl
Rb_69_60 bit_69_60 bit_69_61 R_bl
Rbb_69_60 bitb_69_60 bitb_69_61 R_bl
Cb_69_60 bit_69_60 gnd C_bl
Cbb_69_60 bitb_69_60 gnd C_bl
Rb_69_61 bit_69_61 bit_69_62 R_bl
Rbb_69_61 bitb_69_61 bitb_69_62 R_bl
Cb_69_61 bit_69_61 gnd C_bl
Cbb_69_61 bitb_69_61 gnd C_bl
Rb_69_62 bit_69_62 bit_69_63 R_bl
Rbb_69_62 bitb_69_62 bitb_69_63 R_bl
Cb_69_62 bit_69_62 gnd C_bl
Cbb_69_62 bitb_69_62 gnd C_bl
Rb_69_63 bit_69_63 bit_69_64 R_bl
Rbb_69_63 bitb_69_63 bitb_69_64 R_bl
Cb_69_63 bit_69_63 gnd C_bl
Cbb_69_63 bitb_69_63 gnd C_bl
Rb_69_64 bit_69_64 bit_69_65 R_bl
Rbb_69_64 bitb_69_64 bitb_69_65 R_bl
Cb_69_64 bit_69_64 gnd C_bl
Cbb_69_64 bitb_69_64 gnd C_bl
Rb_69_65 bit_69_65 bit_69_66 R_bl
Rbb_69_65 bitb_69_65 bitb_69_66 R_bl
Cb_69_65 bit_69_65 gnd C_bl
Cbb_69_65 bitb_69_65 gnd C_bl
Rb_69_66 bit_69_66 bit_69_67 R_bl
Rbb_69_66 bitb_69_66 bitb_69_67 R_bl
Cb_69_66 bit_69_66 gnd C_bl
Cbb_69_66 bitb_69_66 gnd C_bl
Rb_69_67 bit_69_67 bit_69_68 R_bl
Rbb_69_67 bitb_69_67 bitb_69_68 R_bl
Cb_69_67 bit_69_67 gnd C_bl
Cbb_69_67 bitb_69_67 gnd C_bl
Rb_69_68 bit_69_68 bit_69_69 R_bl
Rbb_69_68 bitb_69_68 bitb_69_69 R_bl
Cb_69_68 bit_69_68 gnd C_bl
Cbb_69_68 bitb_69_68 gnd C_bl
Rb_69_69 bit_69_69 bit_69_70 R_bl
Rbb_69_69 bitb_69_69 bitb_69_70 R_bl
Cb_69_69 bit_69_69 gnd C_bl
Cbb_69_69 bitb_69_69 gnd C_bl
Rb_69_70 bit_69_70 bit_69_71 R_bl
Rbb_69_70 bitb_69_70 bitb_69_71 R_bl
Cb_69_70 bit_69_70 gnd C_bl
Cbb_69_70 bitb_69_70 gnd C_bl
Rb_69_71 bit_69_71 bit_69_72 R_bl
Rbb_69_71 bitb_69_71 bitb_69_72 R_bl
Cb_69_71 bit_69_71 gnd C_bl
Cbb_69_71 bitb_69_71 gnd C_bl
Rb_69_72 bit_69_72 bit_69_73 R_bl
Rbb_69_72 bitb_69_72 bitb_69_73 R_bl
Cb_69_72 bit_69_72 gnd C_bl
Cbb_69_72 bitb_69_72 gnd C_bl
Rb_69_73 bit_69_73 bit_69_74 R_bl
Rbb_69_73 bitb_69_73 bitb_69_74 R_bl
Cb_69_73 bit_69_73 gnd C_bl
Cbb_69_73 bitb_69_73 gnd C_bl
Rb_69_74 bit_69_74 bit_69_75 R_bl
Rbb_69_74 bitb_69_74 bitb_69_75 R_bl
Cb_69_74 bit_69_74 gnd C_bl
Cbb_69_74 bitb_69_74 gnd C_bl
Rb_69_75 bit_69_75 bit_69_76 R_bl
Rbb_69_75 bitb_69_75 bitb_69_76 R_bl
Cb_69_75 bit_69_75 gnd C_bl
Cbb_69_75 bitb_69_75 gnd C_bl
Rb_69_76 bit_69_76 bit_69_77 R_bl
Rbb_69_76 bitb_69_76 bitb_69_77 R_bl
Cb_69_76 bit_69_76 gnd C_bl
Cbb_69_76 bitb_69_76 gnd C_bl
Rb_69_77 bit_69_77 bit_69_78 R_bl
Rbb_69_77 bitb_69_77 bitb_69_78 R_bl
Cb_69_77 bit_69_77 gnd C_bl
Cbb_69_77 bitb_69_77 gnd C_bl
Rb_69_78 bit_69_78 bit_69_79 R_bl
Rbb_69_78 bitb_69_78 bitb_69_79 R_bl
Cb_69_78 bit_69_78 gnd C_bl
Cbb_69_78 bitb_69_78 gnd C_bl
Rb_69_79 bit_69_79 bit_69_80 R_bl
Rbb_69_79 bitb_69_79 bitb_69_80 R_bl
Cb_69_79 bit_69_79 gnd C_bl
Cbb_69_79 bitb_69_79 gnd C_bl
Rb_69_80 bit_69_80 bit_69_81 R_bl
Rbb_69_80 bitb_69_80 bitb_69_81 R_bl
Cb_69_80 bit_69_80 gnd C_bl
Cbb_69_80 bitb_69_80 gnd C_bl
Rb_69_81 bit_69_81 bit_69_82 R_bl
Rbb_69_81 bitb_69_81 bitb_69_82 R_bl
Cb_69_81 bit_69_81 gnd C_bl
Cbb_69_81 bitb_69_81 gnd C_bl
Rb_69_82 bit_69_82 bit_69_83 R_bl
Rbb_69_82 bitb_69_82 bitb_69_83 R_bl
Cb_69_82 bit_69_82 gnd C_bl
Cbb_69_82 bitb_69_82 gnd C_bl
Rb_69_83 bit_69_83 bit_69_84 R_bl
Rbb_69_83 bitb_69_83 bitb_69_84 R_bl
Cb_69_83 bit_69_83 gnd C_bl
Cbb_69_83 bitb_69_83 gnd C_bl
Rb_69_84 bit_69_84 bit_69_85 R_bl
Rbb_69_84 bitb_69_84 bitb_69_85 R_bl
Cb_69_84 bit_69_84 gnd C_bl
Cbb_69_84 bitb_69_84 gnd C_bl
Rb_69_85 bit_69_85 bit_69_86 R_bl
Rbb_69_85 bitb_69_85 bitb_69_86 R_bl
Cb_69_85 bit_69_85 gnd C_bl
Cbb_69_85 bitb_69_85 gnd C_bl
Rb_69_86 bit_69_86 bit_69_87 R_bl
Rbb_69_86 bitb_69_86 bitb_69_87 R_bl
Cb_69_86 bit_69_86 gnd C_bl
Cbb_69_86 bitb_69_86 gnd C_bl
Rb_69_87 bit_69_87 bit_69_88 R_bl
Rbb_69_87 bitb_69_87 bitb_69_88 R_bl
Cb_69_87 bit_69_87 gnd C_bl
Cbb_69_87 bitb_69_87 gnd C_bl
Rb_69_88 bit_69_88 bit_69_89 R_bl
Rbb_69_88 bitb_69_88 bitb_69_89 R_bl
Cb_69_88 bit_69_88 gnd C_bl
Cbb_69_88 bitb_69_88 gnd C_bl
Rb_69_89 bit_69_89 bit_69_90 R_bl
Rbb_69_89 bitb_69_89 bitb_69_90 R_bl
Cb_69_89 bit_69_89 gnd C_bl
Cbb_69_89 bitb_69_89 gnd C_bl
Rb_69_90 bit_69_90 bit_69_91 R_bl
Rbb_69_90 bitb_69_90 bitb_69_91 R_bl
Cb_69_90 bit_69_90 gnd C_bl
Cbb_69_90 bitb_69_90 gnd C_bl
Rb_69_91 bit_69_91 bit_69_92 R_bl
Rbb_69_91 bitb_69_91 bitb_69_92 R_bl
Cb_69_91 bit_69_91 gnd C_bl
Cbb_69_91 bitb_69_91 gnd C_bl
Rb_69_92 bit_69_92 bit_69_93 R_bl
Rbb_69_92 bitb_69_92 bitb_69_93 R_bl
Cb_69_92 bit_69_92 gnd C_bl
Cbb_69_92 bitb_69_92 gnd C_bl
Rb_69_93 bit_69_93 bit_69_94 R_bl
Rbb_69_93 bitb_69_93 bitb_69_94 R_bl
Cb_69_93 bit_69_93 gnd C_bl
Cbb_69_93 bitb_69_93 gnd C_bl
Rb_69_94 bit_69_94 bit_69_95 R_bl
Rbb_69_94 bitb_69_94 bitb_69_95 R_bl
Cb_69_94 bit_69_94 gnd C_bl
Cbb_69_94 bitb_69_94 gnd C_bl
Rb_69_95 bit_69_95 bit_69_96 R_bl
Rbb_69_95 bitb_69_95 bitb_69_96 R_bl
Cb_69_95 bit_69_95 gnd C_bl
Cbb_69_95 bitb_69_95 gnd C_bl
Rb_69_96 bit_69_96 bit_69_97 R_bl
Rbb_69_96 bitb_69_96 bitb_69_97 R_bl
Cb_69_96 bit_69_96 gnd C_bl
Cbb_69_96 bitb_69_96 gnd C_bl
Rb_69_97 bit_69_97 bit_69_98 R_bl
Rbb_69_97 bitb_69_97 bitb_69_98 R_bl
Cb_69_97 bit_69_97 gnd C_bl
Cbb_69_97 bitb_69_97 gnd C_bl
Rb_69_98 bit_69_98 bit_69_99 R_bl
Rbb_69_98 bitb_69_98 bitb_69_99 R_bl
Cb_69_98 bit_69_98 gnd C_bl
Cbb_69_98 bitb_69_98 gnd C_bl
Rb_69_99 bit_69_99 bit_69_100 R_bl
Rbb_69_99 bitb_69_99 bitb_69_100 R_bl
Cb_69_99 bit_69_99 gnd C_bl
Cbb_69_99 bitb_69_99 gnd C_bl
Rb_70_0 bit_70_0 bit_70_1 R_bl
Rbb_70_0 bitb_70_0 bitb_70_1 R_bl
Cb_70_0 bit_70_0 gnd C_bl
Cbb_70_0 bitb_70_0 gnd C_bl
Rb_70_1 bit_70_1 bit_70_2 R_bl
Rbb_70_1 bitb_70_1 bitb_70_2 R_bl
Cb_70_1 bit_70_1 gnd C_bl
Cbb_70_1 bitb_70_1 gnd C_bl
Rb_70_2 bit_70_2 bit_70_3 R_bl
Rbb_70_2 bitb_70_2 bitb_70_3 R_bl
Cb_70_2 bit_70_2 gnd C_bl
Cbb_70_2 bitb_70_2 gnd C_bl
Rb_70_3 bit_70_3 bit_70_4 R_bl
Rbb_70_3 bitb_70_3 bitb_70_4 R_bl
Cb_70_3 bit_70_3 gnd C_bl
Cbb_70_3 bitb_70_3 gnd C_bl
Rb_70_4 bit_70_4 bit_70_5 R_bl
Rbb_70_4 bitb_70_4 bitb_70_5 R_bl
Cb_70_4 bit_70_4 gnd C_bl
Cbb_70_4 bitb_70_4 gnd C_bl
Rb_70_5 bit_70_5 bit_70_6 R_bl
Rbb_70_5 bitb_70_5 bitb_70_6 R_bl
Cb_70_5 bit_70_5 gnd C_bl
Cbb_70_5 bitb_70_5 gnd C_bl
Rb_70_6 bit_70_6 bit_70_7 R_bl
Rbb_70_6 bitb_70_6 bitb_70_7 R_bl
Cb_70_6 bit_70_6 gnd C_bl
Cbb_70_6 bitb_70_6 gnd C_bl
Rb_70_7 bit_70_7 bit_70_8 R_bl
Rbb_70_7 bitb_70_7 bitb_70_8 R_bl
Cb_70_7 bit_70_7 gnd C_bl
Cbb_70_7 bitb_70_7 gnd C_bl
Rb_70_8 bit_70_8 bit_70_9 R_bl
Rbb_70_8 bitb_70_8 bitb_70_9 R_bl
Cb_70_8 bit_70_8 gnd C_bl
Cbb_70_8 bitb_70_8 gnd C_bl
Rb_70_9 bit_70_9 bit_70_10 R_bl
Rbb_70_9 bitb_70_9 bitb_70_10 R_bl
Cb_70_9 bit_70_9 gnd C_bl
Cbb_70_9 bitb_70_9 gnd C_bl
Rb_70_10 bit_70_10 bit_70_11 R_bl
Rbb_70_10 bitb_70_10 bitb_70_11 R_bl
Cb_70_10 bit_70_10 gnd C_bl
Cbb_70_10 bitb_70_10 gnd C_bl
Rb_70_11 bit_70_11 bit_70_12 R_bl
Rbb_70_11 bitb_70_11 bitb_70_12 R_bl
Cb_70_11 bit_70_11 gnd C_bl
Cbb_70_11 bitb_70_11 gnd C_bl
Rb_70_12 bit_70_12 bit_70_13 R_bl
Rbb_70_12 bitb_70_12 bitb_70_13 R_bl
Cb_70_12 bit_70_12 gnd C_bl
Cbb_70_12 bitb_70_12 gnd C_bl
Rb_70_13 bit_70_13 bit_70_14 R_bl
Rbb_70_13 bitb_70_13 bitb_70_14 R_bl
Cb_70_13 bit_70_13 gnd C_bl
Cbb_70_13 bitb_70_13 gnd C_bl
Rb_70_14 bit_70_14 bit_70_15 R_bl
Rbb_70_14 bitb_70_14 bitb_70_15 R_bl
Cb_70_14 bit_70_14 gnd C_bl
Cbb_70_14 bitb_70_14 gnd C_bl
Rb_70_15 bit_70_15 bit_70_16 R_bl
Rbb_70_15 bitb_70_15 bitb_70_16 R_bl
Cb_70_15 bit_70_15 gnd C_bl
Cbb_70_15 bitb_70_15 gnd C_bl
Rb_70_16 bit_70_16 bit_70_17 R_bl
Rbb_70_16 bitb_70_16 bitb_70_17 R_bl
Cb_70_16 bit_70_16 gnd C_bl
Cbb_70_16 bitb_70_16 gnd C_bl
Rb_70_17 bit_70_17 bit_70_18 R_bl
Rbb_70_17 bitb_70_17 bitb_70_18 R_bl
Cb_70_17 bit_70_17 gnd C_bl
Cbb_70_17 bitb_70_17 gnd C_bl
Rb_70_18 bit_70_18 bit_70_19 R_bl
Rbb_70_18 bitb_70_18 bitb_70_19 R_bl
Cb_70_18 bit_70_18 gnd C_bl
Cbb_70_18 bitb_70_18 gnd C_bl
Rb_70_19 bit_70_19 bit_70_20 R_bl
Rbb_70_19 bitb_70_19 bitb_70_20 R_bl
Cb_70_19 bit_70_19 gnd C_bl
Cbb_70_19 bitb_70_19 gnd C_bl
Rb_70_20 bit_70_20 bit_70_21 R_bl
Rbb_70_20 bitb_70_20 bitb_70_21 R_bl
Cb_70_20 bit_70_20 gnd C_bl
Cbb_70_20 bitb_70_20 gnd C_bl
Rb_70_21 bit_70_21 bit_70_22 R_bl
Rbb_70_21 bitb_70_21 bitb_70_22 R_bl
Cb_70_21 bit_70_21 gnd C_bl
Cbb_70_21 bitb_70_21 gnd C_bl
Rb_70_22 bit_70_22 bit_70_23 R_bl
Rbb_70_22 bitb_70_22 bitb_70_23 R_bl
Cb_70_22 bit_70_22 gnd C_bl
Cbb_70_22 bitb_70_22 gnd C_bl
Rb_70_23 bit_70_23 bit_70_24 R_bl
Rbb_70_23 bitb_70_23 bitb_70_24 R_bl
Cb_70_23 bit_70_23 gnd C_bl
Cbb_70_23 bitb_70_23 gnd C_bl
Rb_70_24 bit_70_24 bit_70_25 R_bl
Rbb_70_24 bitb_70_24 bitb_70_25 R_bl
Cb_70_24 bit_70_24 gnd C_bl
Cbb_70_24 bitb_70_24 gnd C_bl
Rb_70_25 bit_70_25 bit_70_26 R_bl
Rbb_70_25 bitb_70_25 bitb_70_26 R_bl
Cb_70_25 bit_70_25 gnd C_bl
Cbb_70_25 bitb_70_25 gnd C_bl
Rb_70_26 bit_70_26 bit_70_27 R_bl
Rbb_70_26 bitb_70_26 bitb_70_27 R_bl
Cb_70_26 bit_70_26 gnd C_bl
Cbb_70_26 bitb_70_26 gnd C_bl
Rb_70_27 bit_70_27 bit_70_28 R_bl
Rbb_70_27 bitb_70_27 bitb_70_28 R_bl
Cb_70_27 bit_70_27 gnd C_bl
Cbb_70_27 bitb_70_27 gnd C_bl
Rb_70_28 bit_70_28 bit_70_29 R_bl
Rbb_70_28 bitb_70_28 bitb_70_29 R_bl
Cb_70_28 bit_70_28 gnd C_bl
Cbb_70_28 bitb_70_28 gnd C_bl
Rb_70_29 bit_70_29 bit_70_30 R_bl
Rbb_70_29 bitb_70_29 bitb_70_30 R_bl
Cb_70_29 bit_70_29 gnd C_bl
Cbb_70_29 bitb_70_29 gnd C_bl
Rb_70_30 bit_70_30 bit_70_31 R_bl
Rbb_70_30 bitb_70_30 bitb_70_31 R_bl
Cb_70_30 bit_70_30 gnd C_bl
Cbb_70_30 bitb_70_30 gnd C_bl
Rb_70_31 bit_70_31 bit_70_32 R_bl
Rbb_70_31 bitb_70_31 bitb_70_32 R_bl
Cb_70_31 bit_70_31 gnd C_bl
Cbb_70_31 bitb_70_31 gnd C_bl
Rb_70_32 bit_70_32 bit_70_33 R_bl
Rbb_70_32 bitb_70_32 bitb_70_33 R_bl
Cb_70_32 bit_70_32 gnd C_bl
Cbb_70_32 bitb_70_32 gnd C_bl
Rb_70_33 bit_70_33 bit_70_34 R_bl
Rbb_70_33 bitb_70_33 bitb_70_34 R_bl
Cb_70_33 bit_70_33 gnd C_bl
Cbb_70_33 bitb_70_33 gnd C_bl
Rb_70_34 bit_70_34 bit_70_35 R_bl
Rbb_70_34 bitb_70_34 bitb_70_35 R_bl
Cb_70_34 bit_70_34 gnd C_bl
Cbb_70_34 bitb_70_34 gnd C_bl
Rb_70_35 bit_70_35 bit_70_36 R_bl
Rbb_70_35 bitb_70_35 bitb_70_36 R_bl
Cb_70_35 bit_70_35 gnd C_bl
Cbb_70_35 bitb_70_35 gnd C_bl
Rb_70_36 bit_70_36 bit_70_37 R_bl
Rbb_70_36 bitb_70_36 bitb_70_37 R_bl
Cb_70_36 bit_70_36 gnd C_bl
Cbb_70_36 bitb_70_36 gnd C_bl
Rb_70_37 bit_70_37 bit_70_38 R_bl
Rbb_70_37 bitb_70_37 bitb_70_38 R_bl
Cb_70_37 bit_70_37 gnd C_bl
Cbb_70_37 bitb_70_37 gnd C_bl
Rb_70_38 bit_70_38 bit_70_39 R_bl
Rbb_70_38 bitb_70_38 bitb_70_39 R_bl
Cb_70_38 bit_70_38 gnd C_bl
Cbb_70_38 bitb_70_38 gnd C_bl
Rb_70_39 bit_70_39 bit_70_40 R_bl
Rbb_70_39 bitb_70_39 bitb_70_40 R_bl
Cb_70_39 bit_70_39 gnd C_bl
Cbb_70_39 bitb_70_39 gnd C_bl
Rb_70_40 bit_70_40 bit_70_41 R_bl
Rbb_70_40 bitb_70_40 bitb_70_41 R_bl
Cb_70_40 bit_70_40 gnd C_bl
Cbb_70_40 bitb_70_40 gnd C_bl
Rb_70_41 bit_70_41 bit_70_42 R_bl
Rbb_70_41 bitb_70_41 bitb_70_42 R_bl
Cb_70_41 bit_70_41 gnd C_bl
Cbb_70_41 bitb_70_41 gnd C_bl
Rb_70_42 bit_70_42 bit_70_43 R_bl
Rbb_70_42 bitb_70_42 bitb_70_43 R_bl
Cb_70_42 bit_70_42 gnd C_bl
Cbb_70_42 bitb_70_42 gnd C_bl
Rb_70_43 bit_70_43 bit_70_44 R_bl
Rbb_70_43 bitb_70_43 bitb_70_44 R_bl
Cb_70_43 bit_70_43 gnd C_bl
Cbb_70_43 bitb_70_43 gnd C_bl
Rb_70_44 bit_70_44 bit_70_45 R_bl
Rbb_70_44 bitb_70_44 bitb_70_45 R_bl
Cb_70_44 bit_70_44 gnd C_bl
Cbb_70_44 bitb_70_44 gnd C_bl
Rb_70_45 bit_70_45 bit_70_46 R_bl
Rbb_70_45 bitb_70_45 bitb_70_46 R_bl
Cb_70_45 bit_70_45 gnd C_bl
Cbb_70_45 bitb_70_45 gnd C_bl
Rb_70_46 bit_70_46 bit_70_47 R_bl
Rbb_70_46 bitb_70_46 bitb_70_47 R_bl
Cb_70_46 bit_70_46 gnd C_bl
Cbb_70_46 bitb_70_46 gnd C_bl
Rb_70_47 bit_70_47 bit_70_48 R_bl
Rbb_70_47 bitb_70_47 bitb_70_48 R_bl
Cb_70_47 bit_70_47 gnd C_bl
Cbb_70_47 bitb_70_47 gnd C_bl
Rb_70_48 bit_70_48 bit_70_49 R_bl
Rbb_70_48 bitb_70_48 bitb_70_49 R_bl
Cb_70_48 bit_70_48 gnd C_bl
Cbb_70_48 bitb_70_48 gnd C_bl
Rb_70_49 bit_70_49 bit_70_50 R_bl
Rbb_70_49 bitb_70_49 bitb_70_50 R_bl
Cb_70_49 bit_70_49 gnd C_bl
Cbb_70_49 bitb_70_49 gnd C_bl
Rb_70_50 bit_70_50 bit_70_51 R_bl
Rbb_70_50 bitb_70_50 bitb_70_51 R_bl
Cb_70_50 bit_70_50 gnd C_bl
Cbb_70_50 bitb_70_50 gnd C_bl
Rb_70_51 bit_70_51 bit_70_52 R_bl
Rbb_70_51 bitb_70_51 bitb_70_52 R_bl
Cb_70_51 bit_70_51 gnd C_bl
Cbb_70_51 bitb_70_51 gnd C_bl
Rb_70_52 bit_70_52 bit_70_53 R_bl
Rbb_70_52 bitb_70_52 bitb_70_53 R_bl
Cb_70_52 bit_70_52 gnd C_bl
Cbb_70_52 bitb_70_52 gnd C_bl
Rb_70_53 bit_70_53 bit_70_54 R_bl
Rbb_70_53 bitb_70_53 bitb_70_54 R_bl
Cb_70_53 bit_70_53 gnd C_bl
Cbb_70_53 bitb_70_53 gnd C_bl
Rb_70_54 bit_70_54 bit_70_55 R_bl
Rbb_70_54 bitb_70_54 bitb_70_55 R_bl
Cb_70_54 bit_70_54 gnd C_bl
Cbb_70_54 bitb_70_54 gnd C_bl
Rb_70_55 bit_70_55 bit_70_56 R_bl
Rbb_70_55 bitb_70_55 bitb_70_56 R_bl
Cb_70_55 bit_70_55 gnd C_bl
Cbb_70_55 bitb_70_55 gnd C_bl
Rb_70_56 bit_70_56 bit_70_57 R_bl
Rbb_70_56 bitb_70_56 bitb_70_57 R_bl
Cb_70_56 bit_70_56 gnd C_bl
Cbb_70_56 bitb_70_56 gnd C_bl
Rb_70_57 bit_70_57 bit_70_58 R_bl
Rbb_70_57 bitb_70_57 bitb_70_58 R_bl
Cb_70_57 bit_70_57 gnd C_bl
Cbb_70_57 bitb_70_57 gnd C_bl
Rb_70_58 bit_70_58 bit_70_59 R_bl
Rbb_70_58 bitb_70_58 bitb_70_59 R_bl
Cb_70_58 bit_70_58 gnd C_bl
Cbb_70_58 bitb_70_58 gnd C_bl
Rb_70_59 bit_70_59 bit_70_60 R_bl
Rbb_70_59 bitb_70_59 bitb_70_60 R_bl
Cb_70_59 bit_70_59 gnd C_bl
Cbb_70_59 bitb_70_59 gnd C_bl
Rb_70_60 bit_70_60 bit_70_61 R_bl
Rbb_70_60 bitb_70_60 bitb_70_61 R_bl
Cb_70_60 bit_70_60 gnd C_bl
Cbb_70_60 bitb_70_60 gnd C_bl
Rb_70_61 bit_70_61 bit_70_62 R_bl
Rbb_70_61 bitb_70_61 bitb_70_62 R_bl
Cb_70_61 bit_70_61 gnd C_bl
Cbb_70_61 bitb_70_61 gnd C_bl
Rb_70_62 bit_70_62 bit_70_63 R_bl
Rbb_70_62 bitb_70_62 bitb_70_63 R_bl
Cb_70_62 bit_70_62 gnd C_bl
Cbb_70_62 bitb_70_62 gnd C_bl
Rb_70_63 bit_70_63 bit_70_64 R_bl
Rbb_70_63 bitb_70_63 bitb_70_64 R_bl
Cb_70_63 bit_70_63 gnd C_bl
Cbb_70_63 bitb_70_63 gnd C_bl
Rb_70_64 bit_70_64 bit_70_65 R_bl
Rbb_70_64 bitb_70_64 bitb_70_65 R_bl
Cb_70_64 bit_70_64 gnd C_bl
Cbb_70_64 bitb_70_64 gnd C_bl
Rb_70_65 bit_70_65 bit_70_66 R_bl
Rbb_70_65 bitb_70_65 bitb_70_66 R_bl
Cb_70_65 bit_70_65 gnd C_bl
Cbb_70_65 bitb_70_65 gnd C_bl
Rb_70_66 bit_70_66 bit_70_67 R_bl
Rbb_70_66 bitb_70_66 bitb_70_67 R_bl
Cb_70_66 bit_70_66 gnd C_bl
Cbb_70_66 bitb_70_66 gnd C_bl
Rb_70_67 bit_70_67 bit_70_68 R_bl
Rbb_70_67 bitb_70_67 bitb_70_68 R_bl
Cb_70_67 bit_70_67 gnd C_bl
Cbb_70_67 bitb_70_67 gnd C_bl
Rb_70_68 bit_70_68 bit_70_69 R_bl
Rbb_70_68 bitb_70_68 bitb_70_69 R_bl
Cb_70_68 bit_70_68 gnd C_bl
Cbb_70_68 bitb_70_68 gnd C_bl
Rb_70_69 bit_70_69 bit_70_70 R_bl
Rbb_70_69 bitb_70_69 bitb_70_70 R_bl
Cb_70_69 bit_70_69 gnd C_bl
Cbb_70_69 bitb_70_69 gnd C_bl
Rb_70_70 bit_70_70 bit_70_71 R_bl
Rbb_70_70 bitb_70_70 bitb_70_71 R_bl
Cb_70_70 bit_70_70 gnd C_bl
Cbb_70_70 bitb_70_70 gnd C_bl
Rb_70_71 bit_70_71 bit_70_72 R_bl
Rbb_70_71 bitb_70_71 bitb_70_72 R_bl
Cb_70_71 bit_70_71 gnd C_bl
Cbb_70_71 bitb_70_71 gnd C_bl
Rb_70_72 bit_70_72 bit_70_73 R_bl
Rbb_70_72 bitb_70_72 bitb_70_73 R_bl
Cb_70_72 bit_70_72 gnd C_bl
Cbb_70_72 bitb_70_72 gnd C_bl
Rb_70_73 bit_70_73 bit_70_74 R_bl
Rbb_70_73 bitb_70_73 bitb_70_74 R_bl
Cb_70_73 bit_70_73 gnd C_bl
Cbb_70_73 bitb_70_73 gnd C_bl
Rb_70_74 bit_70_74 bit_70_75 R_bl
Rbb_70_74 bitb_70_74 bitb_70_75 R_bl
Cb_70_74 bit_70_74 gnd C_bl
Cbb_70_74 bitb_70_74 gnd C_bl
Rb_70_75 bit_70_75 bit_70_76 R_bl
Rbb_70_75 bitb_70_75 bitb_70_76 R_bl
Cb_70_75 bit_70_75 gnd C_bl
Cbb_70_75 bitb_70_75 gnd C_bl
Rb_70_76 bit_70_76 bit_70_77 R_bl
Rbb_70_76 bitb_70_76 bitb_70_77 R_bl
Cb_70_76 bit_70_76 gnd C_bl
Cbb_70_76 bitb_70_76 gnd C_bl
Rb_70_77 bit_70_77 bit_70_78 R_bl
Rbb_70_77 bitb_70_77 bitb_70_78 R_bl
Cb_70_77 bit_70_77 gnd C_bl
Cbb_70_77 bitb_70_77 gnd C_bl
Rb_70_78 bit_70_78 bit_70_79 R_bl
Rbb_70_78 bitb_70_78 bitb_70_79 R_bl
Cb_70_78 bit_70_78 gnd C_bl
Cbb_70_78 bitb_70_78 gnd C_bl
Rb_70_79 bit_70_79 bit_70_80 R_bl
Rbb_70_79 bitb_70_79 bitb_70_80 R_bl
Cb_70_79 bit_70_79 gnd C_bl
Cbb_70_79 bitb_70_79 gnd C_bl
Rb_70_80 bit_70_80 bit_70_81 R_bl
Rbb_70_80 bitb_70_80 bitb_70_81 R_bl
Cb_70_80 bit_70_80 gnd C_bl
Cbb_70_80 bitb_70_80 gnd C_bl
Rb_70_81 bit_70_81 bit_70_82 R_bl
Rbb_70_81 bitb_70_81 bitb_70_82 R_bl
Cb_70_81 bit_70_81 gnd C_bl
Cbb_70_81 bitb_70_81 gnd C_bl
Rb_70_82 bit_70_82 bit_70_83 R_bl
Rbb_70_82 bitb_70_82 bitb_70_83 R_bl
Cb_70_82 bit_70_82 gnd C_bl
Cbb_70_82 bitb_70_82 gnd C_bl
Rb_70_83 bit_70_83 bit_70_84 R_bl
Rbb_70_83 bitb_70_83 bitb_70_84 R_bl
Cb_70_83 bit_70_83 gnd C_bl
Cbb_70_83 bitb_70_83 gnd C_bl
Rb_70_84 bit_70_84 bit_70_85 R_bl
Rbb_70_84 bitb_70_84 bitb_70_85 R_bl
Cb_70_84 bit_70_84 gnd C_bl
Cbb_70_84 bitb_70_84 gnd C_bl
Rb_70_85 bit_70_85 bit_70_86 R_bl
Rbb_70_85 bitb_70_85 bitb_70_86 R_bl
Cb_70_85 bit_70_85 gnd C_bl
Cbb_70_85 bitb_70_85 gnd C_bl
Rb_70_86 bit_70_86 bit_70_87 R_bl
Rbb_70_86 bitb_70_86 bitb_70_87 R_bl
Cb_70_86 bit_70_86 gnd C_bl
Cbb_70_86 bitb_70_86 gnd C_bl
Rb_70_87 bit_70_87 bit_70_88 R_bl
Rbb_70_87 bitb_70_87 bitb_70_88 R_bl
Cb_70_87 bit_70_87 gnd C_bl
Cbb_70_87 bitb_70_87 gnd C_bl
Rb_70_88 bit_70_88 bit_70_89 R_bl
Rbb_70_88 bitb_70_88 bitb_70_89 R_bl
Cb_70_88 bit_70_88 gnd C_bl
Cbb_70_88 bitb_70_88 gnd C_bl
Rb_70_89 bit_70_89 bit_70_90 R_bl
Rbb_70_89 bitb_70_89 bitb_70_90 R_bl
Cb_70_89 bit_70_89 gnd C_bl
Cbb_70_89 bitb_70_89 gnd C_bl
Rb_70_90 bit_70_90 bit_70_91 R_bl
Rbb_70_90 bitb_70_90 bitb_70_91 R_bl
Cb_70_90 bit_70_90 gnd C_bl
Cbb_70_90 bitb_70_90 gnd C_bl
Rb_70_91 bit_70_91 bit_70_92 R_bl
Rbb_70_91 bitb_70_91 bitb_70_92 R_bl
Cb_70_91 bit_70_91 gnd C_bl
Cbb_70_91 bitb_70_91 gnd C_bl
Rb_70_92 bit_70_92 bit_70_93 R_bl
Rbb_70_92 bitb_70_92 bitb_70_93 R_bl
Cb_70_92 bit_70_92 gnd C_bl
Cbb_70_92 bitb_70_92 gnd C_bl
Rb_70_93 bit_70_93 bit_70_94 R_bl
Rbb_70_93 bitb_70_93 bitb_70_94 R_bl
Cb_70_93 bit_70_93 gnd C_bl
Cbb_70_93 bitb_70_93 gnd C_bl
Rb_70_94 bit_70_94 bit_70_95 R_bl
Rbb_70_94 bitb_70_94 bitb_70_95 R_bl
Cb_70_94 bit_70_94 gnd C_bl
Cbb_70_94 bitb_70_94 gnd C_bl
Rb_70_95 bit_70_95 bit_70_96 R_bl
Rbb_70_95 bitb_70_95 bitb_70_96 R_bl
Cb_70_95 bit_70_95 gnd C_bl
Cbb_70_95 bitb_70_95 gnd C_bl
Rb_70_96 bit_70_96 bit_70_97 R_bl
Rbb_70_96 bitb_70_96 bitb_70_97 R_bl
Cb_70_96 bit_70_96 gnd C_bl
Cbb_70_96 bitb_70_96 gnd C_bl
Rb_70_97 bit_70_97 bit_70_98 R_bl
Rbb_70_97 bitb_70_97 bitb_70_98 R_bl
Cb_70_97 bit_70_97 gnd C_bl
Cbb_70_97 bitb_70_97 gnd C_bl
Rb_70_98 bit_70_98 bit_70_99 R_bl
Rbb_70_98 bitb_70_98 bitb_70_99 R_bl
Cb_70_98 bit_70_98 gnd C_bl
Cbb_70_98 bitb_70_98 gnd C_bl
Rb_70_99 bit_70_99 bit_70_100 R_bl
Rbb_70_99 bitb_70_99 bitb_70_100 R_bl
Cb_70_99 bit_70_99 gnd C_bl
Cbb_70_99 bitb_70_99 gnd C_bl
Rb_71_0 bit_71_0 bit_71_1 R_bl
Rbb_71_0 bitb_71_0 bitb_71_1 R_bl
Cb_71_0 bit_71_0 gnd C_bl
Cbb_71_0 bitb_71_0 gnd C_bl
Rb_71_1 bit_71_1 bit_71_2 R_bl
Rbb_71_1 bitb_71_1 bitb_71_2 R_bl
Cb_71_1 bit_71_1 gnd C_bl
Cbb_71_1 bitb_71_1 gnd C_bl
Rb_71_2 bit_71_2 bit_71_3 R_bl
Rbb_71_2 bitb_71_2 bitb_71_3 R_bl
Cb_71_2 bit_71_2 gnd C_bl
Cbb_71_2 bitb_71_2 gnd C_bl
Rb_71_3 bit_71_3 bit_71_4 R_bl
Rbb_71_3 bitb_71_3 bitb_71_4 R_bl
Cb_71_3 bit_71_3 gnd C_bl
Cbb_71_3 bitb_71_3 gnd C_bl
Rb_71_4 bit_71_4 bit_71_5 R_bl
Rbb_71_4 bitb_71_4 bitb_71_5 R_bl
Cb_71_4 bit_71_4 gnd C_bl
Cbb_71_4 bitb_71_4 gnd C_bl
Rb_71_5 bit_71_5 bit_71_6 R_bl
Rbb_71_5 bitb_71_5 bitb_71_6 R_bl
Cb_71_5 bit_71_5 gnd C_bl
Cbb_71_5 bitb_71_5 gnd C_bl
Rb_71_6 bit_71_6 bit_71_7 R_bl
Rbb_71_6 bitb_71_6 bitb_71_7 R_bl
Cb_71_6 bit_71_6 gnd C_bl
Cbb_71_6 bitb_71_6 gnd C_bl
Rb_71_7 bit_71_7 bit_71_8 R_bl
Rbb_71_7 bitb_71_7 bitb_71_8 R_bl
Cb_71_7 bit_71_7 gnd C_bl
Cbb_71_7 bitb_71_7 gnd C_bl
Rb_71_8 bit_71_8 bit_71_9 R_bl
Rbb_71_8 bitb_71_8 bitb_71_9 R_bl
Cb_71_8 bit_71_8 gnd C_bl
Cbb_71_8 bitb_71_8 gnd C_bl
Rb_71_9 bit_71_9 bit_71_10 R_bl
Rbb_71_9 bitb_71_9 bitb_71_10 R_bl
Cb_71_9 bit_71_9 gnd C_bl
Cbb_71_9 bitb_71_9 gnd C_bl
Rb_71_10 bit_71_10 bit_71_11 R_bl
Rbb_71_10 bitb_71_10 bitb_71_11 R_bl
Cb_71_10 bit_71_10 gnd C_bl
Cbb_71_10 bitb_71_10 gnd C_bl
Rb_71_11 bit_71_11 bit_71_12 R_bl
Rbb_71_11 bitb_71_11 bitb_71_12 R_bl
Cb_71_11 bit_71_11 gnd C_bl
Cbb_71_11 bitb_71_11 gnd C_bl
Rb_71_12 bit_71_12 bit_71_13 R_bl
Rbb_71_12 bitb_71_12 bitb_71_13 R_bl
Cb_71_12 bit_71_12 gnd C_bl
Cbb_71_12 bitb_71_12 gnd C_bl
Rb_71_13 bit_71_13 bit_71_14 R_bl
Rbb_71_13 bitb_71_13 bitb_71_14 R_bl
Cb_71_13 bit_71_13 gnd C_bl
Cbb_71_13 bitb_71_13 gnd C_bl
Rb_71_14 bit_71_14 bit_71_15 R_bl
Rbb_71_14 bitb_71_14 bitb_71_15 R_bl
Cb_71_14 bit_71_14 gnd C_bl
Cbb_71_14 bitb_71_14 gnd C_bl
Rb_71_15 bit_71_15 bit_71_16 R_bl
Rbb_71_15 bitb_71_15 bitb_71_16 R_bl
Cb_71_15 bit_71_15 gnd C_bl
Cbb_71_15 bitb_71_15 gnd C_bl
Rb_71_16 bit_71_16 bit_71_17 R_bl
Rbb_71_16 bitb_71_16 bitb_71_17 R_bl
Cb_71_16 bit_71_16 gnd C_bl
Cbb_71_16 bitb_71_16 gnd C_bl
Rb_71_17 bit_71_17 bit_71_18 R_bl
Rbb_71_17 bitb_71_17 bitb_71_18 R_bl
Cb_71_17 bit_71_17 gnd C_bl
Cbb_71_17 bitb_71_17 gnd C_bl
Rb_71_18 bit_71_18 bit_71_19 R_bl
Rbb_71_18 bitb_71_18 bitb_71_19 R_bl
Cb_71_18 bit_71_18 gnd C_bl
Cbb_71_18 bitb_71_18 gnd C_bl
Rb_71_19 bit_71_19 bit_71_20 R_bl
Rbb_71_19 bitb_71_19 bitb_71_20 R_bl
Cb_71_19 bit_71_19 gnd C_bl
Cbb_71_19 bitb_71_19 gnd C_bl
Rb_71_20 bit_71_20 bit_71_21 R_bl
Rbb_71_20 bitb_71_20 bitb_71_21 R_bl
Cb_71_20 bit_71_20 gnd C_bl
Cbb_71_20 bitb_71_20 gnd C_bl
Rb_71_21 bit_71_21 bit_71_22 R_bl
Rbb_71_21 bitb_71_21 bitb_71_22 R_bl
Cb_71_21 bit_71_21 gnd C_bl
Cbb_71_21 bitb_71_21 gnd C_bl
Rb_71_22 bit_71_22 bit_71_23 R_bl
Rbb_71_22 bitb_71_22 bitb_71_23 R_bl
Cb_71_22 bit_71_22 gnd C_bl
Cbb_71_22 bitb_71_22 gnd C_bl
Rb_71_23 bit_71_23 bit_71_24 R_bl
Rbb_71_23 bitb_71_23 bitb_71_24 R_bl
Cb_71_23 bit_71_23 gnd C_bl
Cbb_71_23 bitb_71_23 gnd C_bl
Rb_71_24 bit_71_24 bit_71_25 R_bl
Rbb_71_24 bitb_71_24 bitb_71_25 R_bl
Cb_71_24 bit_71_24 gnd C_bl
Cbb_71_24 bitb_71_24 gnd C_bl
Rb_71_25 bit_71_25 bit_71_26 R_bl
Rbb_71_25 bitb_71_25 bitb_71_26 R_bl
Cb_71_25 bit_71_25 gnd C_bl
Cbb_71_25 bitb_71_25 gnd C_bl
Rb_71_26 bit_71_26 bit_71_27 R_bl
Rbb_71_26 bitb_71_26 bitb_71_27 R_bl
Cb_71_26 bit_71_26 gnd C_bl
Cbb_71_26 bitb_71_26 gnd C_bl
Rb_71_27 bit_71_27 bit_71_28 R_bl
Rbb_71_27 bitb_71_27 bitb_71_28 R_bl
Cb_71_27 bit_71_27 gnd C_bl
Cbb_71_27 bitb_71_27 gnd C_bl
Rb_71_28 bit_71_28 bit_71_29 R_bl
Rbb_71_28 bitb_71_28 bitb_71_29 R_bl
Cb_71_28 bit_71_28 gnd C_bl
Cbb_71_28 bitb_71_28 gnd C_bl
Rb_71_29 bit_71_29 bit_71_30 R_bl
Rbb_71_29 bitb_71_29 bitb_71_30 R_bl
Cb_71_29 bit_71_29 gnd C_bl
Cbb_71_29 bitb_71_29 gnd C_bl
Rb_71_30 bit_71_30 bit_71_31 R_bl
Rbb_71_30 bitb_71_30 bitb_71_31 R_bl
Cb_71_30 bit_71_30 gnd C_bl
Cbb_71_30 bitb_71_30 gnd C_bl
Rb_71_31 bit_71_31 bit_71_32 R_bl
Rbb_71_31 bitb_71_31 bitb_71_32 R_bl
Cb_71_31 bit_71_31 gnd C_bl
Cbb_71_31 bitb_71_31 gnd C_bl
Rb_71_32 bit_71_32 bit_71_33 R_bl
Rbb_71_32 bitb_71_32 bitb_71_33 R_bl
Cb_71_32 bit_71_32 gnd C_bl
Cbb_71_32 bitb_71_32 gnd C_bl
Rb_71_33 bit_71_33 bit_71_34 R_bl
Rbb_71_33 bitb_71_33 bitb_71_34 R_bl
Cb_71_33 bit_71_33 gnd C_bl
Cbb_71_33 bitb_71_33 gnd C_bl
Rb_71_34 bit_71_34 bit_71_35 R_bl
Rbb_71_34 bitb_71_34 bitb_71_35 R_bl
Cb_71_34 bit_71_34 gnd C_bl
Cbb_71_34 bitb_71_34 gnd C_bl
Rb_71_35 bit_71_35 bit_71_36 R_bl
Rbb_71_35 bitb_71_35 bitb_71_36 R_bl
Cb_71_35 bit_71_35 gnd C_bl
Cbb_71_35 bitb_71_35 gnd C_bl
Rb_71_36 bit_71_36 bit_71_37 R_bl
Rbb_71_36 bitb_71_36 bitb_71_37 R_bl
Cb_71_36 bit_71_36 gnd C_bl
Cbb_71_36 bitb_71_36 gnd C_bl
Rb_71_37 bit_71_37 bit_71_38 R_bl
Rbb_71_37 bitb_71_37 bitb_71_38 R_bl
Cb_71_37 bit_71_37 gnd C_bl
Cbb_71_37 bitb_71_37 gnd C_bl
Rb_71_38 bit_71_38 bit_71_39 R_bl
Rbb_71_38 bitb_71_38 bitb_71_39 R_bl
Cb_71_38 bit_71_38 gnd C_bl
Cbb_71_38 bitb_71_38 gnd C_bl
Rb_71_39 bit_71_39 bit_71_40 R_bl
Rbb_71_39 bitb_71_39 bitb_71_40 R_bl
Cb_71_39 bit_71_39 gnd C_bl
Cbb_71_39 bitb_71_39 gnd C_bl
Rb_71_40 bit_71_40 bit_71_41 R_bl
Rbb_71_40 bitb_71_40 bitb_71_41 R_bl
Cb_71_40 bit_71_40 gnd C_bl
Cbb_71_40 bitb_71_40 gnd C_bl
Rb_71_41 bit_71_41 bit_71_42 R_bl
Rbb_71_41 bitb_71_41 bitb_71_42 R_bl
Cb_71_41 bit_71_41 gnd C_bl
Cbb_71_41 bitb_71_41 gnd C_bl
Rb_71_42 bit_71_42 bit_71_43 R_bl
Rbb_71_42 bitb_71_42 bitb_71_43 R_bl
Cb_71_42 bit_71_42 gnd C_bl
Cbb_71_42 bitb_71_42 gnd C_bl
Rb_71_43 bit_71_43 bit_71_44 R_bl
Rbb_71_43 bitb_71_43 bitb_71_44 R_bl
Cb_71_43 bit_71_43 gnd C_bl
Cbb_71_43 bitb_71_43 gnd C_bl
Rb_71_44 bit_71_44 bit_71_45 R_bl
Rbb_71_44 bitb_71_44 bitb_71_45 R_bl
Cb_71_44 bit_71_44 gnd C_bl
Cbb_71_44 bitb_71_44 gnd C_bl
Rb_71_45 bit_71_45 bit_71_46 R_bl
Rbb_71_45 bitb_71_45 bitb_71_46 R_bl
Cb_71_45 bit_71_45 gnd C_bl
Cbb_71_45 bitb_71_45 gnd C_bl
Rb_71_46 bit_71_46 bit_71_47 R_bl
Rbb_71_46 bitb_71_46 bitb_71_47 R_bl
Cb_71_46 bit_71_46 gnd C_bl
Cbb_71_46 bitb_71_46 gnd C_bl
Rb_71_47 bit_71_47 bit_71_48 R_bl
Rbb_71_47 bitb_71_47 bitb_71_48 R_bl
Cb_71_47 bit_71_47 gnd C_bl
Cbb_71_47 bitb_71_47 gnd C_bl
Rb_71_48 bit_71_48 bit_71_49 R_bl
Rbb_71_48 bitb_71_48 bitb_71_49 R_bl
Cb_71_48 bit_71_48 gnd C_bl
Cbb_71_48 bitb_71_48 gnd C_bl
Rb_71_49 bit_71_49 bit_71_50 R_bl
Rbb_71_49 bitb_71_49 bitb_71_50 R_bl
Cb_71_49 bit_71_49 gnd C_bl
Cbb_71_49 bitb_71_49 gnd C_bl
Rb_71_50 bit_71_50 bit_71_51 R_bl
Rbb_71_50 bitb_71_50 bitb_71_51 R_bl
Cb_71_50 bit_71_50 gnd C_bl
Cbb_71_50 bitb_71_50 gnd C_bl
Rb_71_51 bit_71_51 bit_71_52 R_bl
Rbb_71_51 bitb_71_51 bitb_71_52 R_bl
Cb_71_51 bit_71_51 gnd C_bl
Cbb_71_51 bitb_71_51 gnd C_bl
Rb_71_52 bit_71_52 bit_71_53 R_bl
Rbb_71_52 bitb_71_52 bitb_71_53 R_bl
Cb_71_52 bit_71_52 gnd C_bl
Cbb_71_52 bitb_71_52 gnd C_bl
Rb_71_53 bit_71_53 bit_71_54 R_bl
Rbb_71_53 bitb_71_53 bitb_71_54 R_bl
Cb_71_53 bit_71_53 gnd C_bl
Cbb_71_53 bitb_71_53 gnd C_bl
Rb_71_54 bit_71_54 bit_71_55 R_bl
Rbb_71_54 bitb_71_54 bitb_71_55 R_bl
Cb_71_54 bit_71_54 gnd C_bl
Cbb_71_54 bitb_71_54 gnd C_bl
Rb_71_55 bit_71_55 bit_71_56 R_bl
Rbb_71_55 bitb_71_55 bitb_71_56 R_bl
Cb_71_55 bit_71_55 gnd C_bl
Cbb_71_55 bitb_71_55 gnd C_bl
Rb_71_56 bit_71_56 bit_71_57 R_bl
Rbb_71_56 bitb_71_56 bitb_71_57 R_bl
Cb_71_56 bit_71_56 gnd C_bl
Cbb_71_56 bitb_71_56 gnd C_bl
Rb_71_57 bit_71_57 bit_71_58 R_bl
Rbb_71_57 bitb_71_57 bitb_71_58 R_bl
Cb_71_57 bit_71_57 gnd C_bl
Cbb_71_57 bitb_71_57 gnd C_bl
Rb_71_58 bit_71_58 bit_71_59 R_bl
Rbb_71_58 bitb_71_58 bitb_71_59 R_bl
Cb_71_58 bit_71_58 gnd C_bl
Cbb_71_58 bitb_71_58 gnd C_bl
Rb_71_59 bit_71_59 bit_71_60 R_bl
Rbb_71_59 bitb_71_59 bitb_71_60 R_bl
Cb_71_59 bit_71_59 gnd C_bl
Cbb_71_59 bitb_71_59 gnd C_bl
Rb_71_60 bit_71_60 bit_71_61 R_bl
Rbb_71_60 bitb_71_60 bitb_71_61 R_bl
Cb_71_60 bit_71_60 gnd C_bl
Cbb_71_60 bitb_71_60 gnd C_bl
Rb_71_61 bit_71_61 bit_71_62 R_bl
Rbb_71_61 bitb_71_61 bitb_71_62 R_bl
Cb_71_61 bit_71_61 gnd C_bl
Cbb_71_61 bitb_71_61 gnd C_bl
Rb_71_62 bit_71_62 bit_71_63 R_bl
Rbb_71_62 bitb_71_62 bitb_71_63 R_bl
Cb_71_62 bit_71_62 gnd C_bl
Cbb_71_62 bitb_71_62 gnd C_bl
Rb_71_63 bit_71_63 bit_71_64 R_bl
Rbb_71_63 bitb_71_63 bitb_71_64 R_bl
Cb_71_63 bit_71_63 gnd C_bl
Cbb_71_63 bitb_71_63 gnd C_bl
Rb_71_64 bit_71_64 bit_71_65 R_bl
Rbb_71_64 bitb_71_64 bitb_71_65 R_bl
Cb_71_64 bit_71_64 gnd C_bl
Cbb_71_64 bitb_71_64 gnd C_bl
Rb_71_65 bit_71_65 bit_71_66 R_bl
Rbb_71_65 bitb_71_65 bitb_71_66 R_bl
Cb_71_65 bit_71_65 gnd C_bl
Cbb_71_65 bitb_71_65 gnd C_bl
Rb_71_66 bit_71_66 bit_71_67 R_bl
Rbb_71_66 bitb_71_66 bitb_71_67 R_bl
Cb_71_66 bit_71_66 gnd C_bl
Cbb_71_66 bitb_71_66 gnd C_bl
Rb_71_67 bit_71_67 bit_71_68 R_bl
Rbb_71_67 bitb_71_67 bitb_71_68 R_bl
Cb_71_67 bit_71_67 gnd C_bl
Cbb_71_67 bitb_71_67 gnd C_bl
Rb_71_68 bit_71_68 bit_71_69 R_bl
Rbb_71_68 bitb_71_68 bitb_71_69 R_bl
Cb_71_68 bit_71_68 gnd C_bl
Cbb_71_68 bitb_71_68 gnd C_bl
Rb_71_69 bit_71_69 bit_71_70 R_bl
Rbb_71_69 bitb_71_69 bitb_71_70 R_bl
Cb_71_69 bit_71_69 gnd C_bl
Cbb_71_69 bitb_71_69 gnd C_bl
Rb_71_70 bit_71_70 bit_71_71 R_bl
Rbb_71_70 bitb_71_70 bitb_71_71 R_bl
Cb_71_70 bit_71_70 gnd C_bl
Cbb_71_70 bitb_71_70 gnd C_bl
Rb_71_71 bit_71_71 bit_71_72 R_bl
Rbb_71_71 bitb_71_71 bitb_71_72 R_bl
Cb_71_71 bit_71_71 gnd C_bl
Cbb_71_71 bitb_71_71 gnd C_bl
Rb_71_72 bit_71_72 bit_71_73 R_bl
Rbb_71_72 bitb_71_72 bitb_71_73 R_bl
Cb_71_72 bit_71_72 gnd C_bl
Cbb_71_72 bitb_71_72 gnd C_bl
Rb_71_73 bit_71_73 bit_71_74 R_bl
Rbb_71_73 bitb_71_73 bitb_71_74 R_bl
Cb_71_73 bit_71_73 gnd C_bl
Cbb_71_73 bitb_71_73 gnd C_bl
Rb_71_74 bit_71_74 bit_71_75 R_bl
Rbb_71_74 bitb_71_74 bitb_71_75 R_bl
Cb_71_74 bit_71_74 gnd C_bl
Cbb_71_74 bitb_71_74 gnd C_bl
Rb_71_75 bit_71_75 bit_71_76 R_bl
Rbb_71_75 bitb_71_75 bitb_71_76 R_bl
Cb_71_75 bit_71_75 gnd C_bl
Cbb_71_75 bitb_71_75 gnd C_bl
Rb_71_76 bit_71_76 bit_71_77 R_bl
Rbb_71_76 bitb_71_76 bitb_71_77 R_bl
Cb_71_76 bit_71_76 gnd C_bl
Cbb_71_76 bitb_71_76 gnd C_bl
Rb_71_77 bit_71_77 bit_71_78 R_bl
Rbb_71_77 bitb_71_77 bitb_71_78 R_bl
Cb_71_77 bit_71_77 gnd C_bl
Cbb_71_77 bitb_71_77 gnd C_bl
Rb_71_78 bit_71_78 bit_71_79 R_bl
Rbb_71_78 bitb_71_78 bitb_71_79 R_bl
Cb_71_78 bit_71_78 gnd C_bl
Cbb_71_78 bitb_71_78 gnd C_bl
Rb_71_79 bit_71_79 bit_71_80 R_bl
Rbb_71_79 bitb_71_79 bitb_71_80 R_bl
Cb_71_79 bit_71_79 gnd C_bl
Cbb_71_79 bitb_71_79 gnd C_bl
Rb_71_80 bit_71_80 bit_71_81 R_bl
Rbb_71_80 bitb_71_80 bitb_71_81 R_bl
Cb_71_80 bit_71_80 gnd C_bl
Cbb_71_80 bitb_71_80 gnd C_bl
Rb_71_81 bit_71_81 bit_71_82 R_bl
Rbb_71_81 bitb_71_81 bitb_71_82 R_bl
Cb_71_81 bit_71_81 gnd C_bl
Cbb_71_81 bitb_71_81 gnd C_bl
Rb_71_82 bit_71_82 bit_71_83 R_bl
Rbb_71_82 bitb_71_82 bitb_71_83 R_bl
Cb_71_82 bit_71_82 gnd C_bl
Cbb_71_82 bitb_71_82 gnd C_bl
Rb_71_83 bit_71_83 bit_71_84 R_bl
Rbb_71_83 bitb_71_83 bitb_71_84 R_bl
Cb_71_83 bit_71_83 gnd C_bl
Cbb_71_83 bitb_71_83 gnd C_bl
Rb_71_84 bit_71_84 bit_71_85 R_bl
Rbb_71_84 bitb_71_84 bitb_71_85 R_bl
Cb_71_84 bit_71_84 gnd C_bl
Cbb_71_84 bitb_71_84 gnd C_bl
Rb_71_85 bit_71_85 bit_71_86 R_bl
Rbb_71_85 bitb_71_85 bitb_71_86 R_bl
Cb_71_85 bit_71_85 gnd C_bl
Cbb_71_85 bitb_71_85 gnd C_bl
Rb_71_86 bit_71_86 bit_71_87 R_bl
Rbb_71_86 bitb_71_86 bitb_71_87 R_bl
Cb_71_86 bit_71_86 gnd C_bl
Cbb_71_86 bitb_71_86 gnd C_bl
Rb_71_87 bit_71_87 bit_71_88 R_bl
Rbb_71_87 bitb_71_87 bitb_71_88 R_bl
Cb_71_87 bit_71_87 gnd C_bl
Cbb_71_87 bitb_71_87 gnd C_bl
Rb_71_88 bit_71_88 bit_71_89 R_bl
Rbb_71_88 bitb_71_88 bitb_71_89 R_bl
Cb_71_88 bit_71_88 gnd C_bl
Cbb_71_88 bitb_71_88 gnd C_bl
Rb_71_89 bit_71_89 bit_71_90 R_bl
Rbb_71_89 bitb_71_89 bitb_71_90 R_bl
Cb_71_89 bit_71_89 gnd C_bl
Cbb_71_89 bitb_71_89 gnd C_bl
Rb_71_90 bit_71_90 bit_71_91 R_bl
Rbb_71_90 bitb_71_90 bitb_71_91 R_bl
Cb_71_90 bit_71_90 gnd C_bl
Cbb_71_90 bitb_71_90 gnd C_bl
Rb_71_91 bit_71_91 bit_71_92 R_bl
Rbb_71_91 bitb_71_91 bitb_71_92 R_bl
Cb_71_91 bit_71_91 gnd C_bl
Cbb_71_91 bitb_71_91 gnd C_bl
Rb_71_92 bit_71_92 bit_71_93 R_bl
Rbb_71_92 bitb_71_92 bitb_71_93 R_bl
Cb_71_92 bit_71_92 gnd C_bl
Cbb_71_92 bitb_71_92 gnd C_bl
Rb_71_93 bit_71_93 bit_71_94 R_bl
Rbb_71_93 bitb_71_93 bitb_71_94 R_bl
Cb_71_93 bit_71_93 gnd C_bl
Cbb_71_93 bitb_71_93 gnd C_bl
Rb_71_94 bit_71_94 bit_71_95 R_bl
Rbb_71_94 bitb_71_94 bitb_71_95 R_bl
Cb_71_94 bit_71_94 gnd C_bl
Cbb_71_94 bitb_71_94 gnd C_bl
Rb_71_95 bit_71_95 bit_71_96 R_bl
Rbb_71_95 bitb_71_95 bitb_71_96 R_bl
Cb_71_95 bit_71_95 gnd C_bl
Cbb_71_95 bitb_71_95 gnd C_bl
Rb_71_96 bit_71_96 bit_71_97 R_bl
Rbb_71_96 bitb_71_96 bitb_71_97 R_bl
Cb_71_96 bit_71_96 gnd C_bl
Cbb_71_96 bitb_71_96 gnd C_bl
Rb_71_97 bit_71_97 bit_71_98 R_bl
Rbb_71_97 bitb_71_97 bitb_71_98 R_bl
Cb_71_97 bit_71_97 gnd C_bl
Cbb_71_97 bitb_71_97 gnd C_bl
Rb_71_98 bit_71_98 bit_71_99 R_bl
Rbb_71_98 bitb_71_98 bitb_71_99 R_bl
Cb_71_98 bit_71_98 gnd C_bl
Cbb_71_98 bitb_71_98 gnd C_bl
Rb_71_99 bit_71_99 bit_71_100 R_bl
Rbb_71_99 bitb_71_99 bitb_71_100 R_bl
Cb_71_99 bit_71_99 gnd C_bl
Cbb_71_99 bitb_71_99 gnd C_bl
Rb_72_0 bit_72_0 bit_72_1 R_bl
Rbb_72_0 bitb_72_0 bitb_72_1 R_bl
Cb_72_0 bit_72_0 gnd C_bl
Cbb_72_0 bitb_72_0 gnd C_bl
Rb_72_1 bit_72_1 bit_72_2 R_bl
Rbb_72_1 bitb_72_1 bitb_72_2 R_bl
Cb_72_1 bit_72_1 gnd C_bl
Cbb_72_1 bitb_72_1 gnd C_bl
Rb_72_2 bit_72_2 bit_72_3 R_bl
Rbb_72_2 bitb_72_2 bitb_72_3 R_bl
Cb_72_2 bit_72_2 gnd C_bl
Cbb_72_2 bitb_72_2 gnd C_bl
Rb_72_3 bit_72_3 bit_72_4 R_bl
Rbb_72_3 bitb_72_3 bitb_72_4 R_bl
Cb_72_3 bit_72_3 gnd C_bl
Cbb_72_3 bitb_72_3 gnd C_bl
Rb_72_4 bit_72_4 bit_72_5 R_bl
Rbb_72_4 bitb_72_4 bitb_72_5 R_bl
Cb_72_4 bit_72_4 gnd C_bl
Cbb_72_4 bitb_72_4 gnd C_bl
Rb_72_5 bit_72_5 bit_72_6 R_bl
Rbb_72_5 bitb_72_5 bitb_72_6 R_bl
Cb_72_5 bit_72_5 gnd C_bl
Cbb_72_5 bitb_72_5 gnd C_bl
Rb_72_6 bit_72_6 bit_72_7 R_bl
Rbb_72_6 bitb_72_6 bitb_72_7 R_bl
Cb_72_6 bit_72_6 gnd C_bl
Cbb_72_6 bitb_72_6 gnd C_bl
Rb_72_7 bit_72_7 bit_72_8 R_bl
Rbb_72_7 bitb_72_7 bitb_72_8 R_bl
Cb_72_7 bit_72_7 gnd C_bl
Cbb_72_7 bitb_72_7 gnd C_bl
Rb_72_8 bit_72_8 bit_72_9 R_bl
Rbb_72_8 bitb_72_8 bitb_72_9 R_bl
Cb_72_8 bit_72_8 gnd C_bl
Cbb_72_8 bitb_72_8 gnd C_bl
Rb_72_9 bit_72_9 bit_72_10 R_bl
Rbb_72_9 bitb_72_9 bitb_72_10 R_bl
Cb_72_9 bit_72_9 gnd C_bl
Cbb_72_9 bitb_72_9 gnd C_bl
Rb_72_10 bit_72_10 bit_72_11 R_bl
Rbb_72_10 bitb_72_10 bitb_72_11 R_bl
Cb_72_10 bit_72_10 gnd C_bl
Cbb_72_10 bitb_72_10 gnd C_bl
Rb_72_11 bit_72_11 bit_72_12 R_bl
Rbb_72_11 bitb_72_11 bitb_72_12 R_bl
Cb_72_11 bit_72_11 gnd C_bl
Cbb_72_11 bitb_72_11 gnd C_bl
Rb_72_12 bit_72_12 bit_72_13 R_bl
Rbb_72_12 bitb_72_12 bitb_72_13 R_bl
Cb_72_12 bit_72_12 gnd C_bl
Cbb_72_12 bitb_72_12 gnd C_bl
Rb_72_13 bit_72_13 bit_72_14 R_bl
Rbb_72_13 bitb_72_13 bitb_72_14 R_bl
Cb_72_13 bit_72_13 gnd C_bl
Cbb_72_13 bitb_72_13 gnd C_bl
Rb_72_14 bit_72_14 bit_72_15 R_bl
Rbb_72_14 bitb_72_14 bitb_72_15 R_bl
Cb_72_14 bit_72_14 gnd C_bl
Cbb_72_14 bitb_72_14 gnd C_bl
Rb_72_15 bit_72_15 bit_72_16 R_bl
Rbb_72_15 bitb_72_15 bitb_72_16 R_bl
Cb_72_15 bit_72_15 gnd C_bl
Cbb_72_15 bitb_72_15 gnd C_bl
Rb_72_16 bit_72_16 bit_72_17 R_bl
Rbb_72_16 bitb_72_16 bitb_72_17 R_bl
Cb_72_16 bit_72_16 gnd C_bl
Cbb_72_16 bitb_72_16 gnd C_bl
Rb_72_17 bit_72_17 bit_72_18 R_bl
Rbb_72_17 bitb_72_17 bitb_72_18 R_bl
Cb_72_17 bit_72_17 gnd C_bl
Cbb_72_17 bitb_72_17 gnd C_bl
Rb_72_18 bit_72_18 bit_72_19 R_bl
Rbb_72_18 bitb_72_18 bitb_72_19 R_bl
Cb_72_18 bit_72_18 gnd C_bl
Cbb_72_18 bitb_72_18 gnd C_bl
Rb_72_19 bit_72_19 bit_72_20 R_bl
Rbb_72_19 bitb_72_19 bitb_72_20 R_bl
Cb_72_19 bit_72_19 gnd C_bl
Cbb_72_19 bitb_72_19 gnd C_bl
Rb_72_20 bit_72_20 bit_72_21 R_bl
Rbb_72_20 bitb_72_20 bitb_72_21 R_bl
Cb_72_20 bit_72_20 gnd C_bl
Cbb_72_20 bitb_72_20 gnd C_bl
Rb_72_21 bit_72_21 bit_72_22 R_bl
Rbb_72_21 bitb_72_21 bitb_72_22 R_bl
Cb_72_21 bit_72_21 gnd C_bl
Cbb_72_21 bitb_72_21 gnd C_bl
Rb_72_22 bit_72_22 bit_72_23 R_bl
Rbb_72_22 bitb_72_22 bitb_72_23 R_bl
Cb_72_22 bit_72_22 gnd C_bl
Cbb_72_22 bitb_72_22 gnd C_bl
Rb_72_23 bit_72_23 bit_72_24 R_bl
Rbb_72_23 bitb_72_23 bitb_72_24 R_bl
Cb_72_23 bit_72_23 gnd C_bl
Cbb_72_23 bitb_72_23 gnd C_bl
Rb_72_24 bit_72_24 bit_72_25 R_bl
Rbb_72_24 bitb_72_24 bitb_72_25 R_bl
Cb_72_24 bit_72_24 gnd C_bl
Cbb_72_24 bitb_72_24 gnd C_bl
Rb_72_25 bit_72_25 bit_72_26 R_bl
Rbb_72_25 bitb_72_25 bitb_72_26 R_bl
Cb_72_25 bit_72_25 gnd C_bl
Cbb_72_25 bitb_72_25 gnd C_bl
Rb_72_26 bit_72_26 bit_72_27 R_bl
Rbb_72_26 bitb_72_26 bitb_72_27 R_bl
Cb_72_26 bit_72_26 gnd C_bl
Cbb_72_26 bitb_72_26 gnd C_bl
Rb_72_27 bit_72_27 bit_72_28 R_bl
Rbb_72_27 bitb_72_27 bitb_72_28 R_bl
Cb_72_27 bit_72_27 gnd C_bl
Cbb_72_27 bitb_72_27 gnd C_bl
Rb_72_28 bit_72_28 bit_72_29 R_bl
Rbb_72_28 bitb_72_28 bitb_72_29 R_bl
Cb_72_28 bit_72_28 gnd C_bl
Cbb_72_28 bitb_72_28 gnd C_bl
Rb_72_29 bit_72_29 bit_72_30 R_bl
Rbb_72_29 bitb_72_29 bitb_72_30 R_bl
Cb_72_29 bit_72_29 gnd C_bl
Cbb_72_29 bitb_72_29 gnd C_bl
Rb_72_30 bit_72_30 bit_72_31 R_bl
Rbb_72_30 bitb_72_30 bitb_72_31 R_bl
Cb_72_30 bit_72_30 gnd C_bl
Cbb_72_30 bitb_72_30 gnd C_bl
Rb_72_31 bit_72_31 bit_72_32 R_bl
Rbb_72_31 bitb_72_31 bitb_72_32 R_bl
Cb_72_31 bit_72_31 gnd C_bl
Cbb_72_31 bitb_72_31 gnd C_bl
Rb_72_32 bit_72_32 bit_72_33 R_bl
Rbb_72_32 bitb_72_32 bitb_72_33 R_bl
Cb_72_32 bit_72_32 gnd C_bl
Cbb_72_32 bitb_72_32 gnd C_bl
Rb_72_33 bit_72_33 bit_72_34 R_bl
Rbb_72_33 bitb_72_33 bitb_72_34 R_bl
Cb_72_33 bit_72_33 gnd C_bl
Cbb_72_33 bitb_72_33 gnd C_bl
Rb_72_34 bit_72_34 bit_72_35 R_bl
Rbb_72_34 bitb_72_34 bitb_72_35 R_bl
Cb_72_34 bit_72_34 gnd C_bl
Cbb_72_34 bitb_72_34 gnd C_bl
Rb_72_35 bit_72_35 bit_72_36 R_bl
Rbb_72_35 bitb_72_35 bitb_72_36 R_bl
Cb_72_35 bit_72_35 gnd C_bl
Cbb_72_35 bitb_72_35 gnd C_bl
Rb_72_36 bit_72_36 bit_72_37 R_bl
Rbb_72_36 bitb_72_36 bitb_72_37 R_bl
Cb_72_36 bit_72_36 gnd C_bl
Cbb_72_36 bitb_72_36 gnd C_bl
Rb_72_37 bit_72_37 bit_72_38 R_bl
Rbb_72_37 bitb_72_37 bitb_72_38 R_bl
Cb_72_37 bit_72_37 gnd C_bl
Cbb_72_37 bitb_72_37 gnd C_bl
Rb_72_38 bit_72_38 bit_72_39 R_bl
Rbb_72_38 bitb_72_38 bitb_72_39 R_bl
Cb_72_38 bit_72_38 gnd C_bl
Cbb_72_38 bitb_72_38 gnd C_bl
Rb_72_39 bit_72_39 bit_72_40 R_bl
Rbb_72_39 bitb_72_39 bitb_72_40 R_bl
Cb_72_39 bit_72_39 gnd C_bl
Cbb_72_39 bitb_72_39 gnd C_bl
Rb_72_40 bit_72_40 bit_72_41 R_bl
Rbb_72_40 bitb_72_40 bitb_72_41 R_bl
Cb_72_40 bit_72_40 gnd C_bl
Cbb_72_40 bitb_72_40 gnd C_bl
Rb_72_41 bit_72_41 bit_72_42 R_bl
Rbb_72_41 bitb_72_41 bitb_72_42 R_bl
Cb_72_41 bit_72_41 gnd C_bl
Cbb_72_41 bitb_72_41 gnd C_bl
Rb_72_42 bit_72_42 bit_72_43 R_bl
Rbb_72_42 bitb_72_42 bitb_72_43 R_bl
Cb_72_42 bit_72_42 gnd C_bl
Cbb_72_42 bitb_72_42 gnd C_bl
Rb_72_43 bit_72_43 bit_72_44 R_bl
Rbb_72_43 bitb_72_43 bitb_72_44 R_bl
Cb_72_43 bit_72_43 gnd C_bl
Cbb_72_43 bitb_72_43 gnd C_bl
Rb_72_44 bit_72_44 bit_72_45 R_bl
Rbb_72_44 bitb_72_44 bitb_72_45 R_bl
Cb_72_44 bit_72_44 gnd C_bl
Cbb_72_44 bitb_72_44 gnd C_bl
Rb_72_45 bit_72_45 bit_72_46 R_bl
Rbb_72_45 bitb_72_45 bitb_72_46 R_bl
Cb_72_45 bit_72_45 gnd C_bl
Cbb_72_45 bitb_72_45 gnd C_bl
Rb_72_46 bit_72_46 bit_72_47 R_bl
Rbb_72_46 bitb_72_46 bitb_72_47 R_bl
Cb_72_46 bit_72_46 gnd C_bl
Cbb_72_46 bitb_72_46 gnd C_bl
Rb_72_47 bit_72_47 bit_72_48 R_bl
Rbb_72_47 bitb_72_47 bitb_72_48 R_bl
Cb_72_47 bit_72_47 gnd C_bl
Cbb_72_47 bitb_72_47 gnd C_bl
Rb_72_48 bit_72_48 bit_72_49 R_bl
Rbb_72_48 bitb_72_48 bitb_72_49 R_bl
Cb_72_48 bit_72_48 gnd C_bl
Cbb_72_48 bitb_72_48 gnd C_bl
Rb_72_49 bit_72_49 bit_72_50 R_bl
Rbb_72_49 bitb_72_49 bitb_72_50 R_bl
Cb_72_49 bit_72_49 gnd C_bl
Cbb_72_49 bitb_72_49 gnd C_bl
Rb_72_50 bit_72_50 bit_72_51 R_bl
Rbb_72_50 bitb_72_50 bitb_72_51 R_bl
Cb_72_50 bit_72_50 gnd C_bl
Cbb_72_50 bitb_72_50 gnd C_bl
Rb_72_51 bit_72_51 bit_72_52 R_bl
Rbb_72_51 bitb_72_51 bitb_72_52 R_bl
Cb_72_51 bit_72_51 gnd C_bl
Cbb_72_51 bitb_72_51 gnd C_bl
Rb_72_52 bit_72_52 bit_72_53 R_bl
Rbb_72_52 bitb_72_52 bitb_72_53 R_bl
Cb_72_52 bit_72_52 gnd C_bl
Cbb_72_52 bitb_72_52 gnd C_bl
Rb_72_53 bit_72_53 bit_72_54 R_bl
Rbb_72_53 bitb_72_53 bitb_72_54 R_bl
Cb_72_53 bit_72_53 gnd C_bl
Cbb_72_53 bitb_72_53 gnd C_bl
Rb_72_54 bit_72_54 bit_72_55 R_bl
Rbb_72_54 bitb_72_54 bitb_72_55 R_bl
Cb_72_54 bit_72_54 gnd C_bl
Cbb_72_54 bitb_72_54 gnd C_bl
Rb_72_55 bit_72_55 bit_72_56 R_bl
Rbb_72_55 bitb_72_55 bitb_72_56 R_bl
Cb_72_55 bit_72_55 gnd C_bl
Cbb_72_55 bitb_72_55 gnd C_bl
Rb_72_56 bit_72_56 bit_72_57 R_bl
Rbb_72_56 bitb_72_56 bitb_72_57 R_bl
Cb_72_56 bit_72_56 gnd C_bl
Cbb_72_56 bitb_72_56 gnd C_bl
Rb_72_57 bit_72_57 bit_72_58 R_bl
Rbb_72_57 bitb_72_57 bitb_72_58 R_bl
Cb_72_57 bit_72_57 gnd C_bl
Cbb_72_57 bitb_72_57 gnd C_bl
Rb_72_58 bit_72_58 bit_72_59 R_bl
Rbb_72_58 bitb_72_58 bitb_72_59 R_bl
Cb_72_58 bit_72_58 gnd C_bl
Cbb_72_58 bitb_72_58 gnd C_bl
Rb_72_59 bit_72_59 bit_72_60 R_bl
Rbb_72_59 bitb_72_59 bitb_72_60 R_bl
Cb_72_59 bit_72_59 gnd C_bl
Cbb_72_59 bitb_72_59 gnd C_bl
Rb_72_60 bit_72_60 bit_72_61 R_bl
Rbb_72_60 bitb_72_60 bitb_72_61 R_bl
Cb_72_60 bit_72_60 gnd C_bl
Cbb_72_60 bitb_72_60 gnd C_bl
Rb_72_61 bit_72_61 bit_72_62 R_bl
Rbb_72_61 bitb_72_61 bitb_72_62 R_bl
Cb_72_61 bit_72_61 gnd C_bl
Cbb_72_61 bitb_72_61 gnd C_bl
Rb_72_62 bit_72_62 bit_72_63 R_bl
Rbb_72_62 bitb_72_62 bitb_72_63 R_bl
Cb_72_62 bit_72_62 gnd C_bl
Cbb_72_62 bitb_72_62 gnd C_bl
Rb_72_63 bit_72_63 bit_72_64 R_bl
Rbb_72_63 bitb_72_63 bitb_72_64 R_bl
Cb_72_63 bit_72_63 gnd C_bl
Cbb_72_63 bitb_72_63 gnd C_bl
Rb_72_64 bit_72_64 bit_72_65 R_bl
Rbb_72_64 bitb_72_64 bitb_72_65 R_bl
Cb_72_64 bit_72_64 gnd C_bl
Cbb_72_64 bitb_72_64 gnd C_bl
Rb_72_65 bit_72_65 bit_72_66 R_bl
Rbb_72_65 bitb_72_65 bitb_72_66 R_bl
Cb_72_65 bit_72_65 gnd C_bl
Cbb_72_65 bitb_72_65 gnd C_bl
Rb_72_66 bit_72_66 bit_72_67 R_bl
Rbb_72_66 bitb_72_66 bitb_72_67 R_bl
Cb_72_66 bit_72_66 gnd C_bl
Cbb_72_66 bitb_72_66 gnd C_bl
Rb_72_67 bit_72_67 bit_72_68 R_bl
Rbb_72_67 bitb_72_67 bitb_72_68 R_bl
Cb_72_67 bit_72_67 gnd C_bl
Cbb_72_67 bitb_72_67 gnd C_bl
Rb_72_68 bit_72_68 bit_72_69 R_bl
Rbb_72_68 bitb_72_68 bitb_72_69 R_bl
Cb_72_68 bit_72_68 gnd C_bl
Cbb_72_68 bitb_72_68 gnd C_bl
Rb_72_69 bit_72_69 bit_72_70 R_bl
Rbb_72_69 bitb_72_69 bitb_72_70 R_bl
Cb_72_69 bit_72_69 gnd C_bl
Cbb_72_69 bitb_72_69 gnd C_bl
Rb_72_70 bit_72_70 bit_72_71 R_bl
Rbb_72_70 bitb_72_70 bitb_72_71 R_bl
Cb_72_70 bit_72_70 gnd C_bl
Cbb_72_70 bitb_72_70 gnd C_bl
Rb_72_71 bit_72_71 bit_72_72 R_bl
Rbb_72_71 bitb_72_71 bitb_72_72 R_bl
Cb_72_71 bit_72_71 gnd C_bl
Cbb_72_71 bitb_72_71 gnd C_bl
Rb_72_72 bit_72_72 bit_72_73 R_bl
Rbb_72_72 bitb_72_72 bitb_72_73 R_bl
Cb_72_72 bit_72_72 gnd C_bl
Cbb_72_72 bitb_72_72 gnd C_bl
Rb_72_73 bit_72_73 bit_72_74 R_bl
Rbb_72_73 bitb_72_73 bitb_72_74 R_bl
Cb_72_73 bit_72_73 gnd C_bl
Cbb_72_73 bitb_72_73 gnd C_bl
Rb_72_74 bit_72_74 bit_72_75 R_bl
Rbb_72_74 bitb_72_74 bitb_72_75 R_bl
Cb_72_74 bit_72_74 gnd C_bl
Cbb_72_74 bitb_72_74 gnd C_bl
Rb_72_75 bit_72_75 bit_72_76 R_bl
Rbb_72_75 bitb_72_75 bitb_72_76 R_bl
Cb_72_75 bit_72_75 gnd C_bl
Cbb_72_75 bitb_72_75 gnd C_bl
Rb_72_76 bit_72_76 bit_72_77 R_bl
Rbb_72_76 bitb_72_76 bitb_72_77 R_bl
Cb_72_76 bit_72_76 gnd C_bl
Cbb_72_76 bitb_72_76 gnd C_bl
Rb_72_77 bit_72_77 bit_72_78 R_bl
Rbb_72_77 bitb_72_77 bitb_72_78 R_bl
Cb_72_77 bit_72_77 gnd C_bl
Cbb_72_77 bitb_72_77 gnd C_bl
Rb_72_78 bit_72_78 bit_72_79 R_bl
Rbb_72_78 bitb_72_78 bitb_72_79 R_bl
Cb_72_78 bit_72_78 gnd C_bl
Cbb_72_78 bitb_72_78 gnd C_bl
Rb_72_79 bit_72_79 bit_72_80 R_bl
Rbb_72_79 bitb_72_79 bitb_72_80 R_bl
Cb_72_79 bit_72_79 gnd C_bl
Cbb_72_79 bitb_72_79 gnd C_bl
Rb_72_80 bit_72_80 bit_72_81 R_bl
Rbb_72_80 bitb_72_80 bitb_72_81 R_bl
Cb_72_80 bit_72_80 gnd C_bl
Cbb_72_80 bitb_72_80 gnd C_bl
Rb_72_81 bit_72_81 bit_72_82 R_bl
Rbb_72_81 bitb_72_81 bitb_72_82 R_bl
Cb_72_81 bit_72_81 gnd C_bl
Cbb_72_81 bitb_72_81 gnd C_bl
Rb_72_82 bit_72_82 bit_72_83 R_bl
Rbb_72_82 bitb_72_82 bitb_72_83 R_bl
Cb_72_82 bit_72_82 gnd C_bl
Cbb_72_82 bitb_72_82 gnd C_bl
Rb_72_83 bit_72_83 bit_72_84 R_bl
Rbb_72_83 bitb_72_83 bitb_72_84 R_bl
Cb_72_83 bit_72_83 gnd C_bl
Cbb_72_83 bitb_72_83 gnd C_bl
Rb_72_84 bit_72_84 bit_72_85 R_bl
Rbb_72_84 bitb_72_84 bitb_72_85 R_bl
Cb_72_84 bit_72_84 gnd C_bl
Cbb_72_84 bitb_72_84 gnd C_bl
Rb_72_85 bit_72_85 bit_72_86 R_bl
Rbb_72_85 bitb_72_85 bitb_72_86 R_bl
Cb_72_85 bit_72_85 gnd C_bl
Cbb_72_85 bitb_72_85 gnd C_bl
Rb_72_86 bit_72_86 bit_72_87 R_bl
Rbb_72_86 bitb_72_86 bitb_72_87 R_bl
Cb_72_86 bit_72_86 gnd C_bl
Cbb_72_86 bitb_72_86 gnd C_bl
Rb_72_87 bit_72_87 bit_72_88 R_bl
Rbb_72_87 bitb_72_87 bitb_72_88 R_bl
Cb_72_87 bit_72_87 gnd C_bl
Cbb_72_87 bitb_72_87 gnd C_bl
Rb_72_88 bit_72_88 bit_72_89 R_bl
Rbb_72_88 bitb_72_88 bitb_72_89 R_bl
Cb_72_88 bit_72_88 gnd C_bl
Cbb_72_88 bitb_72_88 gnd C_bl
Rb_72_89 bit_72_89 bit_72_90 R_bl
Rbb_72_89 bitb_72_89 bitb_72_90 R_bl
Cb_72_89 bit_72_89 gnd C_bl
Cbb_72_89 bitb_72_89 gnd C_bl
Rb_72_90 bit_72_90 bit_72_91 R_bl
Rbb_72_90 bitb_72_90 bitb_72_91 R_bl
Cb_72_90 bit_72_90 gnd C_bl
Cbb_72_90 bitb_72_90 gnd C_bl
Rb_72_91 bit_72_91 bit_72_92 R_bl
Rbb_72_91 bitb_72_91 bitb_72_92 R_bl
Cb_72_91 bit_72_91 gnd C_bl
Cbb_72_91 bitb_72_91 gnd C_bl
Rb_72_92 bit_72_92 bit_72_93 R_bl
Rbb_72_92 bitb_72_92 bitb_72_93 R_bl
Cb_72_92 bit_72_92 gnd C_bl
Cbb_72_92 bitb_72_92 gnd C_bl
Rb_72_93 bit_72_93 bit_72_94 R_bl
Rbb_72_93 bitb_72_93 bitb_72_94 R_bl
Cb_72_93 bit_72_93 gnd C_bl
Cbb_72_93 bitb_72_93 gnd C_bl
Rb_72_94 bit_72_94 bit_72_95 R_bl
Rbb_72_94 bitb_72_94 bitb_72_95 R_bl
Cb_72_94 bit_72_94 gnd C_bl
Cbb_72_94 bitb_72_94 gnd C_bl
Rb_72_95 bit_72_95 bit_72_96 R_bl
Rbb_72_95 bitb_72_95 bitb_72_96 R_bl
Cb_72_95 bit_72_95 gnd C_bl
Cbb_72_95 bitb_72_95 gnd C_bl
Rb_72_96 bit_72_96 bit_72_97 R_bl
Rbb_72_96 bitb_72_96 bitb_72_97 R_bl
Cb_72_96 bit_72_96 gnd C_bl
Cbb_72_96 bitb_72_96 gnd C_bl
Rb_72_97 bit_72_97 bit_72_98 R_bl
Rbb_72_97 bitb_72_97 bitb_72_98 R_bl
Cb_72_97 bit_72_97 gnd C_bl
Cbb_72_97 bitb_72_97 gnd C_bl
Rb_72_98 bit_72_98 bit_72_99 R_bl
Rbb_72_98 bitb_72_98 bitb_72_99 R_bl
Cb_72_98 bit_72_98 gnd C_bl
Cbb_72_98 bitb_72_98 gnd C_bl
Rb_72_99 bit_72_99 bit_72_100 R_bl
Rbb_72_99 bitb_72_99 bitb_72_100 R_bl
Cb_72_99 bit_72_99 gnd C_bl
Cbb_72_99 bitb_72_99 gnd C_bl
Rb_73_0 bit_73_0 bit_73_1 R_bl
Rbb_73_0 bitb_73_0 bitb_73_1 R_bl
Cb_73_0 bit_73_0 gnd C_bl
Cbb_73_0 bitb_73_0 gnd C_bl
Rb_73_1 bit_73_1 bit_73_2 R_bl
Rbb_73_1 bitb_73_1 bitb_73_2 R_bl
Cb_73_1 bit_73_1 gnd C_bl
Cbb_73_1 bitb_73_1 gnd C_bl
Rb_73_2 bit_73_2 bit_73_3 R_bl
Rbb_73_2 bitb_73_2 bitb_73_3 R_bl
Cb_73_2 bit_73_2 gnd C_bl
Cbb_73_2 bitb_73_2 gnd C_bl
Rb_73_3 bit_73_3 bit_73_4 R_bl
Rbb_73_3 bitb_73_3 bitb_73_4 R_bl
Cb_73_3 bit_73_3 gnd C_bl
Cbb_73_3 bitb_73_3 gnd C_bl
Rb_73_4 bit_73_4 bit_73_5 R_bl
Rbb_73_4 bitb_73_4 bitb_73_5 R_bl
Cb_73_4 bit_73_4 gnd C_bl
Cbb_73_4 bitb_73_4 gnd C_bl
Rb_73_5 bit_73_5 bit_73_6 R_bl
Rbb_73_5 bitb_73_5 bitb_73_6 R_bl
Cb_73_5 bit_73_5 gnd C_bl
Cbb_73_5 bitb_73_5 gnd C_bl
Rb_73_6 bit_73_6 bit_73_7 R_bl
Rbb_73_6 bitb_73_6 bitb_73_7 R_bl
Cb_73_6 bit_73_6 gnd C_bl
Cbb_73_6 bitb_73_6 gnd C_bl
Rb_73_7 bit_73_7 bit_73_8 R_bl
Rbb_73_7 bitb_73_7 bitb_73_8 R_bl
Cb_73_7 bit_73_7 gnd C_bl
Cbb_73_7 bitb_73_7 gnd C_bl
Rb_73_8 bit_73_8 bit_73_9 R_bl
Rbb_73_8 bitb_73_8 bitb_73_9 R_bl
Cb_73_8 bit_73_8 gnd C_bl
Cbb_73_8 bitb_73_8 gnd C_bl
Rb_73_9 bit_73_9 bit_73_10 R_bl
Rbb_73_9 bitb_73_9 bitb_73_10 R_bl
Cb_73_9 bit_73_9 gnd C_bl
Cbb_73_9 bitb_73_9 gnd C_bl
Rb_73_10 bit_73_10 bit_73_11 R_bl
Rbb_73_10 bitb_73_10 bitb_73_11 R_bl
Cb_73_10 bit_73_10 gnd C_bl
Cbb_73_10 bitb_73_10 gnd C_bl
Rb_73_11 bit_73_11 bit_73_12 R_bl
Rbb_73_11 bitb_73_11 bitb_73_12 R_bl
Cb_73_11 bit_73_11 gnd C_bl
Cbb_73_11 bitb_73_11 gnd C_bl
Rb_73_12 bit_73_12 bit_73_13 R_bl
Rbb_73_12 bitb_73_12 bitb_73_13 R_bl
Cb_73_12 bit_73_12 gnd C_bl
Cbb_73_12 bitb_73_12 gnd C_bl
Rb_73_13 bit_73_13 bit_73_14 R_bl
Rbb_73_13 bitb_73_13 bitb_73_14 R_bl
Cb_73_13 bit_73_13 gnd C_bl
Cbb_73_13 bitb_73_13 gnd C_bl
Rb_73_14 bit_73_14 bit_73_15 R_bl
Rbb_73_14 bitb_73_14 bitb_73_15 R_bl
Cb_73_14 bit_73_14 gnd C_bl
Cbb_73_14 bitb_73_14 gnd C_bl
Rb_73_15 bit_73_15 bit_73_16 R_bl
Rbb_73_15 bitb_73_15 bitb_73_16 R_bl
Cb_73_15 bit_73_15 gnd C_bl
Cbb_73_15 bitb_73_15 gnd C_bl
Rb_73_16 bit_73_16 bit_73_17 R_bl
Rbb_73_16 bitb_73_16 bitb_73_17 R_bl
Cb_73_16 bit_73_16 gnd C_bl
Cbb_73_16 bitb_73_16 gnd C_bl
Rb_73_17 bit_73_17 bit_73_18 R_bl
Rbb_73_17 bitb_73_17 bitb_73_18 R_bl
Cb_73_17 bit_73_17 gnd C_bl
Cbb_73_17 bitb_73_17 gnd C_bl
Rb_73_18 bit_73_18 bit_73_19 R_bl
Rbb_73_18 bitb_73_18 bitb_73_19 R_bl
Cb_73_18 bit_73_18 gnd C_bl
Cbb_73_18 bitb_73_18 gnd C_bl
Rb_73_19 bit_73_19 bit_73_20 R_bl
Rbb_73_19 bitb_73_19 bitb_73_20 R_bl
Cb_73_19 bit_73_19 gnd C_bl
Cbb_73_19 bitb_73_19 gnd C_bl
Rb_73_20 bit_73_20 bit_73_21 R_bl
Rbb_73_20 bitb_73_20 bitb_73_21 R_bl
Cb_73_20 bit_73_20 gnd C_bl
Cbb_73_20 bitb_73_20 gnd C_bl
Rb_73_21 bit_73_21 bit_73_22 R_bl
Rbb_73_21 bitb_73_21 bitb_73_22 R_bl
Cb_73_21 bit_73_21 gnd C_bl
Cbb_73_21 bitb_73_21 gnd C_bl
Rb_73_22 bit_73_22 bit_73_23 R_bl
Rbb_73_22 bitb_73_22 bitb_73_23 R_bl
Cb_73_22 bit_73_22 gnd C_bl
Cbb_73_22 bitb_73_22 gnd C_bl
Rb_73_23 bit_73_23 bit_73_24 R_bl
Rbb_73_23 bitb_73_23 bitb_73_24 R_bl
Cb_73_23 bit_73_23 gnd C_bl
Cbb_73_23 bitb_73_23 gnd C_bl
Rb_73_24 bit_73_24 bit_73_25 R_bl
Rbb_73_24 bitb_73_24 bitb_73_25 R_bl
Cb_73_24 bit_73_24 gnd C_bl
Cbb_73_24 bitb_73_24 gnd C_bl
Rb_73_25 bit_73_25 bit_73_26 R_bl
Rbb_73_25 bitb_73_25 bitb_73_26 R_bl
Cb_73_25 bit_73_25 gnd C_bl
Cbb_73_25 bitb_73_25 gnd C_bl
Rb_73_26 bit_73_26 bit_73_27 R_bl
Rbb_73_26 bitb_73_26 bitb_73_27 R_bl
Cb_73_26 bit_73_26 gnd C_bl
Cbb_73_26 bitb_73_26 gnd C_bl
Rb_73_27 bit_73_27 bit_73_28 R_bl
Rbb_73_27 bitb_73_27 bitb_73_28 R_bl
Cb_73_27 bit_73_27 gnd C_bl
Cbb_73_27 bitb_73_27 gnd C_bl
Rb_73_28 bit_73_28 bit_73_29 R_bl
Rbb_73_28 bitb_73_28 bitb_73_29 R_bl
Cb_73_28 bit_73_28 gnd C_bl
Cbb_73_28 bitb_73_28 gnd C_bl
Rb_73_29 bit_73_29 bit_73_30 R_bl
Rbb_73_29 bitb_73_29 bitb_73_30 R_bl
Cb_73_29 bit_73_29 gnd C_bl
Cbb_73_29 bitb_73_29 gnd C_bl
Rb_73_30 bit_73_30 bit_73_31 R_bl
Rbb_73_30 bitb_73_30 bitb_73_31 R_bl
Cb_73_30 bit_73_30 gnd C_bl
Cbb_73_30 bitb_73_30 gnd C_bl
Rb_73_31 bit_73_31 bit_73_32 R_bl
Rbb_73_31 bitb_73_31 bitb_73_32 R_bl
Cb_73_31 bit_73_31 gnd C_bl
Cbb_73_31 bitb_73_31 gnd C_bl
Rb_73_32 bit_73_32 bit_73_33 R_bl
Rbb_73_32 bitb_73_32 bitb_73_33 R_bl
Cb_73_32 bit_73_32 gnd C_bl
Cbb_73_32 bitb_73_32 gnd C_bl
Rb_73_33 bit_73_33 bit_73_34 R_bl
Rbb_73_33 bitb_73_33 bitb_73_34 R_bl
Cb_73_33 bit_73_33 gnd C_bl
Cbb_73_33 bitb_73_33 gnd C_bl
Rb_73_34 bit_73_34 bit_73_35 R_bl
Rbb_73_34 bitb_73_34 bitb_73_35 R_bl
Cb_73_34 bit_73_34 gnd C_bl
Cbb_73_34 bitb_73_34 gnd C_bl
Rb_73_35 bit_73_35 bit_73_36 R_bl
Rbb_73_35 bitb_73_35 bitb_73_36 R_bl
Cb_73_35 bit_73_35 gnd C_bl
Cbb_73_35 bitb_73_35 gnd C_bl
Rb_73_36 bit_73_36 bit_73_37 R_bl
Rbb_73_36 bitb_73_36 bitb_73_37 R_bl
Cb_73_36 bit_73_36 gnd C_bl
Cbb_73_36 bitb_73_36 gnd C_bl
Rb_73_37 bit_73_37 bit_73_38 R_bl
Rbb_73_37 bitb_73_37 bitb_73_38 R_bl
Cb_73_37 bit_73_37 gnd C_bl
Cbb_73_37 bitb_73_37 gnd C_bl
Rb_73_38 bit_73_38 bit_73_39 R_bl
Rbb_73_38 bitb_73_38 bitb_73_39 R_bl
Cb_73_38 bit_73_38 gnd C_bl
Cbb_73_38 bitb_73_38 gnd C_bl
Rb_73_39 bit_73_39 bit_73_40 R_bl
Rbb_73_39 bitb_73_39 bitb_73_40 R_bl
Cb_73_39 bit_73_39 gnd C_bl
Cbb_73_39 bitb_73_39 gnd C_bl
Rb_73_40 bit_73_40 bit_73_41 R_bl
Rbb_73_40 bitb_73_40 bitb_73_41 R_bl
Cb_73_40 bit_73_40 gnd C_bl
Cbb_73_40 bitb_73_40 gnd C_bl
Rb_73_41 bit_73_41 bit_73_42 R_bl
Rbb_73_41 bitb_73_41 bitb_73_42 R_bl
Cb_73_41 bit_73_41 gnd C_bl
Cbb_73_41 bitb_73_41 gnd C_bl
Rb_73_42 bit_73_42 bit_73_43 R_bl
Rbb_73_42 bitb_73_42 bitb_73_43 R_bl
Cb_73_42 bit_73_42 gnd C_bl
Cbb_73_42 bitb_73_42 gnd C_bl
Rb_73_43 bit_73_43 bit_73_44 R_bl
Rbb_73_43 bitb_73_43 bitb_73_44 R_bl
Cb_73_43 bit_73_43 gnd C_bl
Cbb_73_43 bitb_73_43 gnd C_bl
Rb_73_44 bit_73_44 bit_73_45 R_bl
Rbb_73_44 bitb_73_44 bitb_73_45 R_bl
Cb_73_44 bit_73_44 gnd C_bl
Cbb_73_44 bitb_73_44 gnd C_bl
Rb_73_45 bit_73_45 bit_73_46 R_bl
Rbb_73_45 bitb_73_45 bitb_73_46 R_bl
Cb_73_45 bit_73_45 gnd C_bl
Cbb_73_45 bitb_73_45 gnd C_bl
Rb_73_46 bit_73_46 bit_73_47 R_bl
Rbb_73_46 bitb_73_46 bitb_73_47 R_bl
Cb_73_46 bit_73_46 gnd C_bl
Cbb_73_46 bitb_73_46 gnd C_bl
Rb_73_47 bit_73_47 bit_73_48 R_bl
Rbb_73_47 bitb_73_47 bitb_73_48 R_bl
Cb_73_47 bit_73_47 gnd C_bl
Cbb_73_47 bitb_73_47 gnd C_bl
Rb_73_48 bit_73_48 bit_73_49 R_bl
Rbb_73_48 bitb_73_48 bitb_73_49 R_bl
Cb_73_48 bit_73_48 gnd C_bl
Cbb_73_48 bitb_73_48 gnd C_bl
Rb_73_49 bit_73_49 bit_73_50 R_bl
Rbb_73_49 bitb_73_49 bitb_73_50 R_bl
Cb_73_49 bit_73_49 gnd C_bl
Cbb_73_49 bitb_73_49 gnd C_bl
Rb_73_50 bit_73_50 bit_73_51 R_bl
Rbb_73_50 bitb_73_50 bitb_73_51 R_bl
Cb_73_50 bit_73_50 gnd C_bl
Cbb_73_50 bitb_73_50 gnd C_bl
Rb_73_51 bit_73_51 bit_73_52 R_bl
Rbb_73_51 bitb_73_51 bitb_73_52 R_bl
Cb_73_51 bit_73_51 gnd C_bl
Cbb_73_51 bitb_73_51 gnd C_bl
Rb_73_52 bit_73_52 bit_73_53 R_bl
Rbb_73_52 bitb_73_52 bitb_73_53 R_bl
Cb_73_52 bit_73_52 gnd C_bl
Cbb_73_52 bitb_73_52 gnd C_bl
Rb_73_53 bit_73_53 bit_73_54 R_bl
Rbb_73_53 bitb_73_53 bitb_73_54 R_bl
Cb_73_53 bit_73_53 gnd C_bl
Cbb_73_53 bitb_73_53 gnd C_bl
Rb_73_54 bit_73_54 bit_73_55 R_bl
Rbb_73_54 bitb_73_54 bitb_73_55 R_bl
Cb_73_54 bit_73_54 gnd C_bl
Cbb_73_54 bitb_73_54 gnd C_bl
Rb_73_55 bit_73_55 bit_73_56 R_bl
Rbb_73_55 bitb_73_55 bitb_73_56 R_bl
Cb_73_55 bit_73_55 gnd C_bl
Cbb_73_55 bitb_73_55 gnd C_bl
Rb_73_56 bit_73_56 bit_73_57 R_bl
Rbb_73_56 bitb_73_56 bitb_73_57 R_bl
Cb_73_56 bit_73_56 gnd C_bl
Cbb_73_56 bitb_73_56 gnd C_bl
Rb_73_57 bit_73_57 bit_73_58 R_bl
Rbb_73_57 bitb_73_57 bitb_73_58 R_bl
Cb_73_57 bit_73_57 gnd C_bl
Cbb_73_57 bitb_73_57 gnd C_bl
Rb_73_58 bit_73_58 bit_73_59 R_bl
Rbb_73_58 bitb_73_58 bitb_73_59 R_bl
Cb_73_58 bit_73_58 gnd C_bl
Cbb_73_58 bitb_73_58 gnd C_bl
Rb_73_59 bit_73_59 bit_73_60 R_bl
Rbb_73_59 bitb_73_59 bitb_73_60 R_bl
Cb_73_59 bit_73_59 gnd C_bl
Cbb_73_59 bitb_73_59 gnd C_bl
Rb_73_60 bit_73_60 bit_73_61 R_bl
Rbb_73_60 bitb_73_60 bitb_73_61 R_bl
Cb_73_60 bit_73_60 gnd C_bl
Cbb_73_60 bitb_73_60 gnd C_bl
Rb_73_61 bit_73_61 bit_73_62 R_bl
Rbb_73_61 bitb_73_61 bitb_73_62 R_bl
Cb_73_61 bit_73_61 gnd C_bl
Cbb_73_61 bitb_73_61 gnd C_bl
Rb_73_62 bit_73_62 bit_73_63 R_bl
Rbb_73_62 bitb_73_62 bitb_73_63 R_bl
Cb_73_62 bit_73_62 gnd C_bl
Cbb_73_62 bitb_73_62 gnd C_bl
Rb_73_63 bit_73_63 bit_73_64 R_bl
Rbb_73_63 bitb_73_63 bitb_73_64 R_bl
Cb_73_63 bit_73_63 gnd C_bl
Cbb_73_63 bitb_73_63 gnd C_bl
Rb_73_64 bit_73_64 bit_73_65 R_bl
Rbb_73_64 bitb_73_64 bitb_73_65 R_bl
Cb_73_64 bit_73_64 gnd C_bl
Cbb_73_64 bitb_73_64 gnd C_bl
Rb_73_65 bit_73_65 bit_73_66 R_bl
Rbb_73_65 bitb_73_65 bitb_73_66 R_bl
Cb_73_65 bit_73_65 gnd C_bl
Cbb_73_65 bitb_73_65 gnd C_bl
Rb_73_66 bit_73_66 bit_73_67 R_bl
Rbb_73_66 bitb_73_66 bitb_73_67 R_bl
Cb_73_66 bit_73_66 gnd C_bl
Cbb_73_66 bitb_73_66 gnd C_bl
Rb_73_67 bit_73_67 bit_73_68 R_bl
Rbb_73_67 bitb_73_67 bitb_73_68 R_bl
Cb_73_67 bit_73_67 gnd C_bl
Cbb_73_67 bitb_73_67 gnd C_bl
Rb_73_68 bit_73_68 bit_73_69 R_bl
Rbb_73_68 bitb_73_68 bitb_73_69 R_bl
Cb_73_68 bit_73_68 gnd C_bl
Cbb_73_68 bitb_73_68 gnd C_bl
Rb_73_69 bit_73_69 bit_73_70 R_bl
Rbb_73_69 bitb_73_69 bitb_73_70 R_bl
Cb_73_69 bit_73_69 gnd C_bl
Cbb_73_69 bitb_73_69 gnd C_bl
Rb_73_70 bit_73_70 bit_73_71 R_bl
Rbb_73_70 bitb_73_70 bitb_73_71 R_bl
Cb_73_70 bit_73_70 gnd C_bl
Cbb_73_70 bitb_73_70 gnd C_bl
Rb_73_71 bit_73_71 bit_73_72 R_bl
Rbb_73_71 bitb_73_71 bitb_73_72 R_bl
Cb_73_71 bit_73_71 gnd C_bl
Cbb_73_71 bitb_73_71 gnd C_bl
Rb_73_72 bit_73_72 bit_73_73 R_bl
Rbb_73_72 bitb_73_72 bitb_73_73 R_bl
Cb_73_72 bit_73_72 gnd C_bl
Cbb_73_72 bitb_73_72 gnd C_bl
Rb_73_73 bit_73_73 bit_73_74 R_bl
Rbb_73_73 bitb_73_73 bitb_73_74 R_bl
Cb_73_73 bit_73_73 gnd C_bl
Cbb_73_73 bitb_73_73 gnd C_bl
Rb_73_74 bit_73_74 bit_73_75 R_bl
Rbb_73_74 bitb_73_74 bitb_73_75 R_bl
Cb_73_74 bit_73_74 gnd C_bl
Cbb_73_74 bitb_73_74 gnd C_bl
Rb_73_75 bit_73_75 bit_73_76 R_bl
Rbb_73_75 bitb_73_75 bitb_73_76 R_bl
Cb_73_75 bit_73_75 gnd C_bl
Cbb_73_75 bitb_73_75 gnd C_bl
Rb_73_76 bit_73_76 bit_73_77 R_bl
Rbb_73_76 bitb_73_76 bitb_73_77 R_bl
Cb_73_76 bit_73_76 gnd C_bl
Cbb_73_76 bitb_73_76 gnd C_bl
Rb_73_77 bit_73_77 bit_73_78 R_bl
Rbb_73_77 bitb_73_77 bitb_73_78 R_bl
Cb_73_77 bit_73_77 gnd C_bl
Cbb_73_77 bitb_73_77 gnd C_bl
Rb_73_78 bit_73_78 bit_73_79 R_bl
Rbb_73_78 bitb_73_78 bitb_73_79 R_bl
Cb_73_78 bit_73_78 gnd C_bl
Cbb_73_78 bitb_73_78 gnd C_bl
Rb_73_79 bit_73_79 bit_73_80 R_bl
Rbb_73_79 bitb_73_79 bitb_73_80 R_bl
Cb_73_79 bit_73_79 gnd C_bl
Cbb_73_79 bitb_73_79 gnd C_bl
Rb_73_80 bit_73_80 bit_73_81 R_bl
Rbb_73_80 bitb_73_80 bitb_73_81 R_bl
Cb_73_80 bit_73_80 gnd C_bl
Cbb_73_80 bitb_73_80 gnd C_bl
Rb_73_81 bit_73_81 bit_73_82 R_bl
Rbb_73_81 bitb_73_81 bitb_73_82 R_bl
Cb_73_81 bit_73_81 gnd C_bl
Cbb_73_81 bitb_73_81 gnd C_bl
Rb_73_82 bit_73_82 bit_73_83 R_bl
Rbb_73_82 bitb_73_82 bitb_73_83 R_bl
Cb_73_82 bit_73_82 gnd C_bl
Cbb_73_82 bitb_73_82 gnd C_bl
Rb_73_83 bit_73_83 bit_73_84 R_bl
Rbb_73_83 bitb_73_83 bitb_73_84 R_bl
Cb_73_83 bit_73_83 gnd C_bl
Cbb_73_83 bitb_73_83 gnd C_bl
Rb_73_84 bit_73_84 bit_73_85 R_bl
Rbb_73_84 bitb_73_84 bitb_73_85 R_bl
Cb_73_84 bit_73_84 gnd C_bl
Cbb_73_84 bitb_73_84 gnd C_bl
Rb_73_85 bit_73_85 bit_73_86 R_bl
Rbb_73_85 bitb_73_85 bitb_73_86 R_bl
Cb_73_85 bit_73_85 gnd C_bl
Cbb_73_85 bitb_73_85 gnd C_bl
Rb_73_86 bit_73_86 bit_73_87 R_bl
Rbb_73_86 bitb_73_86 bitb_73_87 R_bl
Cb_73_86 bit_73_86 gnd C_bl
Cbb_73_86 bitb_73_86 gnd C_bl
Rb_73_87 bit_73_87 bit_73_88 R_bl
Rbb_73_87 bitb_73_87 bitb_73_88 R_bl
Cb_73_87 bit_73_87 gnd C_bl
Cbb_73_87 bitb_73_87 gnd C_bl
Rb_73_88 bit_73_88 bit_73_89 R_bl
Rbb_73_88 bitb_73_88 bitb_73_89 R_bl
Cb_73_88 bit_73_88 gnd C_bl
Cbb_73_88 bitb_73_88 gnd C_bl
Rb_73_89 bit_73_89 bit_73_90 R_bl
Rbb_73_89 bitb_73_89 bitb_73_90 R_bl
Cb_73_89 bit_73_89 gnd C_bl
Cbb_73_89 bitb_73_89 gnd C_bl
Rb_73_90 bit_73_90 bit_73_91 R_bl
Rbb_73_90 bitb_73_90 bitb_73_91 R_bl
Cb_73_90 bit_73_90 gnd C_bl
Cbb_73_90 bitb_73_90 gnd C_bl
Rb_73_91 bit_73_91 bit_73_92 R_bl
Rbb_73_91 bitb_73_91 bitb_73_92 R_bl
Cb_73_91 bit_73_91 gnd C_bl
Cbb_73_91 bitb_73_91 gnd C_bl
Rb_73_92 bit_73_92 bit_73_93 R_bl
Rbb_73_92 bitb_73_92 bitb_73_93 R_bl
Cb_73_92 bit_73_92 gnd C_bl
Cbb_73_92 bitb_73_92 gnd C_bl
Rb_73_93 bit_73_93 bit_73_94 R_bl
Rbb_73_93 bitb_73_93 bitb_73_94 R_bl
Cb_73_93 bit_73_93 gnd C_bl
Cbb_73_93 bitb_73_93 gnd C_bl
Rb_73_94 bit_73_94 bit_73_95 R_bl
Rbb_73_94 bitb_73_94 bitb_73_95 R_bl
Cb_73_94 bit_73_94 gnd C_bl
Cbb_73_94 bitb_73_94 gnd C_bl
Rb_73_95 bit_73_95 bit_73_96 R_bl
Rbb_73_95 bitb_73_95 bitb_73_96 R_bl
Cb_73_95 bit_73_95 gnd C_bl
Cbb_73_95 bitb_73_95 gnd C_bl
Rb_73_96 bit_73_96 bit_73_97 R_bl
Rbb_73_96 bitb_73_96 bitb_73_97 R_bl
Cb_73_96 bit_73_96 gnd C_bl
Cbb_73_96 bitb_73_96 gnd C_bl
Rb_73_97 bit_73_97 bit_73_98 R_bl
Rbb_73_97 bitb_73_97 bitb_73_98 R_bl
Cb_73_97 bit_73_97 gnd C_bl
Cbb_73_97 bitb_73_97 gnd C_bl
Rb_73_98 bit_73_98 bit_73_99 R_bl
Rbb_73_98 bitb_73_98 bitb_73_99 R_bl
Cb_73_98 bit_73_98 gnd C_bl
Cbb_73_98 bitb_73_98 gnd C_bl
Rb_73_99 bit_73_99 bit_73_100 R_bl
Rbb_73_99 bitb_73_99 bitb_73_100 R_bl
Cb_73_99 bit_73_99 gnd C_bl
Cbb_73_99 bitb_73_99 gnd C_bl
Rb_74_0 bit_74_0 bit_74_1 R_bl
Rbb_74_0 bitb_74_0 bitb_74_1 R_bl
Cb_74_0 bit_74_0 gnd C_bl
Cbb_74_0 bitb_74_0 gnd C_bl
Rb_74_1 bit_74_1 bit_74_2 R_bl
Rbb_74_1 bitb_74_1 bitb_74_2 R_bl
Cb_74_1 bit_74_1 gnd C_bl
Cbb_74_1 bitb_74_1 gnd C_bl
Rb_74_2 bit_74_2 bit_74_3 R_bl
Rbb_74_2 bitb_74_2 bitb_74_3 R_bl
Cb_74_2 bit_74_2 gnd C_bl
Cbb_74_2 bitb_74_2 gnd C_bl
Rb_74_3 bit_74_3 bit_74_4 R_bl
Rbb_74_3 bitb_74_3 bitb_74_4 R_bl
Cb_74_3 bit_74_3 gnd C_bl
Cbb_74_3 bitb_74_3 gnd C_bl
Rb_74_4 bit_74_4 bit_74_5 R_bl
Rbb_74_4 bitb_74_4 bitb_74_5 R_bl
Cb_74_4 bit_74_4 gnd C_bl
Cbb_74_4 bitb_74_4 gnd C_bl
Rb_74_5 bit_74_5 bit_74_6 R_bl
Rbb_74_5 bitb_74_5 bitb_74_6 R_bl
Cb_74_5 bit_74_5 gnd C_bl
Cbb_74_5 bitb_74_5 gnd C_bl
Rb_74_6 bit_74_6 bit_74_7 R_bl
Rbb_74_6 bitb_74_6 bitb_74_7 R_bl
Cb_74_6 bit_74_6 gnd C_bl
Cbb_74_6 bitb_74_6 gnd C_bl
Rb_74_7 bit_74_7 bit_74_8 R_bl
Rbb_74_7 bitb_74_7 bitb_74_8 R_bl
Cb_74_7 bit_74_7 gnd C_bl
Cbb_74_7 bitb_74_7 gnd C_bl
Rb_74_8 bit_74_8 bit_74_9 R_bl
Rbb_74_8 bitb_74_8 bitb_74_9 R_bl
Cb_74_8 bit_74_8 gnd C_bl
Cbb_74_8 bitb_74_8 gnd C_bl
Rb_74_9 bit_74_9 bit_74_10 R_bl
Rbb_74_9 bitb_74_9 bitb_74_10 R_bl
Cb_74_9 bit_74_9 gnd C_bl
Cbb_74_9 bitb_74_9 gnd C_bl
Rb_74_10 bit_74_10 bit_74_11 R_bl
Rbb_74_10 bitb_74_10 bitb_74_11 R_bl
Cb_74_10 bit_74_10 gnd C_bl
Cbb_74_10 bitb_74_10 gnd C_bl
Rb_74_11 bit_74_11 bit_74_12 R_bl
Rbb_74_11 bitb_74_11 bitb_74_12 R_bl
Cb_74_11 bit_74_11 gnd C_bl
Cbb_74_11 bitb_74_11 gnd C_bl
Rb_74_12 bit_74_12 bit_74_13 R_bl
Rbb_74_12 bitb_74_12 bitb_74_13 R_bl
Cb_74_12 bit_74_12 gnd C_bl
Cbb_74_12 bitb_74_12 gnd C_bl
Rb_74_13 bit_74_13 bit_74_14 R_bl
Rbb_74_13 bitb_74_13 bitb_74_14 R_bl
Cb_74_13 bit_74_13 gnd C_bl
Cbb_74_13 bitb_74_13 gnd C_bl
Rb_74_14 bit_74_14 bit_74_15 R_bl
Rbb_74_14 bitb_74_14 bitb_74_15 R_bl
Cb_74_14 bit_74_14 gnd C_bl
Cbb_74_14 bitb_74_14 gnd C_bl
Rb_74_15 bit_74_15 bit_74_16 R_bl
Rbb_74_15 bitb_74_15 bitb_74_16 R_bl
Cb_74_15 bit_74_15 gnd C_bl
Cbb_74_15 bitb_74_15 gnd C_bl
Rb_74_16 bit_74_16 bit_74_17 R_bl
Rbb_74_16 bitb_74_16 bitb_74_17 R_bl
Cb_74_16 bit_74_16 gnd C_bl
Cbb_74_16 bitb_74_16 gnd C_bl
Rb_74_17 bit_74_17 bit_74_18 R_bl
Rbb_74_17 bitb_74_17 bitb_74_18 R_bl
Cb_74_17 bit_74_17 gnd C_bl
Cbb_74_17 bitb_74_17 gnd C_bl
Rb_74_18 bit_74_18 bit_74_19 R_bl
Rbb_74_18 bitb_74_18 bitb_74_19 R_bl
Cb_74_18 bit_74_18 gnd C_bl
Cbb_74_18 bitb_74_18 gnd C_bl
Rb_74_19 bit_74_19 bit_74_20 R_bl
Rbb_74_19 bitb_74_19 bitb_74_20 R_bl
Cb_74_19 bit_74_19 gnd C_bl
Cbb_74_19 bitb_74_19 gnd C_bl
Rb_74_20 bit_74_20 bit_74_21 R_bl
Rbb_74_20 bitb_74_20 bitb_74_21 R_bl
Cb_74_20 bit_74_20 gnd C_bl
Cbb_74_20 bitb_74_20 gnd C_bl
Rb_74_21 bit_74_21 bit_74_22 R_bl
Rbb_74_21 bitb_74_21 bitb_74_22 R_bl
Cb_74_21 bit_74_21 gnd C_bl
Cbb_74_21 bitb_74_21 gnd C_bl
Rb_74_22 bit_74_22 bit_74_23 R_bl
Rbb_74_22 bitb_74_22 bitb_74_23 R_bl
Cb_74_22 bit_74_22 gnd C_bl
Cbb_74_22 bitb_74_22 gnd C_bl
Rb_74_23 bit_74_23 bit_74_24 R_bl
Rbb_74_23 bitb_74_23 bitb_74_24 R_bl
Cb_74_23 bit_74_23 gnd C_bl
Cbb_74_23 bitb_74_23 gnd C_bl
Rb_74_24 bit_74_24 bit_74_25 R_bl
Rbb_74_24 bitb_74_24 bitb_74_25 R_bl
Cb_74_24 bit_74_24 gnd C_bl
Cbb_74_24 bitb_74_24 gnd C_bl
Rb_74_25 bit_74_25 bit_74_26 R_bl
Rbb_74_25 bitb_74_25 bitb_74_26 R_bl
Cb_74_25 bit_74_25 gnd C_bl
Cbb_74_25 bitb_74_25 gnd C_bl
Rb_74_26 bit_74_26 bit_74_27 R_bl
Rbb_74_26 bitb_74_26 bitb_74_27 R_bl
Cb_74_26 bit_74_26 gnd C_bl
Cbb_74_26 bitb_74_26 gnd C_bl
Rb_74_27 bit_74_27 bit_74_28 R_bl
Rbb_74_27 bitb_74_27 bitb_74_28 R_bl
Cb_74_27 bit_74_27 gnd C_bl
Cbb_74_27 bitb_74_27 gnd C_bl
Rb_74_28 bit_74_28 bit_74_29 R_bl
Rbb_74_28 bitb_74_28 bitb_74_29 R_bl
Cb_74_28 bit_74_28 gnd C_bl
Cbb_74_28 bitb_74_28 gnd C_bl
Rb_74_29 bit_74_29 bit_74_30 R_bl
Rbb_74_29 bitb_74_29 bitb_74_30 R_bl
Cb_74_29 bit_74_29 gnd C_bl
Cbb_74_29 bitb_74_29 gnd C_bl
Rb_74_30 bit_74_30 bit_74_31 R_bl
Rbb_74_30 bitb_74_30 bitb_74_31 R_bl
Cb_74_30 bit_74_30 gnd C_bl
Cbb_74_30 bitb_74_30 gnd C_bl
Rb_74_31 bit_74_31 bit_74_32 R_bl
Rbb_74_31 bitb_74_31 bitb_74_32 R_bl
Cb_74_31 bit_74_31 gnd C_bl
Cbb_74_31 bitb_74_31 gnd C_bl
Rb_74_32 bit_74_32 bit_74_33 R_bl
Rbb_74_32 bitb_74_32 bitb_74_33 R_bl
Cb_74_32 bit_74_32 gnd C_bl
Cbb_74_32 bitb_74_32 gnd C_bl
Rb_74_33 bit_74_33 bit_74_34 R_bl
Rbb_74_33 bitb_74_33 bitb_74_34 R_bl
Cb_74_33 bit_74_33 gnd C_bl
Cbb_74_33 bitb_74_33 gnd C_bl
Rb_74_34 bit_74_34 bit_74_35 R_bl
Rbb_74_34 bitb_74_34 bitb_74_35 R_bl
Cb_74_34 bit_74_34 gnd C_bl
Cbb_74_34 bitb_74_34 gnd C_bl
Rb_74_35 bit_74_35 bit_74_36 R_bl
Rbb_74_35 bitb_74_35 bitb_74_36 R_bl
Cb_74_35 bit_74_35 gnd C_bl
Cbb_74_35 bitb_74_35 gnd C_bl
Rb_74_36 bit_74_36 bit_74_37 R_bl
Rbb_74_36 bitb_74_36 bitb_74_37 R_bl
Cb_74_36 bit_74_36 gnd C_bl
Cbb_74_36 bitb_74_36 gnd C_bl
Rb_74_37 bit_74_37 bit_74_38 R_bl
Rbb_74_37 bitb_74_37 bitb_74_38 R_bl
Cb_74_37 bit_74_37 gnd C_bl
Cbb_74_37 bitb_74_37 gnd C_bl
Rb_74_38 bit_74_38 bit_74_39 R_bl
Rbb_74_38 bitb_74_38 bitb_74_39 R_bl
Cb_74_38 bit_74_38 gnd C_bl
Cbb_74_38 bitb_74_38 gnd C_bl
Rb_74_39 bit_74_39 bit_74_40 R_bl
Rbb_74_39 bitb_74_39 bitb_74_40 R_bl
Cb_74_39 bit_74_39 gnd C_bl
Cbb_74_39 bitb_74_39 gnd C_bl
Rb_74_40 bit_74_40 bit_74_41 R_bl
Rbb_74_40 bitb_74_40 bitb_74_41 R_bl
Cb_74_40 bit_74_40 gnd C_bl
Cbb_74_40 bitb_74_40 gnd C_bl
Rb_74_41 bit_74_41 bit_74_42 R_bl
Rbb_74_41 bitb_74_41 bitb_74_42 R_bl
Cb_74_41 bit_74_41 gnd C_bl
Cbb_74_41 bitb_74_41 gnd C_bl
Rb_74_42 bit_74_42 bit_74_43 R_bl
Rbb_74_42 bitb_74_42 bitb_74_43 R_bl
Cb_74_42 bit_74_42 gnd C_bl
Cbb_74_42 bitb_74_42 gnd C_bl
Rb_74_43 bit_74_43 bit_74_44 R_bl
Rbb_74_43 bitb_74_43 bitb_74_44 R_bl
Cb_74_43 bit_74_43 gnd C_bl
Cbb_74_43 bitb_74_43 gnd C_bl
Rb_74_44 bit_74_44 bit_74_45 R_bl
Rbb_74_44 bitb_74_44 bitb_74_45 R_bl
Cb_74_44 bit_74_44 gnd C_bl
Cbb_74_44 bitb_74_44 gnd C_bl
Rb_74_45 bit_74_45 bit_74_46 R_bl
Rbb_74_45 bitb_74_45 bitb_74_46 R_bl
Cb_74_45 bit_74_45 gnd C_bl
Cbb_74_45 bitb_74_45 gnd C_bl
Rb_74_46 bit_74_46 bit_74_47 R_bl
Rbb_74_46 bitb_74_46 bitb_74_47 R_bl
Cb_74_46 bit_74_46 gnd C_bl
Cbb_74_46 bitb_74_46 gnd C_bl
Rb_74_47 bit_74_47 bit_74_48 R_bl
Rbb_74_47 bitb_74_47 bitb_74_48 R_bl
Cb_74_47 bit_74_47 gnd C_bl
Cbb_74_47 bitb_74_47 gnd C_bl
Rb_74_48 bit_74_48 bit_74_49 R_bl
Rbb_74_48 bitb_74_48 bitb_74_49 R_bl
Cb_74_48 bit_74_48 gnd C_bl
Cbb_74_48 bitb_74_48 gnd C_bl
Rb_74_49 bit_74_49 bit_74_50 R_bl
Rbb_74_49 bitb_74_49 bitb_74_50 R_bl
Cb_74_49 bit_74_49 gnd C_bl
Cbb_74_49 bitb_74_49 gnd C_bl
Rb_74_50 bit_74_50 bit_74_51 R_bl
Rbb_74_50 bitb_74_50 bitb_74_51 R_bl
Cb_74_50 bit_74_50 gnd C_bl
Cbb_74_50 bitb_74_50 gnd C_bl
Rb_74_51 bit_74_51 bit_74_52 R_bl
Rbb_74_51 bitb_74_51 bitb_74_52 R_bl
Cb_74_51 bit_74_51 gnd C_bl
Cbb_74_51 bitb_74_51 gnd C_bl
Rb_74_52 bit_74_52 bit_74_53 R_bl
Rbb_74_52 bitb_74_52 bitb_74_53 R_bl
Cb_74_52 bit_74_52 gnd C_bl
Cbb_74_52 bitb_74_52 gnd C_bl
Rb_74_53 bit_74_53 bit_74_54 R_bl
Rbb_74_53 bitb_74_53 bitb_74_54 R_bl
Cb_74_53 bit_74_53 gnd C_bl
Cbb_74_53 bitb_74_53 gnd C_bl
Rb_74_54 bit_74_54 bit_74_55 R_bl
Rbb_74_54 bitb_74_54 bitb_74_55 R_bl
Cb_74_54 bit_74_54 gnd C_bl
Cbb_74_54 bitb_74_54 gnd C_bl
Rb_74_55 bit_74_55 bit_74_56 R_bl
Rbb_74_55 bitb_74_55 bitb_74_56 R_bl
Cb_74_55 bit_74_55 gnd C_bl
Cbb_74_55 bitb_74_55 gnd C_bl
Rb_74_56 bit_74_56 bit_74_57 R_bl
Rbb_74_56 bitb_74_56 bitb_74_57 R_bl
Cb_74_56 bit_74_56 gnd C_bl
Cbb_74_56 bitb_74_56 gnd C_bl
Rb_74_57 bit_74_57 bit_74_58 R_bl
Rbb_74_57 bitb_74_57 bitb_74_58 R_bl
Cb_74_57 bit_74_57 gnd C_bl
Cbb_74_57 bitb_74_57 gnd C_bl
Rb_74_58 bit_74_58 bit_74_59 R_bl
Rbb_74_58 bitb_74_58 bitb_74_59 R_bl
Cb_74_58 bit_74_58 gnd C_bl
Cbb_74_58 bitb_74_58 gnd C_bl
Rb_74_59 bit_74_59 bit_74_60 R_bl
Rbb_74_59 bitb_74_59 bitb_74_60 R_bl
Cb_74_59 bit_74_59 gnd C_bl
Cbb_74_59 bitb_74_59 gnd C_bl
Rb_74_60 bit_74_60 bit_74_61 R_bl
Rbb_74_60 bitb_74_60 bitb_74_61 R_bl
Cb_74_60 bit_74_60 gnd C_bl
Cbb_74_60 bitb_74_60 gnd C_bl
Rb_74_61 bit_74_61 bit_74_62 R_bl
Rbb_74_61 bitb_74_61 bitb_74_62 R_bl
Cb_74_61 bit_74_61 gnd C_bl
Cbb_74_61 bitb_74_61 gnd C_bl
Rb_74_62 bit_74_62 bit_74_63 R_bl
Rbb_74_62 bitb_74_62 bitb_74_63 R_bl
Cb_74_62 bit_74_62 gnd C_bl
Cbb_74_62 bitb_74_62 gnd C_bl
Rb_74_63 bit_74_63 bit_74_64 R_bl
Rbb_74_63 bitb_74_63 bitb_74_64 R_bl
Cb_74_63 bit_74_63 gnd C_bl
Cbb_74_63 bitb_74_63 gnd C_bl
Rb_74_64 bit_74_64 bit_74_65 R_bl
Rbb_74_64 bitb_74_64 bitb_74_65 R_bl
Cb_74_64 bit_74_64 gnd C_bl
Cbb_74_64 bitb_74_64 gnd C_bl
Rb_74_65 bit_74_65 bit_74_66 R_bl
Rbb_74_65 bitb_74_65 bitb_74_66 R_bl
Cb_74_65 bit_74_65 gnd C_bl
Cbb_74_65 bitb_74_65 gnd C_bl
Rb_74_66 bit_74_66 bit_74_67 R_bl
Rbb_74_66 bitb_74_66 bitb_74_67 R_bl
Cb_74_66 bit_74_66 gnd C_bl
Cbb_74_66 bitb_74_66 gnd C_bl
Rb_74_67 bit_74_67 bit_74_68 R_bl
Rbb_74_67 bitb_74_67 bitb_74_68 R_bl
Cb_74_67 bit_74_67 gnd C_bl
Cbb_74_67 bitb_74_67 gnd C_bl
Rb_74_68 bit_74_68 bit_74_69 R_bl
Rbb_74_68 bitb_74_68 bitb_74_69 R_bl
Cb_74_68 bit_74_68 gnd C_bl
Cbb_74_68 bitb_74_68 gnd C_bl
Rb_74_69 bit_74_69 bit_74_70 R_bl
Rbb_74_69 bitb_74_69 bitb_74_70 R_bl
Cb_74_69 bit_74_69 gnd C_bl
Cbb_74_69 bitb_74_69 gnd C_bl
Rb_74_70 bit_74_70 bit_74_71 R_bl
Rbb_74_70 bitb_74_70 bitb_74_71 R_bl
Cb_74_70 bit_74_70 gnd C_bl
Cbb_74_70 bitb_74_70 gnd C_bl
Rb_74_71 bit_74_71 bit_74_72 R_bl
Rbb_74_71 bitb_74_71 bitb_74_72 R_bl
Cb_74_71 bit_74_71 gnd C_bl
Cbb_74_71 bitb_74_71 gnd C_bl
Rb_74_72 bit_74_72 bit_74_73 R_bl
Rbb_74_72 bitb_74_72 bitb_74_73 R_bl
Cb_74_72 bit_74_72 gnd C_bl
Cbb_74_72 bitb_74_72 gnd C_bl
Rb_74_73 bit_74_73 bit_74_74 R_bl
Rbb_74_73 bitb_74_73 bitb_74_74 R_bl
Cb_74_73 bit_74_73 gnd C_bl
Cbb_74_73 bitb_74_73 gnd C_bl
Rb_74_74 bit_74_74 bit_74_75 R_bl
Rbb_74_74 bitb_74_74 bitb_74_75 R_bl
Cb_74_74 bit_74_74 gnd C_bl
Cbb_74_74 bitb_74_74 gnd C_bl
Rb_74_75 bit_74_75 bit_74_76 R_bl
Rbb_74_75 bitb_74_75 bitb_74_76 R_bl
Cb_74_75 bit_74_75 gnd C_bl
Cbb_74_75 bitb_74_75 gnd C_bl
Rb_74_76 bit_74_76 bit_74_77 R_bl
Rbb_74_76 bitb_74_76 bitb_74_77 R_bl
Cb_74_76 bit_74_76 gnd C_bl
Cbb_74_76 bitb_74_76 gnd C_bl
Rb_74_77 bit_74_77 bit_74_78 R_bl
Rbb_74_77 bitb_74_77 bitb_74_78 R_bl
Cb_74_77 bit_74_77 gnd C_bl
Cbb_74_77 bitb_74_77 gnd C_bl
Rb_74_78 bit_74_78 bit_74_79 R_bl
Rbb_74_78 bitb_74_78 bitb_74_79 R_bl
Cb_74_78 bit_74_78 gnd C_bl
Cbb_74_78 bitb_74_78 gnd C_bl
Rb_74_79 bit_74_79 bit_74_80 R_bl
Rbb_74_79 bitb_74_79 bitb_74_80 R_bl
Cb_74_79 bit_74_79 gnd C_bl
Cbb_74_79 bitb_74_79 gnd C_bl
Rb_74_80 bit_74_80 bit_74_81 R_bl
Rbb_74_80 bitb_74_80 bitb_74_81 R_bl
Cb_74_80 bit_74_80 gnd C_bl
Cbb_74_80 bitb_74_80 gnd C_bl
Rb_74_81 bit_74_81 bit_74_82 R_bl
Rbb_74_81 bitb_74_81 bitb_74_82 R_bl
Cb_74_81 bit_74_81 gnd C_bl
Cbb_74_81 bitb_74_81 gnd C_bl
Rb_74_82 bit_74_82 bit_74_83 R_bl
Rbb_74_82 bitb_74_82 bitb_74_83 R_bl
Cb_74_82 bit_74_82 gnd C_bl
Cbb_74_82 bitb_74_82 gnd C_bl
Rb_74_83 bit_74_83 bit_74_84 R_bl
Rbb_74_83 bitb_74_83 bitb_74_84 R_bl
Cb_74_83 bit_74_83 gnd C_bl
Cbb_74_83 bitb_74_83 gnd C_bl
Rb_74_84 bit_74_84 bit_74_85 R_bl
Rbb_74_84 bitb_74_84 bitb_74_85 R_bl
Cb_74_84 bit_74_84 gnd C_bl
Cbb_74_84 bitb_74_84 gnd C_bl
Rb_74_85 bit_74_85 bit_74_86 R_bl
Rbb_74_85 bitb_74_85 bitb_74_86 R_bl
Cb_74_85 bit_74_85 gnd C_bl
Cbb_74_85 bitb_74_85 gnd C_bl
Rb_74_86 bit_74_86 bit_74_87 R_bl
Rbb_74_86 bitb_74_86 bitb_74_87 R_bl
Cb_74_86 bit_74_86 gnd C_bl
Cbb_74_86 bitb_74_86 gnd C_bl
Rb_74_87 bit_74_87 bit_74_88 R_bl
Rbb_74_87 bitb_74_87 bitb_74_88 R_bl
Cb_74_87 bit_74_87 gnd C_bl
Cbb_74_87 bitb_74_87 gnd C_bl
Rb_74_88 bit_74_88 bit_74_89 R_bl
Rbb_74_88 bitb_74_88 bitb_74_89 R_bl
Cb_74_88 bit_74_88 gnd C_bl
Cbb_74_88 bitb_74_88 gnd C_bl
Rb_74_89 bit_74_89 bit_74_90 R_bl
Rbb_74_89 bitb_74_89 bitb_74_90 R_bl
Cb_74_89 bit_74_89 gnd C_bl
Cbb_74_89 bitb_74_89 gnd C_bl
Rb_74_90 bit_74_90 bit_74_91 R_bl
Rbb_74_90 bitb_74_90 bitb_74_91 R_bl
Cb_74_90 bit_74_90 gnd C_bl
Cbb_74_90 bitb_74_90 gnd C_bl
Rb_74_91 bit_74_91 bit_74_92 R_bl
Rbb_74_91 bitb_74_91 bitb_74_92 R_bl
Cb_74_91 bit_74_91 gnd C_bl
Cbb_74_91 bitb_74_91 gnd C_bl
Rb_74_92 bit_74_92 bit_74_93 R_bl
Rbb_74_92 bitb_74_92 bitb_74_93 R_bl
Cb_74_92 bit_74_92 gnd C_bl
Cbb_74_92 bitb_74_92 gnd C_bl
Rb_74_93 bit_74_93 bit_74_94 R_bl
Rbb_74_93 bitb_74_93 bitb_74_94 R_bl
Cb_74_93 bit_74_93 gnd C_bl
Cbb_74_93 bitb_74_93 gnd C_bl
Rb_74_94 bit_74_94 bit_74_95 R_bl
Rbb_74_94 bitb_74_94 bitb_74_95 R_bl
Cb_74_94 bit_74_94 gnd C_bl
Cbb_74_94 bitb_74_94 gnd C_bl
Rb_74_95 bit_74_95 bit_74_96 R_bl
Rbb_74_95 bitb_74_95 bitb_74_96 R_bl
Cb_74_95 bit_74_95 gnd C_bl
Cbb_74_95 bitb_74_95 gnd C_bl
Rb_74_96 bit_74_96 bit_74_97 R_bl
Rbb_74_96 bitb_74_96 bitb_74_97 R_bl
Cb_74_96 bit_74_96 gnd C_bl
Cbb_74_96 bitb_74_96 gnd C_bl
Rb_74_97 bit_74_97 bit_74_98 R_bl
Rbb_74_97 bitb_74_97 bitb_74_98 R_bl
Cb_74_97 bit_74_97 gnd C_bl
Cbb_74_97 bitb_74_97 gnd C_bl
Rb_74_98 bit_74_98 bit_74_99 R_bl
Rbb_74_98 bitb_74_98 bitb_74_99 R_bl
Cb_74_98 bit_74_98 gnd C_bl
Cbb_74_98 bitb_74_98 gnd C_bl
Rb_74_99 bit_74_99 bit_74_100 R_bl
Rbb_74_99 bitb_74_99 bitb_74_100 R_bl
Cb_74_99 bit_74_99 gnd C_bl
Cbb_74_99 bitb_74_99 gnd C_bl
Rb_75_0 bit_75_0 bit_75_1 R_bl
Rbb_75_0 bitb_75_0 bitb_75_1 R_bl
Cb_75_0 bit_75_0 gnd C_bl
Cbb_75_0 bitb_75_0 gnd C_bl
Rb_75_1 bit_75_1 bit_75_2 R_bl
Rbb_75_1 bitb_75_1 bitb_75_2 R_bl
Cb_75_1 bit_75_1 gnd C_bl
Cbb_75_1 bitb_75_1 gnd C_bl
Rb_75_2 bit_75_2 bit_75_3 R_bl
Rbb_75_2 bitb_75_2 bitb_75_3 R_bl
Cb_75_2 bit_75_2 gnd C_bl
Cbb_75_2 bitb_75_2 gnd C_bl
Rb_75_3 bit_75_3 bit_75_4 R_bl
Rbb_75_3 bitb_75_3 bitb_75_4 R_bl
Cb_75_3 bit_75_3 gnd C_bl
Cbb_75_3 bitb_75_3 gnd C_bl
Rb_75_4 bit_75_4 bit_75_5 R_bl
Rbb_75_4 bitb_75_4 bitb_75_5 R_bl
Cb_75_4 bit_75_4 gnd C_bl
Cbb_75_4 bitb_75_4 gnd C_bl
Rb_75_5 bit_75_5 bit_75_6 R_bl
Rbb_75_5 bitb_75_5 bitb_75_6 R_bl
Cb_75_5 bit_75_5 gnd C_bl
Cbb_75_5 bitb_75_5 gnd C_bl
Rb_75_6 bit_75_6 bit_75_7 R_bl
Rbb_75_6 bitb_75_6 bitb_75_7 R_bl
Cb_75_6 bit_75_6 gnd C_bl
Cbb_75_6 bitb_75_6 gnd C_bl
Rb_75_7 bit_75_7 bit_75_8 R_bl
Rbb_75_7 bitb_75_7 bitb_75_8 R_bl
Cb_75_7 bit_75_7 gnd C_bl
Cbb_75_7 bitb_75_7 gnd C_bl
Rb_75_8 bit_75_8 bit_75_9 R_bl
Rbb_75_8 bitb_75_8 bitb_75_9 R_bl
Cb_75_8 bit_75_8 gnd C_bl
Cbb_75_8 bitb_75_8 gnd C_bl
Rb_75_9 bit_75_9 bit_75_10 R_bl
Rbb_75_9 bitb_75_9 bitb_75_10 R_bl
Cb_75_9 bit_75_9 gnd C_bl
Cbb_75_9 bitb_75_9 gnd C_bl
Rb_75_10 bit_75_10 bit_75_11 R_bl
Rbb_75_10 bitb_75_10 bitb_75_11 R_bl
Cb_75_10 bit_75_10 gnd C_bl
Cbb_75_10 bitb_75_10 gnd C_bl
Rb_75_11 bit_75_11 bit_75_12 R_bl
Rbb_75_11 bitb_75_11 bitb_75_12 R_bl
Cb_75_11 bit_75_11 gnd C_bl
Cbb_75_11 bitb_75_11 gnd C_bl
Rb_75_12 bit_75_12 bit_75_13 R_bl
Rbb_75_12 bitb_75_12 bitb_75_13 R_bl
Cb_75_12 bit_75_12 gnd C_bl
Cbb_75_12 bitb_75_12 gnd C_bl
Rb_75_13 bit_75_13 bit_75_14 R_bl
Rbb_75_13 bitb_75_13 bitb_75_14 R_bl
Cb_75_13 bit_75_13 gnd C_bl
Cbb_75_13 bitb_75_13 gnd C_bl
Rb_75_14 bit_75_14 bit_75_15 R_bl
Rbb_75_14 bitb_75_14 bitb_75_15 R_bl
Cb_75_14 bit_75_14 gnd C_bl
Cbb_75_14 bitb_75_14 gnd C_bl
Rb_75_15 bit_75_15 bit_75_16 R_bl
Rbb_75_15 bitb_75_15 bitb_75_16 R_bl
Cb_75_15 bit_75_15 gnd C_bl
Cbb_75_15 bitb_75_15 gnd C_bl
Rb_75_16 bit_75_16 bit_75_17 R_bl
Rbb_75_16 bitb_75_16 bitb_75_17 R_bl
Cb_75_16 bit_75_16 gnd C_bl
Cbb_75_16 bitb_75_16 gnd C_bl
Rb_75_17 bit_75_17 bit_75_18 R_bl
Rbb_75_17 bitb_75_17 bitb_75_18 R_bl
Cb_75_17 bit_75_17 gnd C_bl
Cbb_75_17 bitb_75_17 gnd C_bl
Rb_75_18 bit_75_18 bit_75_19 R_bl
Rbb_75_18 bitb_75_18 bitb_75_19 R_bl
Cb_75_18 bit_75_18 gnd C_bl
Cbb_75_18 bitb_75_18 gnd C_bl
Rb_75_19 bit_75_19 bit_75_20 R_bl
Rbb_75_19 bitb_75_19 bitb_75_20 R_bl
Cb_75_19 bit_75_19 gnd C_bl
Cbb_75_19 bitb_75_19 gnd C_bl
Rb_75_20 bit_75_20 bit_75_21 R_bl
Rbb_75_20 bitb_75_20 bitb_75_21 R_bl
Cb_75_20 bit_75_20 gnd C_bl
Cbb_75_20 bitb_75_20 gnd C_bl
Rb_75_21 bit_75_21 bit_75_22 R_bl
Rbb_75_21 bitb_75_21 bitb_75_22 R_bl
Cb_75_21 bit_75_21 gnd C_bl
Cbb_75_21 bitb_75_21 gnd C_bl
Rb_75_22 bit_75_22 bit_75_23 R_bl
Rbb_75_22 bitb_75_22 bitb_75_23 R_bl
Cb_75_22 bit_75_22 gnd C_bl
Cbb_75_22 bitb_75_22 gnd C_bl
Rb_75_23 bit_75_23 bit_75_24 R_bl
Rbb_75_23 bitb_75_23 bitb_75_24 R_bl
Cb_75_23 bit_75_23 gnd C_bl
Cbb_75_23 bitb_75_23 gnd C_bl
Rb_75_24 bit_75_24 bit_75_25 R_bl
Rbb_75_24 bitb_75_24 bitb_75_25 R_bl
Cb_75_24 bit_75_24 gnd C_bl
Cbb_75_24 bitb_75_24 gnd C_bl
Rb_75_25 bit_75_25 bit_75_26 R_bl
Rbb_75_25 bitb_75_25 bitb_75_26 R_bl
Cb_75_25 bit_75_25 gnd C_bl
Cbb_75_25 bitb_75_25 gnd C_bl
Rb_75_26 bit_75_26 bit_75_27 R_bl
Rbb_75_26 bitb_75_26 bitb_75_27 R_bl
Cb_75_26 bit_75_26 gnd C_bl
Cbb_75_26 bitb_75_26 gnd C_bl
Rb_75_27 bit_75_27 bit_75_28 R_bl
Rbb_75_27 bitb_75_27 bitb_75_28 R_bl
Cb_75_27 bit_75_27 gnd C_bl
Cbb_75_27 bitb_75_27 gnd C_bl
Rb_75_28 bit_75_28 bit_75_29 R_bl
Rbb_75_28 bitb_75_28 bitb_75_29 R_bl
Cb_75_28 bit_75_28 gnd C_bl
Cbb_75_28 bitb_75_28 gnd C_bl
Rb_75_29 bit_75_29 bit_75_30 R_bl
Rbb_75_29 bitb_75_29 bitb_75_30 R_bl
Cb_75_29 bit_75_29 gnd C_bl
Cbb_75_29 bitb_75_29 gnd C_bl
Rb_75_30 bit_75_30 bit_75_31 R_bl
Rbb_75_30 bitb_75_30 bitb_75_31 R_bl
Cb_75_30 bit_75_30 gnd C_bl
Cbb_75_30 bitb_75_30 gnd C_bl
Rb_75_31 bit_75_31 bit_75_32 R_bl
Rbb_75_31 bitb_75_31 bitb_75_32 R_bl
Cb_75_31 bit_75_31 gnd C_bl
Cbb_75_31 bitb_75_31 gnd C_bl
Rb_75_32 bit_75_32 bit_75_33 R_bl
Rbb_75_32 bitb_75_32 bitb_75_33 R_bl
Cb_75_32 bit_75_32 gnd C_bl
Cbb_75_32 bitb_75_32 gnd C_bl
Rb_75_33 bit_75_33 bit_75_34 R_bl
Rbb_75_33 bitb_75_33 bitb_75_34 R_bl
Cb_75_33 bit_75_33 gnd C_bl
Cbb_75_33 bitb_75_33 gnd C_bl
Rb_75_34 bit_75_34 bit_75_35 R_bl
Rbb_75_34 bitb_75_34 bitb_75_35 R_bl
Cb_75_34 bit_75_34 gnd C_bl
Cbb_75_34 bitb_75_34 gnd C_bl
Rb_75_35 bit_75_35 bit_75_36 R_bl
Rbb_75_35 bitb_75_35 bitb_75_36 R_bl
Cb_75_35 bit_75_35 gnd C_bl
Cbb_75_35 bitb_75_35 gnd C_bl
Rb_75_36 bit_75_36 bit_75_37 R_bl
Rbb_75_36 bitb_75_36 bitb_75_37 R_bl
Cb_75_36 bit_75_36 gnd C_bl
Cbb_75_36 bitb_75_36 gnd C_bl
Rb_75_37 bit_75_37 bit_75_38 R_bl
Rbb_75_37 bitb_75_37 bitb_75_38 R_bl
Cb_75_37 bit_75_37 gnd C_bl
Cbb_75_37 bitb_75_37 gnd C_bl
Rb_75_38 bit_75_38 bit_75_39 R_bl
Rbb_75_38 bitb_75_38 bitb_75_39 R_bl
Cb_75_38 bit_75_38 gnd C_bl
Cbb_75_38 bitb_75_38 gnd C_bl
Rb_75_39 bit_75_39 bit_75_40 R_bl
Rbb_75_39 bitb_75_39 bitb_75_40 R_bl
Cb_75_39 bit_75_39 gnd C_bl
Cbb_75_39 bitb_75_39 gnd C_bl
Rb_75_40 bit_75_40 bit_75_41 R_bl
Rbb_75_40 bitb_75_40 bitb_75_41 R_bl
Cb_75_40 bit_75_40 gnd C_bl
Cbb_75_40 bitb_75_40 gnd C_bl
Rb_75_41 bit_75_41 bit_75_42 R_bl
Rbb_75_41 bitb_75_41 bitb_75_42 R_bl
Cb_75_41 bit_75_41 gnd C_bl
Cbb_75_41 bitb_75_41 gnd C_bl
Rb_75_42 bit_75_42 bit_75_43 R_bl
Rbb_75_42 bitb_75_42 bitb_75_43 R_bl
Cb_75_42 bit_75_42 gnd C_bl
Cbb_75_42 bitb_75_42 gnd C_bl
Rb_75_43 bit_75_43 bit_75_44 R_bl
Rbb_75_43 bitb_75_43 bitb_75_44 R_bl
Cb_75_43 bit_75_43 gnd C_bl
Cbb_75_43 bitb_75_43 gnd C_bl
Rb_75_44 bit_75_44 bit_75_45 R_bl
Rbb_75_44 bitb_75_44 bitb_75_45 R_bl
Cb_75_44 bit_75_44 gnd C_bl
Cbb_75_44 bitb_75_44 gnd C_bl
Rb_75_45 bit_75_45 bit_75_46 R_bl
Rbb_75_45 bitb_75_45 bitb_75_46 R_bl
Cb_75_45 bit_75_45 gnd C_bl
Cbb_75_45 bitb_75_45 gnd C_bl
Rb_75_46 bit_75_46 bit_75_47 R_bl
Rbb_75_46 bitb_75_46 bitb_75_47 R_bl
Cb_75_46 bit_75_46 gnd C_bl
Cbb_75_46 bitb_75_46 gnd C_bl
Rb_75_47 bit_75_47 bit_75_48 R_bl
Rbb_75_47 bitb_75_47 bitb_75_48 R_bl
Cb_75_47 bit_75_47 gnd C_bl
Cbb_75_47 bitb_75_47 gnd C_bl
Rb_75_48 bit_75_48 bit_75_49 R_bl
Rbb_75_48 bitb_75_48 bitb_75_49 R_bl
Cb_75_48 bit_75_48 gnd C_bl
Cbb_75_48 bitb_75_48 gnd C_bl
Rb_75_49 bit_75_49 bit_75_50 R_bl
Rbb_75_49 bitb_75_49 bitb_75_50 R_bl
Cb_75_49 bit_75_49 gnd C_bl
Cbb_75_49 bitb_75_49 gnd C_bl
Rb_75_50 bit_75_50 bit_75_51 R_bl
Rbb_75_50 bitb_75_50 bitb_75_51 R_bl
Cb_75_50 bit_75_50 gnd C_bl
Cbb_75_50 bitb_75_50 gnd C_bl
Rb_75_51 bit_75_51 bit_75_52 R_bl
Rbb_75_51 bitb_75_51 bitb_75_52 R_bl
Cb_75_51 bit_75_51 gnd C_bl
Cbb_75_51 bitb_75_51 gnd C_bl
Rb_75_52 bit_75_52 bit_75_53 R_bl
Rbb_75_52 bitb_75_52 bitb_75_53 R_bl
Cb_75_52 bit_75_52 gnd C_bl
Cbb_75_52 bitb_75_52 gnd C_bl
Rb_75_53 bit_75_53 bit_75_54 R_bl
Rbb_75_53 bitb_75_53 bitb_75_54 R_bl
Cb_75_53 bit_75_53 gnd C_bl
Cbb_75_53 bitb_75_53 gnd C_bl
Rb_75_54 bit_75_54 bit_75_55 R_bl
Rbb_75_54 bitb_75_54 bitb_75_55 R_bl
Cb_75_54 bit_75_54 gnd C_bl
Cbb_75_54 bitb_75_54 gnd C_bl
Rb_75_55 bit_75_55 bit_75_56 R_bl
Rbb_75_55 bitb_75_55 bitb_75_56 R_bl
Cb_75_55 bit_75_55 gnd C_bl
Cbb_75_55 bitb_75_55 gnd C_bl
Rb_75_56 bit_75_56 bit_75_57 R_bl
Rbb_75_56 bitb_75_56 bitb_75_57 R_bl
Cb_75_56 bit_75_56 gnd C_bl
Cbb_75_56 bitb_75_56 gnd C_bl
Rb_75_57 bit_75_57 bit_75_58 R_bl
Rbb_75_57 bitb_75_57 bitb_75_58 R_bl
Cb_75_57 bit_75_57 gnd C_bl
Cbb_75_57 bitb_75_57 gnd C_bl
Rb_75_58 bit_75_58 bit_75_59 R_bl
Rbb_75_58 bitb_75_58 bitb_75_59 R_bl
Cb_75_58 bit_75_58 gnd C_bl
Cbb_75_58 bitb_75_58 gnd C_bl
Rb_75_59 bit_75_59 bit_75_60 R_bl
Rbb_75_59 bitb_75_59 bitb_75_60 R_bl
Cb_75_59 bit_75_59 gnd C_bl
Cbb_75_59 bitb_75_59 gnd C_bl
Rb_75_60 bit_75_60 bit_75_61 R_bl
Rbb_75_60 bitb_75_60 bitb_75_61 R_bl
Cb_75_60 bit_75_60 gnd C_bl
Cbb_75_60 bitb_75_60 gnd C_bl
Rb_75_61 bit_75_61 bit_75_62 R_bl
Rbb_75_61 bitb_75_61 bitb_75_62 R_bl
Cb_75_61 bit_75_61 gnd C_bl
Cbb_75_61 bitb_75_61 gnd C_bl
Rb_75_62 bit_75_62 bit_75_63 R_bl
Rbb_75_62 bitb_75_62 bitb_75_63 R_bl
Cb_75_62 bit_75_62 gnd C_bl
Cbb_75_62 bitb_75_62 gnd C_bl
Rb_75_63 bit_75_63 bit_75_64 R_bl
Rbb_75_63 bitb_75_63 bitb_75_64 R_bl
Cb_75_63 bit_75_63 gnd C_bl
Cbb_75_63 bitb_75_63 gnd C_bl
Rb_75_64 bit_75_64 bit_75_65 R_bl
Rbb_75_64 bitb_75_64 bitb_75_65 R_bl
Cb_75_64 bit_75_64 gnd C_bl
Cbb_75_64 bitb_75_64 gnd C_bl
Rb_75_65 bit_75_65 bit_75_66 R_bl
Rbb_75_65 bitb_75_65 bitb_75_66 R_bl
Cb_75_65 bit_75_65 gnd C_bl
Cbb_75_65 bitb_75_65 gnd C_bl
Rb_75_66 bit_75_66 bit_75_67 R_bl
Rbb_75_66 bitb_75_66 bitb_75_67 R_bl
Cb_75_66 bit_75_66 gnd C_bl
Cbb_75_66 bitb_75_66 gnd C_bl
Rb_75_67 bit_75_67 bit_75_68 R_bl
Rbb_75_67 bitb_75_67 bitb_75_68 R_bl
Cb_75_67 bit_75_67 gnd C_bl
Cbb_75_67 bitb_75_67 gnd C_bl
Rb_75_68 bit_75_68 bit_75_69 R_bl
Rbb_75_68 bitb_75_68 bitb_75_69 R_bl
Cb_75_68 bit_75_68 gnd C_bl
Cbb_75_68 bitb_75_68 gnd C_bl
Rb_75_69 bit_75_69 bit_75_70 R_bl
Rbb_75_69 bitb_75_69 bitb_75_70 R_bl
Cb_75_69 bit_75_69 gnd C_bl
Cbb_75_69 bitb_75_69 gnd C_bl
Rb_75_70 bit_75_70 bit_75_71 R_bl
Rbb_75_70 bitb_75_70 bitb_75_71 R_bl
Cb_75_70 bit_75_70 gnd C_bl
Cbb_75_70 bitb_75_70 gnd C_bl
Rb_75_71 bit_75_71 bit_75_72 R_bl
Rbb_75_71 bitb_75_71 bitb_75_72 R_bl
Cb_75_71 bit_75_71 gnd C_bl
Cbb_75_71 bitb_75_71 gnd C_bl
Rb_75_72 bit_75_72 bit_75_73 R_bl
Rbb_75_72 bitb_75_72 bitb_75_73 R_bl
Cb_75_72 bit_75_72 gnd C_bl
Cbb_75_72 bitb_75_72 gnd C_bl
Rb_75_73 bit_75_73 bit_75_74 R_bl
Rbb_75_73 bitb_75_73 bitb_75_74 R_bl
Cb_75_73 bit_75_73 gnd C_bl
Cbb_75_73 bitb_75_73 gnd C_bl
Rb_75_74 bit_75_74 bit_75_75 R_bl
Rbb_75_74 bitb_75_74 bitb_75_75 R_bl
Cb_75_74 bit_75_74 gnd C_bl
Cbb_75_74 bitb_75_74 gnd C_bl
Rb_75_75 bit_75_75 bit_75_76 R_bl
Rbb_75_75 bitb_75_75 bitb_75_76 R_bl
Cb_75_75 bit_75_75 gnd C_bl
Cbb_75_75 bitb_75_75 gnd C_bl
Rb_75_76 bit_75_76 bit_75_77 R_bl
Rbb_75_76 bitb_75_76 bitb_75_77 R_bl
Cb_75_76 bit_75_76 gnd C_bl
Cbb_75_76 bitb_75_76 gnd C_bl
Rb_75_77 bit_75_77 bit_75_78 R_bl
Rbb_75_77 bitb_75_77 bitb_75_78 R_bl
Cb_75_77 bit_75_77 gnd C_bl
Cbb_75_77 bitb_75_77 gnd C_bl
Rb_75_78 bit_75_78 bit_75_79 R_bl
Rbb_75_78 bitb_75_78 bitb_75_79 R_bl
Cb_75_78 bit_75_78 gnd C_bl
Cbb_75_78 bitb_75_78 gnd C_bl
Rb_75_79 bit_75_79 bit_75_80 R_bl
Rbb_75_79 bitb_75_79 bitb_75_80 R_bl
Cb_75_79 bit_75_79 gnd C_bl
Cbb_75_79 bitb_75_79 gnd C_bl
Rb_75_80 bit_75_80 bit_75_81 R_bl
Rbb_75_80 bitb_75_80 bitb_75_81 R_bl
Cb_75_80 bit_75_80 gnd C_bl
Cbb_75_80 bitb_75_80 gnd C_bl
Rb_75_81 bit_75_81 bit_75_82 R_bl
Rbb_75_81 bitb_75_81 bitb_75_82 R_bl
Cb_75_81 bit_75_81 gnd C_bl
Cbb_75_81 bitb_75_81 gnd C_bl
Rb_75_82 bit_75_82 bit_75_83 R_bl
Rbb_75_82 bitb_75_82 bitb_75_83 R_bl
Cb_75_82 bit_75_82 gnd C_bl
Cbb_75_82 bitb_75_82 gnd C_bl
Rb_75_83 bit_75_83 bit_75_84 R_bl
Rbb_75_83 bitb_75_83 bitb_75_84 R_bl
Cb_75_83 bit_75_83 gnd C_bl
Cbb_75_83 bitb_75_83 gnd C_bl
Rb_75_84 bit_75_84 bit_75_85 R_bl
Rbb_75_84 bitb_75_84 bitb_75_85 R_bl
Cb_75_84 bit_75_84 gnd C_bl
Cbb_75_84 bitb_75_84 gnd C_bl
Rb_75_85 bit_75_85 bit_75_86 R_bl
Rbb_75_85 bitb_75_85 bitb_75_86 R_bl
Cb_75_85 bit_75_85 gnd C_bl
Cbb_75_85 bitb_75_85 gnd C_bl
Rb_75_86 bit_75_86 bit_75_87 R_bl
Rbb_75_86 bitb_75_86 bitb_75_87 R_bl
Cb_75_86 bit_75_86 gnd C_bl
Cbb_75_86 bitb_75_86 gnd C_bl
Rb_75_87 bit_75_87 bit_75_88 R_bl
Rbb_75_87 bitb_75_87 bitb_75_88 R_bl
Cb_75_87 bit_75_87 gnd C_bl
Cbb_75_87 bitb_75_87 gnd C_bl
Rb_75_88 bit_75_88 bit_75_89 R_bl
Rbb_75_88 bitb_75_88 bitb_75_89 R_bl
Cb_75_88 bit_75_88 gnd C_bl
Cbb_75_88 bitb_75_88 gnd C_bl
Rb_75_89 bit_75_89 bit_75_90 R_bl
Rbb_75_89 bitb_75_89 bitb_75_90 R_bl
Cb_75_89 bit_75_89 gnd C_bl
Cbb_75_89 bitb_75_89 gnd C_bl
Rb_75_90 bit_75_90 bit_75_91 R_bl
Rbb_75_90 bitb_75_90 bitb_75_91 R_bl
Cb_75_90 bit_75_90 gnd C_bl
Cbb_75_90 bitb_75_90 gnd C_bl
Rb_75_91 bit_75_91 bit_75_92 R_bl
Rbb_75_91 bitb_75_91 bitb_75_92 R_bl
Cb_75_91 bit_75_91 gnd C_bl
Cbb_75_91 bitb_75_91 gnd C_bl
Rb_75_92 bit_75_92 bit_75_93 R_bl
Rbb_75_92 bitb_75_92 bitb_75_93 R_bl
Cb_75_92 bit_75_92 gnd C_bl
Cbb_75_92 bitb_75_92 gnd C_bl
Rb_75_93 bit_75_93 bit_75_94 R_bl
Rbb_75_93 bitb_75_93 bitb_75_94 R_bl
Cb_75_93 bit_75_93 gnd C_bl
Cbb_75_93 bitb_75_93 gnd C_bl
Rb_75_94 bit_75_94 bit_75_95 R_bl
Rbb_75_94 bitb_75_94 bitb_75_95 R_bl
Cb_75_94 bit_75_94 gnd C_bl
Cbb_75_94 bitb_75_94 gnd C_bl
Rb_75_95 bit_75_95 bit_75_96 R_bl
Rbb_75_95 bitb_75_95 bitb_75_96 R_bl
Cb_75_95 bit_75_95 gnd C_bl
Cbb_75_95 bitb_75_95 gnd C_bl
Rb_75_96 bit_75_96 bit_75_97 R_bl
Rbb_75_96 bitb_75_96 bitb_75_97 R_bl
Cb_75_96 bit_75_96 gnd C_bl
Cbb_75_96 bitb_75_96 gnd C_bl
Rb_75_97 bit_75_97 bit_75_98 R_bl
Rbb_75_97 bitb_75_97 bitb_75_98 R_bl
Cb_75_97 bit_75_97 gnd C_bl
Cbb_75_97 bitb_75_97 gnd C_bl
Rb_75_98 bit_75_98 bit_75_99 R_bl
Rbb_75_98 bitb_75_98 bitb_75_99 R_bl
Cb_75_98 bit_75_98 gnd C_bl
Cbb_75_98 bitb_75_98 gnd C_bl
Rb_75_99 bit_75_99 bit_75_100 R_bl
Rbb_75_99 bitb_75_99 bitb_75_100 R_bl
Cb_75_99 bit_75_99 gnd C_bl
Cbb_75_99 bitb_75_99 gnd C_bl
Rb_76_0 bit_76_0 bit_76_1 R_bl
Rbb_76_0 bitb_76_0 bitb_76_1 R_bl
Cb_76_0 bit_76_0 gnd C_bl
Cbb_76_0 bitb_76_0 gnd C_bl
Rb_76_1 bit_76_1 bit_76_2 R_bl
Rbb_76_1 bitb_76_1 bitb_76_2 R_bl
Cb_76_1 bit_76_1 gnd C_bl
Cbb_76_1 bitb_76_1 gnd C_bl
Rb_76_2 bit_76_2 bit_76_3 R_bl
Rbb_76_2 bitb_76_2 bitb_76_3 R_bl
Cb_76_2 bit_76_2 gnd C_bl
Cbb_76_2 bitb_76_2 gnd C_bl
Rb_76_3 bit_76_3 bit_76_4 R_bl
Rbb_76_3 bitb_76_3 bitb_76_4 R_bl
Cb_76_3 bit_76_3 gnd C_bl
Cbb_76_3 bitb_76_3 gnd C_bl
Rb_76_4 bit_76_4 bit_76_5 R_bl
Rbb_76_4 bitb_76_4 bitb_76_5 R_bl
Cb_76_4 bit_76_4 gnd C_bl
Cbb_76_4 bitb_76_4 gnd C_bl
Rb_76_5 bit_76_5 bit_76_6 R_bl
Rbb_76_5 bitb_76_5 bitb_76_6 R_bl
Cb_76_5 bit_76_5 gnd C_bl
Cbb_76_5 bitb_76_5 gnd C_bl
Rb_76_6 bit_76_6 bit_76_7 R_bl
Rbb_76_6 bitb_76_6 bitb_76_7 R_bl
Cb_76_6 bit_76_6 gnd C_bl
Cbb_76_6 bitb_76_6 gnd C_bl
Rb_76_7 bit_76_7 bit_76_8 R_bl
Rbb_76_7 bitb_76_7 bitb_76_8 R_bl
Cb_76_7 bit_76_7 gnd C_bl
Cbb_76_7 bitb_76_7 gnd C_bl
Rb_76_8 bit_76_8 bit_76_9 R_bl
Rbb_76_8 bitb_76_8 bitb_76_9 R_bl
Cb_76_8 bit_76_8 gnd C_bl
Cbb_76_8 bitb_76_8 gnd C_bl
Rb_76_9 bit_76_9 bit_76_10 R_bl
Rbb_76_9 bitb_76_9 bitb_76_10 R_bl
Cb_76_9 bit_76_9 gnd C_bl
Cbb_76_9 bitb_76_9 gnd C_bl
Rb_76_10 bit_76_10 bit_76_11 R_bl
Rbb_76_10 bitb_76_10 bitb_76_11 R_bl
Cb_76_10 bit_76_10 gnd C_bl
Cbb_76_10 bitb_76_10 gnd C_bl
Rb_76_11 bit_76_11 bit_76_12 R_bl
Rbb_76_11 bitb_76_11 bitb_76_12 R_bl
Cb_76_11 bit_76_11 gnd C_bl
Cbb_76_11 bitb_76_11 gnd C_bl
Rb_76_12 bit_76_12 bit_76_13 R_bl
Rbb_76_12 bitb_76_12 bitb_76_13 R_bl
Cb_76_12 bit_76_12 gnd C_bl
Cbb_76_12 bitb_76_12 gnd C_bl
Rb_76_13 bit_76_13 bit_76_14 R_bl
Rbb_76_13 bitb_76_13 bitb_76_14 R_bl
Cb_76_13 bit_76_13 gnd C_bl
Cbb_76_13 bitb_76_13 gnd C_bl
Rb_76_14 bit_76_14 bit_76_15 R_bl
Rbb_76_14 bitb_76_14 bitb_76_15 R_bl
Cb_76_14 bit_76_14 gnd C_bl
Cbb_76_14 bitb_76_14 gnd C_bl
Rb_76_15 bit_76_15 bit_76_16 R_bl
Rbb_76_15 bitb_76_15 bitb_76_16 R_bl
Cb_76_15 bit_76_15 gnd C_bl
Cbb_76_15 bitb_76_15 gnd C_bl
Rb_76_16 bit_76_16 bit_76_17 R_bl
Rbb_76_16 bitb_76_16 bitb_76_17 R_bl
Cb_76_16 bit_76_16 gnd C_bl
Cbb_76_16 bitb_76_16 gnd C_bl
Rb_76_17 bit_76_17 bit_76_18 R_bl
Rbb_76_17 bitb_76_17 bitb_76_18 R_bl
Cb_76_17 bit_76_17 gnd C_bl
Cbb_76_17 bitb_76_17 gnd C_bl
Rb_76_18 bit_76_18 bit_76_19 R_bl
Rbb_76_18 bitb_76_18 bitb_76_19 R_bl
Cb_76_18 bit_76_18 gnd C_bl
Cbb_76_18 bitb_76_18 gnd C_bl
Rb_76_19 bit_76_19 bit_76_20 R_bl
Rbb_76_19 bitb_76_19 bitb_76_20 R_bl
Cb_76_19 bit_76_19 gnd C_bl
Cbb_76_19 bitb_76_19 gnd C_bl
Rb_76_20 bit_76_20 bit_76_21 R_bl
Rbb_76_20 bitb_76_20 bitb_76_21 R_bl
Cb_76_20 bit_76_20 gnd C_bl
Cbb_76_20 bitb_76_20 gnd C_bl
Rb_76_21 bit_76_21 bit_76_22 R_bl
Rbb_76_21 bitb_76_21 bitb_76_22 R_bl
Cb_76_21 bit_76_21 gnd C_bl
Cbb_76_21 bitb_76_21 gnd C_bl
Rb_76_22 bit_76_22 bit_76_23 R_bl
Rbb_76_22 bitb_76_22 bitb_76_23 R_bl
Cb_76_22 bit_76_22 gnd C_bl
Cbb_76_22 bitb_76_22 gnd C_bl
Rb_76_23 bit_76_23 bit_76_24 R_bl
Rbb_76_23 bitb_76_23 bitb_76_24 R_bl
Cb_76_23 bit_76_23 gnd C_bl
Cbb_76_23 bitb_76_23 gnd C_bl
Rb_76_24 bit_76_24 bit_76_25 R_bl
Rbb_76_24 bitb_76_24 bitb_76_25 R_bl
Cb_76_24 bit_76_24 gnd C_bl
Cbb_76_24 bitb_76_24 gnd C_bl
Rb_76_25 bit_76_25 bit_76_26 R_bl
Rbb_76_25 bitb_76_25 bitb_76_26 R_bl
Cb_76_25 bit_76_25 gnd C_bl
Cbb_76_25 bitb_76_25 gnd C_bl
Rb_76_26 bit_76_26 bit_76_27 R_bl
Rbb_76_26 bitb_76_26 bitb_76_27 R_bl
Cb_76_26 bit_76_26 gnd C_bl
Cbb_76_26 bitb_76_26 gnd C_bl
Rb_76_27 bit_76_27 bit_76_28 R_bl
Rbb_76_27 bitb_76_27 bitb_76_28 R_bl
Cb_76_27 bit_76_27 gnd C_bl
Cbb_76_27 bitb_76_27 gnd C_bl
Rb_76_28 bit_76_28 bit_76_29 R_bl
Rbb_76_28 bitb_76_28 bitb_76_29 R_bl
Cb_76_28 bit_76_28 gnd C_bl
Cbb_76_28 bitb_76_28 gnd C_bl
Rb_76_29 bit_76_29 bit_76_30 R_bl
Rbb_76_29 bitb_76_29 bitb_76_30 R_bl
Cb_76_29 bit_76_29 gnd C_bl
Cbb_76_29 bitb_76_29 gnd C_bl
Rb_76_30 bit_76_30 bit_76_31 R_bl
Rbb_76_30 bitb_76_30 bitb_76_31 R_bl
Cb_76_30 bit_76_30 gnd C_bl
Cbb_76_30 bitb_76_30 gnd C_bl
Rb_76_31 bit_76_31 bit_76_32 R_bl
Rbb_76_31 bitb_76_31 bitb_76_32 R_bl
Cb_76_31 bit_76_31 gnd C_bl
Cbb_76_31 bitb_76_31 gnd C_bl
Rb_76_32 bit_76_32 bit_76_33 R_bl
Rbb_76_32 bitb_76_32 bitb_76_33 R_bl
Cb_76_32 bit_76_32 gnd C_bl
Cbb_76_32 bitb_76_32 gnd C_bl
Rb_76_33 bit_76_33 bit_76_34 R_bl
Rbb_76_33 bitb_76_33 bitb_76_34 R_bl
Cb_76_33 bit_76_33 gnd C_bl
Cbb_76_33 bitb_76_33 gnd C_bl
Rb_76_34 bit_76_34 bit_76_35 R_bl
Rbb_76_34 bitb_76_34 bitb_76_35 R_bl
Cb_76_34 bit_76_34 gnd C_bl
Cbb_76_34 bitb_76_34 gnd C_bl
Rb_76_35 bit_76_35 bit_76_36 R_bl
Rbb_76_35 bitb_76_35 bitb_76_36 R_bl
Cb_76_35 bit_76_35 gnd C_bl
Cbb_76_35 bitb_76_35 gnd C_bl
Rb_76_36 bit_76_36 bit_76_37 R_bl
Rbb_76_36 bitb_76_36 bitb_76_37 R_bl
Cb_76_36 bit_76_36 gnd C_bl
Cbb_76_36 bitb_76_36 gnd C_bl
Rb_76_37 bit_76_37 bit_76_38 R_bl
Rbb_76_37 bitb_76_37 bitb_76_38 R_bl
Cb_76_37 bit_76_37 gnd C_bl
Cbb_76_37 bitb_76_37 gnd C_bl
Rb_76_38 bit_76_38 bit_76_39 R_bl
Rbb_76_38 bitb_76_38 bitb_76_39 R_bl
Cb_76_38 bit_76_38 gnd C_bl
Cbb_76_38 bitb_76_38 gnd C_bl
Rb_76_39 bit_76_39 bit_76_40 R_bl
Rbb_76_39 bitb_76_39 bitb_76_40 R_bl
Cb_76_39 bit_76_39 gnd C_bl
Cbb_76_39 bitb_76_39 gnd C_bl
Rb_76_40 bit_76_40 bit_76_41 R_bl
Rbb_76_40 bitb_76_40 bitb_76_41 R_bl
Cb_76_40 bit_76_40 gnd C_bl
Cbb_76_40 bitb_76_40 gnd C_bl
Rb_76_41 bit_76_41 bit_76_42 R_bl
Rbb_76_41 bitb_76_41 bitb_76_42 R_bl
Cb_76_41 bit_76_41 gnd C_bl
Cbb_76_41 bitb_76_41 gnd C_bl
Rb_76_42 bit_76_42 bit_76_43 R_bl
Rbb_76_42 bitb_76_42 bitb_76_43 R_bl
Cb_76_42 bit_76_42 gnd C_bl
Cbb_76_42 bitb_76_42 gnd C_bl
Rb_76_43 bit_76_43 bit_76_44 R_bl
Rbb_76_43 bitb_76_43 bitb_76_44 R_bl
Cb_76_43 bit_76_43 gnd C_bl
Cbb_76_43 bitb_76_43 gnd C_bl
Rb_76_44 bit_76_44 bit_76_45 R_bl
Rbb_76_44 bitb_76_44 bitb_76_45 R_bl
Cb_76_44 bit_76_44 gnd C_bl
Cbb_76_44 bitb_76_44 gnd C_bl
Rb_76_45 bit_76_45 bit_76_46 R_bl
Rbb_76_45 bitb_76_45 bitb_76_46 R_bl
Cb_76_45 bit_76_45 gnd C_bl
Cbb_76_45 bitb_76_45 gnd C_bl
Rb_76_46 bit_76_46 bit_76_47 R_bl
Rbb_76_46 bitb_76_46 bitb_76_47 R_bl
Cb_76_46 bit_76_46 gnd C_bl
Cbb_76_46 bitb_76_46 gnd C_bl
Rb_76_47 bit_76_47 bit_76_48 R_bl
Rbb_76_47 bitb_76_47 bitb_76_48 R_bl
Cb_76_47 bit_76_47 gnd C_bl
Cbb_76_47 bitb_76_47 gnd C_bl
Rb_76_48 bit_76_48 bit_76_49 R_bl
Rbb_76_48 bitb_76_48 bitb_76_49 R_bl
Cb_76_48 bit_76_48 gnd C_bl
Cbb_76_48 bitb_76_48 gnd C_bl
Rb_76_49 bit_76_49 bit_76_50 R_bl
Rbb_76_49 bitb_76_49 bitb_76_50 R_bl
Cb_76_49 bit_76_49 gnd C_bl
Cbb_76_49 bitb_76_49 gnd C_bl
Rb_76_50 bit_76_50 bit_76_51 R_bl
Rbb_76_50 bitb_76_50 bitb_76_51 R_bl
Cb_76_50 bit_76_50 gnd C_bl
Cbb_76_50 bitb_76_50 gnd C_bl
Rb_76_51 bit_76_51 bit_76_52 R_bl
Rbb_76_51 bitb_76_51 bitb_76_52 R_bl
Cb_76_51 bit_76_51 gnd C_bl
Cbb_76_51 bitb_76_51 gnd C_bl
Rb_76_52 bit_76_52 bit_76_53 R_bl
Rbb_76_52 bitb_76_52 bitb_76_53 R_bl
Cb_76_52 bit_76_52 gnd C_bl
Cbb_76_52 bitb_76_52 gnd C_bl
Rb_76_53 bit_76_53 bit_76_54 R_bl
Rbb_76_53 bitb_76_53 bitb_76_54 R_bl
Cb_76_53 bit_76_53 gnd C_bl
Cbb_76_53 bitb_76_53 gnd C_bl
Rb_76_54 bit_76_54 bit_76_55 R_bl
Rbb_76_54 bitb_76_54 bitb_76_55 R_bl
Cb_76_54 bit_76_54 gnd C_bl
Cbb_76_54 bitb_76_54 gnd C_bl
Rb_76_55 bit_76_55 bit_76_56 R_bl
Rbb_76_55 bitb_76_55 bitb_76_56 R_bl
Cb_76_55 bit_76_55 gnd C_bl
Cbb_76_55 bitb_76_55 gnd C_bl
Rb_76_56 bit_76_56 bit_76_57 R_bl
Rbb_76_56 bitb_76_56 bitb_76_57 R_bl
Cb_76_56 bit_76_56 gnd C_bl
Cbb_76_56 bitb_76_56 gnd C_bl
Rb_76_57 bit_76_57 bit_76_58 R_bl
Rbb_76_57 bitb_76_57 bitb_76_58 R_bl
Cb_76_57 bit_76_57 gnd C_bl
Cbb_76_57 bitb_76_57 gnd C_bl
Rb_76_58 bit_76_58 bit_76_59 R_bl
Rbb_76_58 bitb_76_58 bitb_76_59 R_bl
Cb_76_58 bit_76_58 gnd C_bl
Cbb_76_58 bitb_76_58 gnd C_bl
Rb_76_59 bit_76_59 bit_76_60 R_bl
Rbb_76_59 bitb_76_59 bitb_76_60 R_bl
Cb_76_59 bit_76_59 gnd C_bl
Cbb_76_59 bitb_76_59 gnd C_bl
Rb_76_60 bit_76_60 bit_76_61 R_bl
Rbb_76_60 bitb_76_60 bitb_76_61 R_bl
Cb_76_60 bit_76_60 gnd C_bl
Cbb_76_60 bitb_76_60 gnd C_bl
Rb_76_61 bit_76_61 bit_76_62 R_bl
Rbb_76_61 bitb_76_61 bitb_76_62 R_bl
Cb_76_61 bit_76_61 gnd C_bl
Cbb_76_61 bitb_76_61 gnd C_bl
Rb_76_62 bit_76_62 bit_76_63 R_bl
Rbb_76_62 bitb_76_62 bitb_76_63 R_bl
Cb_76_62 bit_76_62 gnd C_bl
Cbb_76_62 bitb_76_62 gnd C_bl
Rb_76_63 bit_76_63 bit_76_64 R_bl
Rbb_76_63 bitb_76_63 bitb_76_64 R_bl
Cb_76_63 bit_76_63 gnd C_bl
Cbb_76_63 bitb_76_63 gnd C_bl
Rb_76_64 bit_76_64 bit_76_65 R_bl
Rbb_76_64 bitb_76_64 bitb_76_65 R_bl
Cb_76_64 bit_76_64 gnd C_bl
Cbb_76_64 bitb_76_64 gnd C_bl
Rb_76_65 bit_76_65 bit_76_66 R_bl
Rbb_76_65 bitb_76_65 bitb_76_66 R_bl
Cb_76_65 bit_76_65 gnd C_bl
Cbb_76_65 bitb_76_65 gnd C_bl
Rb_76_66 bit_76_66 bit_76_67 R_bl
Rbb_76_66 bitb_76_66 bitb_76_67 R_bl
Cb_76_66 bit_76_66 gnd C_bl
Cbb_76_66 bitb_76_66 gnd C_bl
Rb_76_67 bit_76_67 bit_76_68 R_bl
Rbb_76_67 bitb_76_67 bitb_76_68 R_bl
Cb_76_67 bit_76_67 gnd C_bl
Cbb_76_67 bitb_76_67 gnd C_bl
Rb_76_68 bit_76_68 bit_76_69 R_bl
Rbb_76_68 bitb_76_68 bitb_76_69 R_bl
Cb_76_68 bit_76_68 gnd C_bl
Cbb_76_68 bitb_76_68 gnd C_bl
Rb_76_69 bit_76_69 bit_76_70 R_bl
Rbb_76_69 bitb_76_69 bitb_76_70 R_bl
Cb_76_69 bit_76_69 gnd C_bl
Cbb_76_69 bitb_76_69 gnd C_bl
Rb_76_70 bit_76_70 bit_76_71 R_bl
Rbb_76_70 bitb_76_70 bitb_76_71 R_bl
Cb_76_70 bit_76_70 gnd C_bl
Cbb_76_70 bitb_76_70 gnd C_bl
Rb_76_71 bit_76_71 bit_76_72 R_bl
Rbb_76_71 bitb_76_71 bitb_76_72 R_bl
Cb_76_71 bit_76_71 gnd C_bl
Cbb_76_71 bitb_76_71 gnd C_bl
Rb_76_72 bit_76_72 bit_76_73 R_bl
Rbb_76_72 bitb_76_72 bitb_76_73 R_bl
Cb_76_72 bit_76_72 gnd C_bl
Cbb_76_72 bitb_76_72 gnd C_bl
Rb_76_73 bit_76_73 bit_76_74 R_bl
Rbb_76_73 bitb_76_73 bitb_76_74 R_bl
Cb_76_73 bit_76_73 gnd C_bl
Cbb_76_73 bitb_76_73 gnd C_bl
Rb_76_74 bit_76_74 bit_76_75 R_bl
Rbb_76_74 bitb_76_74 bitb_76_75 R_bl
Cb_76_74 bit_76_74 gnd C_bl
Cbb_76_74 bitb_76_74 gnd C_bl
Rb_76_75 bit_76_75 bit_76_76 R_bl
Rbb_76_75 bitb_76_75 bitb_76_76 R_bl
Cb_76_75 bit_76_75 gnd C_bl
Cbb_76_75 bitb_76_75 gnd C_bl
Rb_76_76 bit_76_76 bit_76_77 R_bl
Rbb_76_76 bitb_76_76 bitb_76_77 R_bl
Cb_76_76 bit_76_76 gnd C_bl
Cbb_76_76 bitb_76_76 gnd C_bl
Rb_76_77 bit_76_77 bit_76_78 R_bl
Rbb_76_77 bitb_76_77 bitb_76_78 R_bl
Cb_76_77 bit_76_77 gnd C_bl
Cbb_76_77 bitb_76_77 gnd C_bl
Rb_76_78 bit_76_78 bit_76_79 R_bl
Rbb_76_78 bitb_76_78 bitb_76_79 R_bl
Cb_76_78 bit_76_78 gnd C_bl
Cbb_76_78 bitb_76_78 gnd C_bl
Rb_76_79 bit_76_79 bit_76_80 R_bl
Rbb_76_79 bitb_76_79 bitb_76_80 R_bl
Cb_76_79 bit_76_79 gnd C_bl
Cbb_76_79 bitb_76_79 gnd C_bl
Rb_76_80 bit_76_80 bit_76_81 R_bl
Rbb_76_80 bitb_76_80 bitb_76_81 R_bl
Cb_76_80 bit_76_80 gnd C_bl
Cbb_76_80 bitb_76_80 gnd C_bl
Rb_76_81 bit_76_81 bit_76_82 R_bl
Rbb_76_81 bitb_76_81 bitb_76_82 R_bl
Cb_76_81 bit_76_81 gnd C_bl
Cbb_76_81 bitb_76_81 gnd C_bl
Rb_76_82 bit_76_82 bit_76_83 R_bl
Rbb_76_82 bitb_76_82 bitb_76_83 R_bl
Cb_76_82 bit_76_82 gnd C_bl
Cbb_76_82 bitb_76_82 gnd C_bl
Rb_76_83 bit_76_83 bit_76_84 R_bl
Rbb_76_83 bitb_76_83 bitb_76_84 R_bl
Cb_76_83 bit_76_83 gnd C_bl
Cbb_76_83 bitb_76_83 gnd C_bl
Rb_76_84 bit_76_84 bit_76_85 R_bl
Rbb_76_84 bitb_76_84 bitb_76_85 R_bl
Cb_76_84 bit_76_84 gnd C_bl
Cbb_76_84 bitb_76_84 gnd C_bl
Rb_76_85 bit_76_85 bit_76_86 R_bl
Rbb_76_85 bitb_76_85 bitb_76_86 R_bl
Cb_76_85 bit_76_85 gnd C_bl
Cbb_76_85 bitb_76_85 gnd C_bl
Rb_76_86 bit_76_86 bit_76_87 R_bl
Rbb_76_86 bitb_76_86 bitb_76_87 R_bl
Cb_76_86 bit_76_86 gnd C_bl
Cbb_76_86 bitb_76_86 gnd C_bl
Rb_76_87 bit_76_87 bit_76_88 R_bl
Rbb_76_87 bitb_76_87 bitb_76_88 R_bl
Cb_76_87 bit_76_87 gnd C_bl
Cbb_76_87 bitb_76_87 gnd C_bl
Rb_76_88 bit_76_88 bit_76_89 R_bl
Rbb_76_88 bitb_76_88 bitb_76_89 R_bl
Cb_76_88 bit_76_88 gnd C_bl
Cbb_76_88 bitb_76_88 gnd C_bl
Rb_76_89 bit_76_89 bit_76_90 R_bl
Rbb_76_89 bitb_76_89 bitb_76_90 R_bl
Cb_76_89 bit_76_89 gnd C_bl
Cbb_76_89 bitb_76_89 gnd C_bl
Rb_76_90 bit_76_90 bit_76_91 R_bl
Rbb_76_90 bitb_76_90 bitb_76_91 R_bl
Cb_76_90 bit_76_90 gnd C_bl
Cbb_76_90 bitb_76_90 gnd C_bl
Rb_76_91 bit_76_91 bit_76_92 R_bl
Rbb_76_91 bitb_76_91 bitb_76_92 R_bl
Cb_76_91 bit_76_91 gnd C_bl
Cbb_76_91 bitb_76_91 gnd C_bl
Rb_76_92 bit_76_92 bit_76_93 R_bl
Rbb_76_92 bitb_76_92 bitb_76_93 R_bl
Cb_76_92 bit_76_92 gnd C_bl
Cbb_76_92 bitb_76_92 gnd C_bl
Rb_76_93 bit_76_93 bit_76_94 R_bl
Rbb_76_93 bitb_76_93 bitb_76_94 R_bl
Cb_76_93 bit_76_93 gnd C_bl
Cbb_76_93 bitb_76_93 gnd C_bl
Rb_76_94 bit_76_94 bit_76_95 R_bl
Rbb_76_94 bitb_76_94 bitb_76_95 R_bl
Cb_76_94 bit_76_94 gnd C_bl
Cbb_76_94 bitb_76_94 gnd C_bl
Rb_76_95 bit_76_95 bit_76_96 R_bl
Rbb_76_95 bitb_76_95 bitb_76_96 R_bl
Cb_76_95 bit_76_95 gnd C_bl
Cbb_76_95 bitb_76_95 gnd C_bl
Rb_76_96 bit_76_96 bit_76_97 R_bl
Rbb_76_96 bitb_76_96 bitb_76_97 R_bl
Cb_76_96 bit_76_96 gnd C_bl
Cbb_76_96 bitb_76_96 gnd C_bl
Rb_76_97 bit_76_97 bit_76_98 R_bl
Rbb_76_97 bitb_76_97 bitb_76_98 R_bl
Cb_76_97 bit_76_97 gnd C_bl
Cbb_76_97 bitb_76_97 gnd C_bl
Rb_76_98 bit_76_98 bit_76_99 R_bl
Rbb_76_98 bitb_76_98 bitb_76_99 R_bl
Cb_76_98 bit_76_98 gnd C_bl
Cbb_76_98 bitb_76_98 gnd C_bl
Rb_76_99 bit_76_99 bit_76_100 R_bl
Rbb_76_99 bitb_76_99 bitb_76_100 R_bl
Cb_76_99 bit_76_99 gnd C_bl
Cbb_76_99 bitb_76_99 gnd C_bl
Rb_77_0 bit_77_0 bit_77_1 R_bl
Rbb_77_0 bitb_77_0 bitb_77_1 R_bl
Cb_77_0 bit_77_0 gnd C_bl
Cbb_77_0 bitb_77_0 gnd C_bl
Rb_77_1 bit_77_1 bit_77_2 R_bl
Rbb_77_1 bitb_77_1 bitb_77_2 R_bl
Cb_77_1 bit_77_1 gnd C_bl
Cbb_77_1 bitb_77_1 gnd C_bl
Rb_77_2 bit_77_2 bit_77_3 R_bl
Rbb_77_2 bitb_77_2 bitb_77_3 R_bl
Cb_77_2 bit_77_2 gnd C_bl
Cbb_77_2 bitb_77_2 gnd C_bl
Rb_77_3 bit_77_3 bit_77_4 R_bl
Rbb_77_3 bitb_77_3 bitb_77_4 R_bl
Cb_77_3 bit_77_3 gnd C_bl
Cbb_77_3 bitb_77_3 gnd C_bl
Rb_77_4 bit_77_4 bit_77_5 R_bl
Rbb_77_4 bitb_77_4 bitb_77_5 R_bl
Cb_77_4 bit_77_4 gnd C_bl
Cbb_77_4 bitb_77_4 gnd C_bl
Rb_77_5 bit_77_5 bit_77_6 R_bl
Rbb_77_5 bitb_77_5 bitb_77_6 R_bl
Cb_77_5 bit_77_5 gnd C_bl
Cbb_77_5 bitb_77_5 gnd C_bl
Rb_77_6 bit_77_6 bit_77_7 R_bl
Rbb_77_6 bitb_77_6 bitb_77_7 R_bl
Cb_77_6 bit_77_6 gnd C_bl
Cbb_77_6 bitb_77_6 gnd C_bl
Rb_77_7 bit_77_7 bit_77_8 R_bl
Rbb_77_7 bitb_77_7 bitb_77_8 R_bl
Cb_77_7 bit_77_7 gnd C_bl
Cbb_77_7 bitb_77_7 gnd C_bl
Rb_77_8 bit_77_8 bit_77_9 R_bl
Rbb_77_8 bitb_77_8 bitb_77_9 R_bl
Cb_77_8 bit_77_8 gnd C_bl
Cbb_77_8 bitb_77_8 gnd C_bl
Rb_77_9 bit_77_9 bit_77_10 R_bl
Rbb_77_9 bitb_77_9 bitb_77_10 R_bl
Cb_77_9 bit_77_9 gnd C_bl
Cbb_77_9 bitb_77_9 gnd C_bl
Rb_77_10 bit_77_10 bit_77_11 R_bl
Rbb_77_10 bitb_77_10 bitb_77_11 R_bl
Cb_77_10 bit_77_10 gnd C_bl
Cbb_77_10 bitb_77_10 gnd C_bl
Rb_77_11 bit_77_11 bit_77_12 R_bl
Rbb_77_11 bitb_77_11 bitb_77_12 R_bl
Cb_77_11 bit_77_11 gnd C_bl
Cbb_77_11 bitb_77_11 gnd C_bl
Rb_77_12 bit_77_12 bit_77_13 R_bl
Rbb_77_12 bitb_77_12 bitb_77_13 R_bl
Cb_77_12 bit_77_12 gnd C_bl
Cbb_77_12 bitb_77_12 gnd C_bl
Rb_77_13 bit_77_13 bit_77_14 R_bl
Rbb_77_13 bitb_77_13 bitb_77_14 R_bl
Cb_77_13 bit_77_13 gnd C_bl
Cbb_77_13 bitb_77_13 gnd C_bl
Rb_77_14 bit_77_14 bit_77_15 R_bl
Rbb_77_14 bitb_77_14 bitb_77_15 R_bl
Cb_77_14 bit_77_14 gnd C_bl
Cbb_77_14 bitb_77_14 gnd C_bl
Rb_77_15 bit_77_15 bit_77_16 R_bl
Rbb_77_15 bitb_77_15 bitb_77_16 R_bl
Cb_77_15 bit_77_15 gnd C_bl
Cbb_77_15 bitb_77_15 gnd C_bl
Rb_77_16 bit_77_16 bit_77_17 R_bl
Rbb_77_16 bitb_77_16 bitb_77_17 R_bl
Cb_77_16 bit_77_16 gnd C_bl
Cbb_77_16 bitb_77_16 gnd C_bl
Rb_77_17 bit_77_17 bit_77_18 R_bl
Rbb_77_17 bitb_77_17 bitb_77_18 R_bl
Cb_77_17 bit_77_17 gnd C_bl
Cbb_77_17 bitb_77_17 gnd C_bl
Rb_77_18 bit_77_18 bit_77_19 R_bl
Rbb_77_18 bitb_77_18 bitb_77_19 R_bl
Cb_77_18 bit_77_18 gnd C_bl
Cbb_77_18 bitb_77_18 gnd C_bl
Rb_77_19 bit_77_19 bit_77_20 R_bl
Rbb_77_19 bitb_77_19 bitb_77_20 R_bl
Cb_77_19 bit_77_19 gnd C_bl
Cbb_77_19 bitb_77_19 gnd C_bl
Rb_77_20 bit_77_20 bit_77_21 R_bl
Rbb_77_20 bitb_77_20 bitb_77_21 R_bl
Cb_77_20 bit_77_20 gnd C_bl
Cbb_77_20 bitb_77_20 gnd C_bl
Rb_77_21 bit_77_21 bit_77_22 R_bl
Rbb_77_21 bitb_77_21 bitb_77_22 R_bl
Cb_77_21 bit_77_21 gnd C_bl
Cbb_77_21 bitb_77_21 gnd C_bl
Rb_77_22 bit_77_22 bit_77_23 R_bl
Rbb_77_22 bitb_77_22 bitb_77_23 R_bl
Cb_77_22 bit_77_22 gnd C_bl
Cbb_77_22 bitb_77_22 gnd C_bl
Rb_77_23 bit_77_23 bit_77_24 R_bl
Rbb_77_23 bitb_77_23 bitb_77_24 R_bl
Cb_77_23 bit_77_23 gnd C_bl
Cbb_77_23 bitb_77_23 gnd C_bl
Rb_77_24 bit_77_24 bit_77_25 R_bl
Rbb_77_24 bitb_77_24 bitb_77_25 R_bl
Cb_77_24 bit_77_24 gnd C_bl
Cbb_77_24 bitb_77_24 gnd C_bl
Rb_77_25 bit_77_25 bit_77_26 R_bl
Rbb_77_25 bitb_77_25 bitb_77_26 R_bl
Cb_77_25 bit_77_25 gnd C_bl
Cbb_77_25 bitb_77_25 gnd C_bl
Rb_77_26 bit_77_26 bit_77_27 R_bl
Rbb_77_26 bitb_77_26 bitb_77_27 R_bl
Cb_77_26 bit_77_26 gnd C_bl
Cbb_77_26 bitb_77_26 gnd C_bl
Rb_77_27 bit_77_27 bit_77_28 R_bl
Rbb_77_27 bitb_77_27 bitb_77_28 R_bl
Cb_77_27 bit_77_27 gnd C_bl
Cbb_77_27 bitb_77_27 gnd C_bl
Rb_77_28 bit_77_28 bit_77_29 R_bl
Rbb_77_28 bitb_77_28 bitb_77_29 R_bl
Cb_77_28 bit_77_28 gnd C_bl
Cbb_77_28 bitb_77_28 gnd C_bl
Rb_77_29 bit_77_29 bit_77_30 R_bl
Rbb_77_29 bitb_77_29 bitb_77_30 R_bl
Cb_77_29 bit_77_29 gnd C_bl
Cbb_77_29 bitb_77_29 gnd C_bl
Rb_77_30 bit_77_30 bit_77_31 R_bl
Rbb_77_30 bitb_77_30 bitb_77_31 R_bl
Cb_77_30 bit_77_30 gnd C_bl
Cbb_77_30 bitb_77_30 gnd C_bl
Rb_77_31 bit_77_31 bit_77_32 R_bl
Rbb_77_31 bitb_77_31 bitb_77_32 R_bl
Cb_77_31 bit_77_31 gnd C_bl
Cbb_77_31 bitb_77_31 gnd C_bl
Rb_77_32 bit_77_32 bit_77_33 R_bl
Rbb_77_32 bitb_77_32 bitb_77_33 R_bl
Cb_77_32 bit_77_32 gnd C_bl
Cbb_77_32 bitb_77_32 gnd C_bl
Rb_77_33 bit_77_33 bit_77_34 R_bl
Rbb_77_33 bitb_77_33 bitb_77_34 R_bl
Cb_77_33 bit_77_33 gnd C_bl
Cbb_77_33 bitb_77_33 gnd C_bl
Rb_77_34 bit_77_34 bit_77_35 R_bl
Rbb_77_34 bitb_77_34 bitb_77_35 R_bl
Cb_77_34 bit_77_34 gnd C_bl
Cbb_77_34 bitb_77_34 gnd C_bl
Rb_77_35 bit_77_35 bit_77_36 R_bl
Rbb_77_35 bitb_77_35 bitb_77_36 R_bl
Cb_77_35 bit_77_35 gnd C_bl
Cbb_77_35 bitb_77_35 gnd C_bl
Rb_77_36 bit_77_36 bit_77_37 R_bl
Rbb_77_36 bitb_77_36 bitb_77_37 R_bl
Cb_77_36 bit_77_36 gnd C_bl
Cbb_77_36 bitb_77_36 gnd C_bl
Rb_77_37 bit_77_37 bit_77_38 R_bl
Rbb_77_37 bitb_77_37 bitb_77_38 R_bl
Cb_77_37 bit_77_37 gnd C_bl
Cbb_77_37 bitb_77_37 gnd C_bl
Rb_77_38 bit_77_38 bit_77_39 R_bl
Rbb_77_38 bitb_77_38 bitb_77_39 R_bl
Cb_77_38 bit_77_38 gnd C_bl
Cbb_77_38 bitb_77_38 gnd C_bl
Rb_77_39 bit_77_39 bit_77_40 R_bl
Rbb_77_39 bitb_77_39 bitb_77_40 R_bl
Cb_77_39 bit_77_39 gnd C_bl
Cbb_77_39 bitb_77_39 gnd C_bl
Rb_77_40 bit_77_40 bit_77_41 R_bl
Rbb_77_40 bitb_77_40 bitb_77_41 R_bl
Cb_77_40 bit_77_40 gnd C_bl
Cbb_77_40 bitb_77_40 gnd C_bl
Rb_77_41 bit_77_41 bit_77_42 R_bl
Rbb_77_41 bitb_77_41 bitb_77_42 R_bl
Cb_77_41 bit_77_41 gnd C_bl
Cbb_77_41 bitb_77_41 gnd C_bl
Rb_77_42 bit_77_42 bit_77_43 R_bl
Rbb_77_42 bitb_77_42 bitb_77_43 R_bl
Cb_77_42 bit_77_42 gnd C_bl
Cbb_77_42 bitb_77_42 gnd C_bl
Rb_77_43 bit_77_43 bit_77_44 R_bl
Rbb_77_43 bitb_77_43 bitb_77_44 R_bl
Cb_77_43 bit_77_43 gnd C_bl
Cbb_77_43 bitb_77_43 gnd C_bl
Rb_77_44 bit_77_44 bit_77_45 R_bl
Rbb_77_44 bitb_77_44 bitb_77_45 R_bl
Cb_77_44 bit_77_44 gnd C_bl
Cbb_77_44 bitb_77_44 gnd C_bl
Rb_77_45 bit_77_45 bit_77_46 R_bl
Rbb_77_45 bitb_77_45 bitb_77_46 R_bl
Cb_77_45 bit_77_45 gnd C_bl
Cbb_77_45 bitb_77_45 gnd C_bl
Rb_77_46 bit_77_46 bit_77_47 R_bl
Rbb_77_46 bitb_77_46 bitb_77_47 R_bl
Cb_77_46 bit_77_46 gnd C_bl
Cbb_77_46 bitb_77_46 gnd C_bl
Rb_77_47 bit_77_47 bit_77_48 R_bl
Rbb_77_47 bitb_77_47 bitb_77_48 R_bl
Cb_77_47 bit_77_47 gnd C_bl
Cbb_77_47 bitb_77_47 gnd C_bl
Rb_77_48 bit_77_48 bit_77_49 R_bl
Rbb_77_48 bitb_77_48 bitb_77_49 R_bl
Cb_77_48 bit_77_48 gnd C_bl
Cbb_77_48 bitb_77_48 gnd C_bl
Rb_77_49 bit_77_49 bit_77_50 R_bl
Rbb_77_49 bitb_77_49 bitb_77_50 R_bl
Cb_77_49 bit_77_49 gnd C_bl
Cbb_77_49 bitb_77_49 gnd C_bl
Rb_77_50 bit_77_50 bit_77_51 R_bl
Rbb_77_50 bitb_77_50 bitb_77_51 R_bl
Cb_77_50 bit_77_50 gnd C_bl
Cbb_77_50 bitb_77_50 gnd C_bl
Rb_77_51 bit_77_51 bit_77_52 R_bl
Rbb_77_51 bitb_77_51 bitb_77_52 R_bl
Cb_77_51 bit_77_51 gnd C_bl
Cbb_77_51 bitb_77_51 gnd C_bl
Rb_77_52 bit_77_52 bit_77_53 R_bl
Rbb_77_52 bitb_77_52 bitb_77_53 R_bl
Cb_77_52 bit_77_52 gnd C_bl
Cbb_77_52 bitb_77_52 gnd C_bl
Rb_77_53 bit_77_53 bit_77_54 R_bl
Rbb_77_53 bitb_77_53 bitb_77_54 R_bl
Cb_77_53 bit_77_53 gnd C_bl
Cbb_77_53 bitb_77_53 gnd C_bl
Rb_77_54 bit_77_54 bit_77_55 R_bl
Rbb_77_54 bitb_77_54 bitb_77_55 R_bl
Cb_77_54 bit_77_54 gnd C_bl
Cbb_77_54 bitb_77_54 gnd C_bl
Rb_77_55 bit_77_55 bit_77_56 R_bl
Rbb_77_55 bitb_77_55 bitb_77_56 R_bl
Cb_77_55 bit_77_55 gnd C_bl
Cbb_77_55 bitb_77_55 gnd C_bl
Rb_77_56 bit_77_56 bit_77_57 R_bl
Rbb_77_56 bitb_77_56 bitb_77_57 R_bl
Cb_77_56 bit_77_56 gnd C_bl
Cbb_77_56 bitb_77_56 gnd C_bl
Rb_77_57 bit_77_57 bit_77_58 R_bl
Rbb_77_57 bitb_77_57 bitb_77_58 R_bl
Cb_77_57 bit_77_57 gnd C_bl
Cbb_77_57 bitb_77_57 gnd C_bl
Rb_77_58 bit_77_58 bit_77_59 R_bl
Rbb_77_58 bitb_77_58 bitb_77_59 R_bl
Cb_77_58 bit_77_58 gnd C_bl
Cbb_77_58 bitb_77_58 gnd C_bl
Rb_77_59 bit_77_59 bit_77_60 R_bl
Rbb_77_59 bitb_77_59 bitb_77_60 R_bl
Cb_77_59 bit_77_59 gnd C_bl
Cbb_77_59 bitb_77_59 gnd C_bl
Rb_77_60 bit_77_60 bit_77_61 R_bl
Rbb_77_60 bitb_77_60 bitb_77_61 R_bl
Cb_77_60 bit_77_60 gnd C_bl
Cbb_77_60 bitb_77_60 gnd C_bl
Rb_77_61 bit_77_61 bit_77_62 R_bl
Rbb_77_61 bitb_77_61 bitb_77_62 R_bl
Cb_77_61 bit_77_61 gnd C_bl
Cbb_77_61 bitb_77_61 gnd C_bl
Rb_77_62 bit_77_62 bit_77_63 R_bl
Rbb_77_62 bitb_77_62 bitb_77_63 R_bl
Cb_77_62 bit_77_62 gnd C_bl
Cbb_77_62 bitb_77_62 gnd C_bl
Rb_77_63 bit_77_63 bit_77_64 R_bl
Rbb_77_63 bitb_77_63 bitb_77_64 R_bl
Cb_77_63 bit_77_63 gnd C_bl
Cbb_77_63 bitb_77_63 gnd C_bl
Rb_77_64 bit_77_64 bit_77_65 R_bl
Rbb_77_64 bitb_77_64 bitb_77_65 R_bl
Cb_77_64 bit_77_64 gnd C_bl
Cbb_77_64 bitb_77_64 gnd C_bl
Rb_77_65 bit_77_65 bit_77_66 R_bl
Rbb_77_65 bitb_77_65 bitb_77_66 R_bl
Cb_77_65 bit_77_65 gnd C_bl
Cbb_77_65 bitb_77_65 gnd C_bl
Rb_77_66 bit_77_66 bit_77_67 R_bl
Rbb_77_66 bitb_77_66 bitb_77_67 R_bl
Cb_77_66 bit_77_66 gnd C_bl
Cbb_77_66 bitb_77_66 gnd C_bl
Rb_77_67 bit_77_67 bit_77_68 R_bl
Rbb_77_67 bitb_77_67 bitb_77_68 R_bl
Cb_77_67 bit_77_67 gnd C_bl
Cbb_77_67 bitb_77_67 gnd C_bl
Rb_77_68 bit_77_68 bit_77_69 R_bl
Rbb_77_68 bitb_77_68 bitb_77_69 R_bl
Cb_77_68 bit_77_68 gnd C_bl
Cbb_77_68 bitb_77_68 gnd C_bl
Rb_77_69 bit_77_69 bit_77_70 R_bl
Rbb_77_69 bitb_77_69 bitb_77_70 R_bl
Cb_77_69 bit_77_69 gnd C_bl
Cbb_77_69 bitb_77_69 gnd C_bl
Rb_77_70 bit_77_70 bit_77_71 R_bl
Rbb_77_70 bitb_77_70 bitb_77_71 R_bl
Cb_77_70 bit_77_70 gnd C_bl
Cbb_77_70 bitb_77_70 gnd C_bl
Rb_77_71 bit_77_71 bit_77_72 R_bl
Rbb_77_71 bitb_77_71 bitb_77_72 R_bl
Cb_77_71 bit_77_71 gnd C_bl
Cbb_77_71 bitb_77_71 gnd C_bl
Rb_77_72 bit_77_72 bit_77_73 R_bl
Rbb_77_72 bitb_77_72 bitb_77_73 R_bl
Cb_77_72 bit_77_72 gnd C_bl
Cbb_77_72 bitb_77_72 gnd C_bl
Rb_77_73 bit_77_73 bit_77_74 R_bl
Rbb_77_73 bitb_77_73 bitb_77_74 R_bl
Cb_77_73 bit_77_73 gnd C_bl
Cbb_77_73 bitb_77_73 gnd C_bl
Rb_77_74 bit_77_74 bit_77_75 R_bl
Rbb_77_74 bitb_77_74 bitb_77_75 R_bl
Cb_77_74 bit_77_74 gnd C_bl
Cbb_77_74 bitb_77_74 gnd C_bl
Rb_77_75 bit_77_75 bit_77_76 R_bl
Rbb_77_75 bitb_77_75 bitb_77_76 R_bl
Cb_77_75 bit_77_75 gnd C_bl
Cbb_77_75 bitb_77_75 gnd C_bl
Rb_77_76 bit_77_76 bit_77_77 R_bl
Rbb_77_76 bitb_77_76 bitb_77_77 R_bl
Cb_77_76 bit_77_76 gnd C_bl
Cbb_77_76 bitb_77_76 gnd C_bl
Rb_77_77 bit_77_77 bit_77_78 R_bl
Rbb_77_77 bitb_77_77 bitb_77_78 R_bl
Cb_77_77 bit_77_77 gnd C_bl
Cbb_77_77 bitb_77_77 gnd C_bl
Rb_77_78 bit_77_78 bit_77_79 R_bl
Rbb_77_78 bitb_77_78 bitb_77_79 R_bl
Cb_77_78 bit_77_78 gnd C_bl
Cbb_77_78 bitb_77_78 gnd C_bl
Rb_77_79 bit_77_79 bit_77_80 R_bl
Rbb_77_79 bitb_77_79 bitb_77_80 R_bl
Cb_77_79 bit_77_79 gnd C_bl
Cbb_77_79 bitb_77_79 gnd C_bl
Rb_77_80 bit_77_80 bit_77_81 R_bl
Rbb_77_80 bitb_77_80 bitb_77_81 R_bl
Cb_77_80 bit_77_80 gnd C_bl
Cbb_77_80 bitb_77_80 gnd C_bl
Rb_77_81 bit_77_81 bit_77_82 R_bl
Rbb_77_81 bitb_77_81 bitb_77_82 R_bl
Cb_77_81 bit_77_81 gnd C_bl
Cbb_77_81 bitb_77_81 gnd C_bl
Rb_77_82 bit_77_82 bit_77_83 R_bl
Rbb_77_82 bitb_77_82 bitb_77_83 R_bl
Cb_77_82 bit_77_82 gnd C_bl
Cbb_77_82 bitb_77_82 gnd C_bl
Rb_77_83 bit_77_83 bit_77_84 R_bl
Rbb_77_83 bitb_77_83 bitb_77_84 R_bl
Cb_77_83 bit_77_83 gnd C_bl
Cbb_77_83 bitb_77_83 gnd C_bl
Rb_77_84 bit_77_84 bit_77_85 R_bl
Rbb_77_84 bitb_77_84 bitb_77_85 R_bl
Cb_77_84 bit_77_84 gnd C_bl
Cbb_77_84 bitb_77_84 gnd C_bl
Rb_77_85 bit_77_85 bit_77_86 R_bl
Rbb_77_85 bitb_77_85 bitb_77_86 R_bl
Cb_77_85 bit_77_85 gnd C_bl
Cbb_77_85 bitb_77_85 gnd C_bl
Rb_77_86 bit_77_86 bit_77_87 R_bl
Rbb_77_86 bitb_77_86 bitb_77_87 R_bl
Cb_77_86 bit_77_86 gnd C_bl
Cbb_77_86 bitb_77_86 gnd C_bl
Rb_77_87 bit_77_87 bit_77_88 R_bl
Rbb_77_87 bitb_77_87 bitb_77_88 R_bl
Cb_77_87 bit_77_87 gnd C_bl
Cbb_77_87 bitb_77_87 gnd C_bl
Rb_77_88 bit_77_88 bit_77_89 R_bl
Rbb_77_88 bitb_77_88 bitb_77_89 R_bl
Cb_77_88 bit_77_88 gnd C_bl
Cbb_77_88 bitb_77_88 gnd C_bl
Rb_77_89 bit_77_89 bit_77_90 R_bl
Rbb_77_89 bitb_77_89 bitb_77_90 R_bl
Cb_77_89 bit_77_89 gnd C_bl
Cbb_77_89 bitb_77_89 gnd C_bl
Rb_77_90 bit_77_90 bit_77_91 R_bl
Rbb_77_90 bitb_77_90 bitb_77_91 R_bl
Cb_77_90 bit_77_90 gnd C_bl
Cbb_77_90 bitb_77_90 gnd C_bl
Rb_77_91 bit_77_91 bit_77_92 R_bl
Rbb_77_91 bitb_77_91 bitb_77_92 R_bl
Cb_77_91 bit_77_91 gnd C_bl
Cbb_77_91 bitb_77_91 gnd C_bl
Rb_77_92 bit_77_92 bit_77_93 R_bl
Rbb_77_92 bitb_77_92 bitb_77_93 R_bl
Cb_77_92 bit_77_92 gnd C_bl
Cbb_77_92 bitb_77_92 gnd C_bl
Rb_77_93 bit_77_93 bit_77_94 R_bl
Rbb_77_93 bitb_77_93 bitb_77_94 R_bl
Cb_77_93 bit_77_93 gnd C_bl
Cbb_77_93 bitb_77_93 gnd C_bl
Rb_77_94 bit_77_94 bit_77_95 R_bl
Rbb_77_94 bitb_77_94 bitb_77_95 R_bl
Cb_77_94 bit_77_94 gnd C_bl
Cbb_77_94 bitb_77_94 gnd C_bl
Rb_77_95 bit_77_95 bit_77_96 R_bl
Rbb_77_95 bitb_77_95 bitb_77_96 R_bl
Cb_77_95 bit_77_95 gnd C_bl
Cbb_77_95 bitb_77_95 gnd C_bl
Rb_77_96 bit_77_96 bit_77_97 R_bl
Rbb_77_96 bitb_77_96 bitb_77_97 R_bl
Cb_77_96 bit_77_96 gnd C_bl
Cbb_77_96 bitb_77_96 gnd C_bl
Rb_77_97 bit_77_97 bit_77_98 R_bl
Rbb_77_97 bitb_77_97 bitb_77_98 R_bl
Cb_77_97 bit_77_97 gnd C_bl
Cbb_77_97 bitb_77_97 gnd C_bl
Rb_77_98 bit_77_98 bit_77_99 R_bl
Rbb_77_98 bitb_77_98 bitb_77_99 R_bl
Cb_77_98 bit_77_98 gnd C_bl
Cbb_77_98 bitb_77_98 gnd C_bl
Rb_77_99 bit_77_99 bit_77_100 R_bl
Rbb_77_99 bitb_77_99 bitb_77_100 R_bl
Cb_77_99 bit_77_99 gnd C_bl
Cbb_77_99 bitb_77_99 gnd C_bl
Rb_78_0 bit_78_0 bit_78_1 R_bl
Rbb_78_0 bitb_78_0 bitb_78_1 R_bl
Cb_78_0 bit_78_0 gnd C_bl
Cbb_78_0 bitb_78_0 gnd C_bl
Rb_78_1 bit_78_1 bit_78_2 R_bl
Rbb_78_1 bitb_78_1 bitb_78_2 R_bl
Cb_78_1 bit_78_1 gnd C_bl
Cbb_78_1 bitb_78_1 gnd C_bl
Rb_78_2 bit_78_2 bit_78_3 R_bl
Rbb_78_2 bitb_78_2 bitb_78_3 R_bl
Cb_78_2 bit_78_2 gnd C_bl
Cbb_78_2 bitb_78_2 gnd C_bl
Rb_78_3 bit_78_3 bit_78_4 R_bl
Rbb_78_3 bitb_78_3 bitb_78_4 R_bl
Cb_78_3 bit_78_3 gnd C_bl
Cbb_78_3 bitb_78_3 gnd C_bl
Rb_78_4 bit_78_4 bit_78_5 R_bl
Rbb_78_4 bitb_78_4 bitb_78_5 R_bl
Cb_78_4 bit_78_4 gnd C_bl
Cbb_78_4 bitb_78_4 gnd C_bl
Rb_78_5 bit_78_5 bit_78_6 R_bl
Rbb_78_5 bitb_78_5 bitb_78_6 R_bl
Cb_78_5 bit_78_5 gnd C_bl
Cbb_78_5 bitb_78_5 gnd C_bl
Rb_78_6 bit_78_6 bit_78_7 R_bl
Rbb_78_6 bitb_78_6 bitb_78_7 R_bl
Cb_78_6 bit_78_6 gnd C_bl
Cbb_78_6 bitb_78_6 gnd C_bl
Rb_78_7 bit_78_7 bit_78_8 R_bl
Rbb_78_7 bitb_78_7 bitb_78_8 R_bl
Cb_78_7 bit_78_7 gnd C_bl
Cbb_78_7 bitb_78_7 gnd C_bl
Rb_78_8 bit_78_8 bit_78_9 R_bl
Rbb_78_8 bitb_78_8 bitb_78_9 R_bl
Cb_78_8 bit_78_8 gnd C_bl
Cbb_78_8 bitb_78_8 gnd C_bl
Rb_78_9 bit_78_9 bit_78_10 R_bl
Rbb_78_9 bitb_78_9 bitb_78_10 R_bl
Cb_78_9 bit_78_9 gnd C_bl
Cbb_78_9 bitb_78_9 gnd C_bl
Rb_78_10 bit_78_10 bit_78_11 R_bl
Rbb_78_10 bitb_78_10 bitb_78_11 R_bl
Cb_78_10 bit_78_10 gnd C_bl
Cbb_78_10 bitb_78_10 gnd C_bl
Rb_78_11 bit_78_11 bit_78_12 R_bl
Rbb_78_11 bitb_78_11 bitb_78_12 R_bl
Cb_78_11 bit_78_11 gnd C_bl
Cbb_78_11 bitb_78_11 gnd C_bl
Rb_78_12 bit_78_12 bit_78_13 R_bl
Rbb_78_12 bitb_78_12 bitb_78_13 R_bl
Cb_78_12 bit_78_12 gnd C_bl
Cbb_78_12 bitb_78_12 gnd C_bl
Rb_78_13 bit_78_13 bit_78_14 R_bl
Rbb_78_13 bitb_78_13 bitb_78_14 R_bl
Cb_78_13 bit_78_13 gnd C_bl
Cbb_78_13 bitb_78_13 gnd C_bl
Rb_78_14 bit_78_14 bit_78_15 R_bl
Rbb_78_14 bitb_78_14 bitb_78_15 R_bl
Cb_78_14 bit_78_14 gnd C_bl
Cbb_78_14 bitb_78_14 gnd C_bl
Rb_78_15 bit_78_15 bit_78_16 R_bl
Rbb_78_15 bitb_78_15 bitb_78_16 R_bl
Cb_78_15 bit_78_15 gnd C_bl
Cbb_78_15 bitb_78_15 gnd C_bl
Rb_78_16 bit_78_16 bit_78_17 R_bl
Rbb_78_16 bitb_78_16 bitb_78_17 R_bl
Cb_78_16 bit_78_16 gnd C_bl
Cbb_78_16 bitb_78_16 gnd C_bl
Rb_78_17 bit_78_17 bit_78_18 R_bl
Rbb_78_17 bitb_78_17 bitb_78_18 R_bl
Cb_78_17 bit_78_17 gnd C_bl
Cbb_78_17 bitb_78_17 gnd C_bl
Rb_78_18 bit_78_18 bit_78_19 R_bl
Rbb_78_18 bitb_78_18 bitb_78_19 R_bl
Cb_78_18 bit_78_18 gnd C_bl
Cbb_78_18 bitb_78_18 gnd C_bl
Rb_78_19 bit_78_19 bit_78_20 R_bl
Rbb_78_19 bitb_78_19 bitb_78_20 R_bl
Cb_78_19 bit_78_19 gnd C_bl
Cbb_78_19 bitb_78_19 gnd C_bl
Rb_78_20 bit_78_20 bit_78_21 R_bl
Rbb_78_20 bitb_78_20 bitb_78_21 R_bl
Cb_78_20 bit_78_20 gnd C_bl
Cbb_78_20 bitb_78_20 gnd C_bl
Rb_78_21 bit_78_21 bit_78_22 R_bl
Rbb_78_21 bitb_78_21 bitb_78_22 R_bl
Cb_78_21 bit_78_21 gnd C_bl
Cbb_78_21 bitb_78_21 gnd C_bl
Rb_78_22 bit_78_22 bit_78_23 R_bl
Rbb_78_22 bitb_78_22 bitb_78_23 R_bl
Cb_78_22 bit_78_22 gnd C_bl
Cbb_78_22 bitb_78_22 gnd C_bl
Rb_78_23 bit_78_23 bit_78_24 R_bl
Rbb_78_23 bitb_78_23 bitb_78_24 R_bl
Cb_78_23 bit_78_23 gnd C_bl
Cbb_78_23 bitb_78_23 gnd C_bl
Rb_78_24 bit_78_24 bit_78_25 R_bl
Rbb_78_24 bitb_78_24 bitb_78_25 R_bl
Cb_78_24 bit_78_24 gnd C_bl
Cbb_78_24 bitb_78_24 gnd C_bl
Rb_78_25 bit_78_25 bit_78_26 R_bl
Rbb_78_25 bitb_78_25 bitb_78_26 R_bl
Cb_78_25 bit_78_25 gnd C_bl
Cbb_78_25 bitb_78_25 gnd C_bl
Rb_78_26 bit_78_26 bit_78_27 R_bl
Rbb_78_26 bitb_78_26 bitb_78_27 R_bl
Cb_78_26 bit_78_26 gnd C_bl
Cbb_78_26 bitb_78_26 gnd C_bl
Rb_78_27 bit_78_27 bit_78_28 R_bl
Rbb_78_27 bitb_78_27 bitb_78_28 R_bl
Cb_78_27 bit_78_27 gnd C_bl
Cbb_78_27 bitb_78_27 gnd C_bl
Rb_78_28 bit_78_28 bit_78_29 R_bl
Rbb_78_28 bitb_78_28 bitb_78_29 R_bl
Cb_78_28 bit_78_28 gnd C_bl
Cbb_78_28 bitb_78_28 gnd C_bl
Rb_78_29 bit_78_29 bit_78_30 R_bl
Rbb_78_29 bitb_78_29 bitb_78_30 R_bl
Cb_78_29 bit_78_29 gnd C_bl
Cbb_78_29 bitb_78_29 gnd C_bl
Rb_78_30 bit_78_30 bit_78_31 R_bl
Rbb_78_30 bitb_78_30 bitb_78_31 R_bl
Cb_78_30 bit_78_30 gnd C_bl
Cbb_78_30 bitb_78_30 gnd C_bl
Rb_78_31 bit_78_31 bit_78_32 R_bl
Rbb_78_31 bitb_78_31 bitb_78_32 R_bl
Cb_78_31 bit_78_31 gnd C_bl
Cbb_78_31 bitb_78_31 gnd C_bl
Rb_78_32 bit_78_32 bit_78_33 R_bl
Rbb_78_32 bitb_78_32 bitb_78_33 R_bl
Cb_78_32 bit_78_32 gnd C_bl
Cbb_78_32 bitb_78_32 gnd C_bl
Rb_78_33 bit_78_33 bit_78_34 R_bl
Rbb_78_33 bitb_78_33 bitb_78_34 R_bl
Cb_78_33 bit_78_33 gnd C_bl
Cbb_78_33 bitb_78_33 gnd C_bl
Rb_78_34 bit_78_34 bit_78_35 R_bl
Rbb_78_34 bitb_78_34 bitb_78_35 R_bl
Cb_78_34 bit_78_34 gnd C_bl
Cbb_78_34 bitb_78_34 gnd C_bl
Rb_78_35 bit_78_35 bit_78_36 R_bl
Rbb_78_35 bitb_78_35 bitb_78_36 R_bl
Cb_78_35 bit_78_35 gnd C_bl
Cbb_78_35 bitb_78_35 gnd C_bl
Rb_78_36 bit_78_36 bit_78_37 R_bl
Rbb_78_36 bitb_78_36 bitb_78_37 R_bl
Cb_78_36 bit_78_36 gnd C_bl
Cbb_78_36 bitb_78_36 gnd C_bl
Rb_78_37 bit_78_37 bit_78_38 R_bl
Rbb_78_37 bitb_78_37 bitb_78_38 R_bl
Cb_78_37 bit_78_37 gnd C_bl
Cbb_78_37 bitb_78_37 gnd C_bl
Rb_78_38 bit_78_38 bit_78_39 R_bl
Rbb_78_38 bitb_78_38 bitb_78_39 R_bl
Cb_78_38 bit_78_38 gnd C_bl
Cbb_78_38 bitb_78_38 gnd C_bl
Rb_78_39 bit_78_39 bit_78_40 R_bl
Rbb_78_39 bitb_78_39 bitb_78_40 R_bl
Cb_78_39 bit_78_39 gnd C_bl
Cbb_78_39 bitb_78_39 gnd C_bl
Rb_78_40 bit_78_40 bit_78_41 R_bl
Rbb_78_40 bitb_78_40 bitb_78_41 R_bl
Cb_78_40 bit_78_40 gnd C_bl
Cbb_78_40 bitb_78_40 gnd C_bl
Rb_78_41 bit_78_41 bit_78_42 R_bl
Rbb_78_41 bitb_78_41 bitb_78_42 R_bl
Cb_78_41 bit_78_41 gnd C_bl
Cbb_78_41 bitb_78_41 gnd C_bl
Rb_78_42 bit_78_42 bit_78_43 R_bl
Rbb_78_42 bitb_78_42 bitb_78_43 R_bl
Cb_78_42 bit_78_42 gnd C_bl
Cbb_78_42 bitb_78_42 gnd C_bl
Rb_78_43 bit_78_43 bit_78_44 R_bl
Rbb_78_43 bitb_78_43 bitb_78_44 R_bl
Cb_78_43 bit_78_43 gnd C_bl
Cbb_78_43 bitb_78_43 gnd C_bl
Rb_78_44 bit_78_44 bit_78_45 R_bl
Rbb_78_44 bitb_78_44 bitb_78_45 R_bl
Cb_78_44 bit_78_44 gnd C_bl
Cbb_78_44 bitb_78_44 gnd C_bl
Rb_78_45 bit_78_45 bit_78_46 R_bl
Rbb_78_45 bitb_78_45 bitb_78_46 R_bl
Cb_78_45 bit_78_45 gnd C_bl
Cbb_78_45 bitb_78_45 gnd C_bl
Rb_78_46 bit_78_46 bit_78_47 R_bl
Rbb_78_46 bitb_78_46 bitb_78_47 R_bl
Cb_78_46 bit_78_46 gnd C_bl
Cbb_78_46 bitb_78_46 gnd C_bl
Rb_78_47 bit_78_47 bit_78_48 R_bl
Rbb_78_47 bitb_78_47 bitb_78_48 R_bl
Cb_78_47 bit_78_47 gnd C_bl
Cbb_78_47 bitb_78_47 gnd C_bl
Rb_78_48 bit_78_48 bit_78_49 R_bl
Rbb_78_48 bitb_78_48 bitb_78_49 R_bl
Cb_78_48 bit_78_48 gnd C_bl
Cbb_78_48 bitb_78_48 gnd C_bl
Rb_78_49 bit_78_49 bit_78_50 R_bl
Rbb_78_49 bitb_78_49 bitb_78_50 R_bl
Cb_78_49 bit_78_49 gnd C_bl
Cbb_78_49 bitb_78_49 gnd C_bl
Rb_78_50 bit_78_50 bit_78_51 R_bl
Rbb_78_50 bitb_78_50 bitb_78_51 R_bl
Cb_78_50 bit_78_50 gnd C_bl
Cbb_78_50 bitb_78_50 gnd C_bl
Rb_78_51 bit_78_51 bit_78_52 R_bl
Rbb_78_51 bitb_78_51 bitb_78_52 R_bl
Cb_78_51 bit_78_51 gnd C_bl
Cbb_78_51 bitb_78_51 gnd C_bl
Rb_78_52 bit_78_52 bit_78_53 R_bl
Rbb_78_52 bitb_78_52 bitb_78_53 R_bl
Cb_78_52 bit_78_52 gnd C_bl
Cbb_78_52 bitb_78_52 gnd C_bl
Rb_78_53 bit_78_53 bit_78_54 R_bl
Rbb_78_53 bitb_78_53 bitb_78_54 R_bl
Cb_78_53 bit_78_53 gnd C_bl
Cbb_78_53 bitb_78_53 gnd C_bl
Rb_78_54 bit_78_54 bit_78_55 R_bl
Rbb_78_54 bitb_78_54 bitb_78_55 R_bl
Cb_78_54 bit_78_54 gnd C_bl
Cbb_78_54 bitb_78_54 gnd C_bl
Rb_78_55 bit_78_55 bit_78_56 R_bl
Rbb_78_55 bitb_78_55 bitb_78_56 R_bl
Cb_78_55 bit_78_55 gnd C_bl
Cbb_78_55 bitb_78_55 gnd C_bl
Rb_78_56 bit_78_56 bit_78_57 R_bl
Rbb_78_56 bitb_78_56 bitb_78_57 R_bl
Cb_78_56 bit_78_56 gnd C_bl
Cbb_78_56 bitb_78_56 gnd C_bl
Rb_78_57 bit_78_57 bit_78_58 R_bl
Rbb_78_57 bitb_78_57 bitb_78_58 R_bl
Cb_78_57 bit_78_57 gnd C_bl
Cbb_78_57 bitb_78_57 gnd C_bl
Rb_78_58 bit_78_58 bit_78_59 R_bl
Rbb_78_58 bitb_78_58 bitb_78_59 R_bl
Cb_78_58 bit_78_58 gnd C_bl
Cbb_78_58 bitb_78_58 gnd C_bl
Rb_78_59 bit_78_59 bit_78_60 R_bl
Rbb_78_59 bitb_78_59 bitb_78_60 R_bl
Cb_78_59 bit_78_59 gnd C_bl
Cbb_78_59 bitb_78_59 gnd C_bl
Rb_78_60 bit_78_60 bit_78_61 R_bl
Rbb_78_60 bitb_78_60 bitb_78_61 R_bl
Cb_78_60 bit_78_60 gnd C_bl
Cbb_78_60 bitb_78_60 gnd C_bl
Rb_78_61 bit_78_61 bit_78_62 R_bl
Rbb_78_61 bitb_78_61 bitb_78_62 R_bl
Cb_78_61 bit_78_61 gnd C_bl
Cbb_78_61 bitb_78_61 gnd C_bl
Rb_78_62 bit_78_62 bit_78_63 R_bl
Rbb_78_62 bitb_78_62 bitb_78_63 R_bl
Cb_78_62 bit_78_62 gnd C_bl
Cbb_78_62 bitb_78_62 gnd C_bl
Rb_78_63 bit_78_63 bit_78_64 R_bl
Rbb_78_63 bitb_78_63 bitb_78_64 R_bl
Cb_78_63 bit_78_63 gnd C_bl
Cbb_78_63 bitb_78_63 gnd C_bl
Rb_78_64 bit_78_64 bit_78_65 R_bl
Rbb_78_64 bitb_78_64 bitb_78_65 R_bl
Cb_78_64 bit_78_64 gnd C_bl
Cbb_78_64 bitb_78_64 gnd C_bl
Rb_78_65 bit_78_65 bit_78_66 R_bl
Rbb_78_65 bitb_78_65 bitb_78_66 R_bl
Cb_78_65 bit_78_65 gnd C_bl
Cbb_78_65 bitb_78_65 gnd C_bl
Rb_78_66 bit_78_66 bit_78_67 R_bl
Rbb_78_66 bitb_78_66 bitb_78_67 R_bl
Cb_78_66 bit_78_66 gnd C_bl
Cbb_78_66 bitb_78_66 gnd C_bl
Rb_78_67 bit_78_67 bit_78_68 R_bl
Rbb_78_67 bitb_78_67 bitb_78_68 R_bl
Cb_78_67 bit_78_67 gnd C_bl
Cbb_78_67 bitb_78_67 gnd C_bl
Rb_78_68 bit_78_68 bit_78_69 R_bl
Rbb_78_68 bitb_78_68 bitb_78_69 R_bl
Cb_78_68 bit_78_68 gnd C_bl
Cbb_78_68 bitb_78_68 gnd C_bl
Rb_78_69 bit_78_69 bit_78_70 R_bl
Rbb_78_69 bitb_78_69 bitb_78_70 R_bl
Cb_78_69 bit_78_69 gnd C_bl
Cbb_78_69 bitb_78_69 gnd C_bl
Rb_78_70 bit_78_70 bit_78_71 R_bl
Rbb_78_70 bitb_78_70 bitb_78_71 R_bl
Cb_78_70 bit_78_70 gnd C_bl
Cbb_78_70 bitb_78_70 gnd C_bl
Rb_78_71 bit_78_71 bit_78_72 R_bl
Rbb_78_71 bitb_78_71 bitb_78_72 R_bl
Cb_78_71 bit_78_71 gnd C_bl
Cbb_78_71 bitb_78_71 gnd C_bl
Rb_78_72 bit_78_72 bit_78_73 R_bl
Rbb_78_72 bitb_78_72 bitb_78_73 R_bl
Cb_78_72 bit_78_72 gnd C_bl
Cbb_78_72 bitb_78_72 gnd C_bl
Rb_78_73 bit_78_73 bit_78_74 R_bl
Rbb_78_73 bitb_78_73 bitb_78_74 R_bl
Cb_78_73 bit_78_73 gnd C_bl
Cbb_78_73 bitb_78_73 gnd C_bl
Rb_78_74 bit_78_74 bit_78_75 R_bl
Rbb_78_74 bitb_78_74 bitb_78_75 R_bl
Cb_78_74 bit_78_74 gnd C_bl
Cbb_78_74 bitb_78_74 gnd C_bl
Rb_78_75 bit_78_75 bit_78_76 R_bl
Rbb_78_75 bitb_78_75 bitb_78_76 R_bl
Cb_78_75 bit_78_75 gnd C_bl
Cbb_78_75 bitb_78_75 gnd C_bl
Rb_78_76 bit_78_76 bit_78_77 R_bl
Rbb_78_76 bitb_78_76 bitb_78_77 R_bl
Cb_78_76 bit_78_76 gnd C_bl
Cbb_78_76 bitb_78_76 gnd C_bl
Rb_78_77 bit_78_77 bit_78_78 R_bl
Rbb_78_77 bitb_78_77 bitb_78_78 R_bl
Cb_78_77 bit_78_77 gnd C_bl
Cbb_78_77 bitb_78_77 gnd C_bl
Rb_78_78 bit_78_78 bit_78_79 R_bl
Rbb_78_78 bitb_78_78 bitb_78_79 R_bl
Cb_78_78 bit_78_78 gnd C_bl
Cbb_78_78 bitb_78_78 gnd C_bl
Rb_78_79 bit_78_79 bit_78_80 R_bl
Rbb_78_79 bitb_78_79 bitb_78_80 R_bl
Cb_78_79 bit_78_79 gnd C_bl
Cbb_78_79 bitb_78_79 gnd C_bl
Rb_78_80 bit_78_80 bit_78_81 R_bl
Rbb_78_80 bitb_78_80 bitb_78_81 R_bl
Cb_78_80 bit_78_80 gnd C_bl
Cbb_78_80 bitb_78_80 gnd C_bl
Rb_78_81 bit_78_81 bit_78_82 R_bl
Rbb_78_81 bitb_78_81 bitb_78_82 R_bl
Cb_78_81 bit_78_81 gnd C_bl
Cbb_78_81 bitb_78_81 gnd C_bl
Rb_78_82 bit_78_82 bit_78_83 R_bl
Rbb_78_82 bitb_78_82 bitb_78_83 R_bl
Cb_78_82 bit_78_82 gnd C_bl
Cbb_78_82 bitb_78_82 gnd C_bl
Rb_78_83 bit_78_83 bit_78_84 R_bl
Rbb_78_83 bitb_78_83 bitb_78_84 R_bl
Cb_78_83 bit_78_83 gnd C_bl
Cbb_78_83 bitb_78_83 gnd C_bl
Rb_78_84 bit_78_84 bit_78_85 R_bl
Rbb_78_84 bitb_78_84 bitb_78_85 R_bl
Cb_78_84 bit_78_84 gnd C_bl
Cbb_78_84 bitb_78_84 gnd C_bl
Rb_78_85 bit_78_85 bit_78_86 R_bl
Rbb_78_85 bitb_78_85 bitb_78_86 R_bl
Cb_78_85 bit_78_85 gnd C_bl
Cbb_78_85 bitb_78_85 gnd C_bl
Rb_78_86 bit_78_86 bit_78_87 R_bl
Rbb_78_86 bitb_78_86 bitb_78_87 R_bl
Cb_78_86 bit_78_86 gnd C_bl
Cbb_78_86 bitb_78_86 gnd C_bl
Rb_78_87 bit_78_87 bit_78_88 R_bl
Rbb_78_87 bitb_78_87 bitb_78_88 R_bl
Cb_78_87 bit_78_87 gnd C_bl
Cbb_78_87 bitb_78_87 gnd C_bl
Rb_78_88 bit_78_88 bit_78_89 R_bl
Rbb_78_88 bitb_78_88 bitb_78_89 R_bl
Cb_78_88 bit_78_88 gnd C_bl
Cbb_78_88 bitb_78_88 gnd C_bl
Rb_78_89 bit_78_89 bit_78_90 R_bl
Rbb_78_89 bitb_78_89 bitb_78_90 R_bl
Cb_78_89 bit_78_89 gnd C_bl
Cbb_78_89 bitb_78_89 gnd C_bl
Rb_78_90 bit_78_90 bit_78_91 R_bl
Rbb_78_90 bitb_78_90 bitb_78_91 R_bl
Cb_78_90 bit_78_90 gnd C_bl
Cbb_78_90 bitb_78_90 gnd C_bl
Rb_78_91 bit_78_91 bit_78_92 R_bl
Rbb_78_91 bitb_78_91 bitb_78_92 R_bl
Cb_78_91 bit_78_91 gnd C_bl
Cbb_78_91 bitb_78_91 gnd C_bl
Rb_78_92 bit_78_92 bit_78_93 R_bl
Rbb_78_92 bitb_78_92 bitb_78_93 R_bl
Cb_78_92 bit_78_92 gnd C_bl
Cbb_78_92 bitb_78_92 gnd C_bl
Rb_78_93 bit_78_93 bit_78_94 R_bl
Rbb_78_93 bitb_78_93 bitb_78_94 R_bl
Cb_78_93 bit_78_93 gnd C_bl
Cbb_78_93 bitb_78_93 gnd C_bl
Rb_78_94 bit_78_94 bit_78_95 R_bl
Rbb_78_94 bitb_78_94 bitb_78_95 R_bl
Cb_78_94 bit_78_94 gnd C_bl
Cbb_78_94 bitb_78_94 gnd C_bl
Rb_78_95 bit_78_95 bit_78_96 R_bl
Rbb_78_95 bitb_78_95 bitb_78_96 R_bl
Cb_78_95 bit_78_95 gnd C_bl
Cbb_78_95 bitb_78_95 gnd C_bl
Rb_78_96 bit_78_96 bit_78_97 R_bl
Rbb_78_96 bitb_78_96 bitb_78_97 R_bl
Cb_78_96 bit_78_96 gnd C_bl
Cbb_78_96 bitb_78_96 gnd C_bl
Rb_78_97 bit_78_97 bit_78_98 R_bl
Rbb_78_97 bitb_78_97 bitb_78_98 R_bl
Cb_78_97 bit_78_97 gnd C_bl
Cbb_78_97 bitb_78_97 gnd C_bl
Rb_78_98 bit_78_98 bit_78_99 R_bl
Rbb_78_98 bitb_78_98 bitb_78_99 R_bl
Cb_78_98 bit_78_98 gnd C_bl
Cbb_78_98 bitb_78_98 gnd C_bl
Rb_78_99 bit_78_99 bit_78_100 R_bl
Rbb_78_99 bitb_78_99 bitb_78_100 R_bl
Cb_78_99 bit_78_99 gnd C_bl
Cbb_78_99 bitb_78_99 gnd C_bl
Rb_79_0 bit_79_0 bit_79_1 R_bl
Rbb_79_0 bitb_79_0 bitb_79_1 R_bl
Cb_79_0 bit_79_0 gnd C_bl
Cbb_79_0 bitb_79_0 gnd C_bl
Rb_79_1 bit_79_1 bit_79_2 R_bl
Rbb_79_1 bitb_79_1 bitb_79_2 R_bl
Cb_79_1 bit_79_1 gnd C_bl
Cbb_79_1 bitb_79_1 gnd C_bl
Rb_79_2 bit_79_2 bit_79_3 R_bl
Rbb_79_2 bitb_79_2 bitb_79_3 R_bl
Cb_79_2 bit_79_2 gnd C_bl
Cbb_79_2 bitb_79_2 gnd C_bl
Rb_79_3 bit_79_3 bit_79_4 R_bl
Rbb_79_3 bitb_79_3 bitb_79_4 R_bl
Cb_79_3 bit_79_3 gnd C_bl
Cbb_79_3 bitb_79_3 gnd C_bl
Rb_79_4 bit_79_4 bit_79_5 R_bl
Rbb_79_4 bitb_79_4 bitb_79_5 R_bl
Cb_79_4 bit_79_4 gnd C_bl
Cbb_79_4 bitb_79_4 gnd C_bl
Rb_79_5 bit_79_5 bit_79_6 R_bl
Rbb_79_5 bitb_79_5 bitb_79_6 R_bl
Cb_79_5 bit_79_5 gnd C_bl
Cbb_79_5 bitb_79_5 gnd C_bl
Rb_79_6 bit_79_6 bit_79_7 R_bl
Rbb_79_6 bitb_79_6 bitb_79_7 R_bl
Cb_79_6 bit_79_6 gnd C_bl
Cbb_79_6 bitb_79_6 gnd C_bl
Rb_79_7 bit_79_7 bit_79_8 R_bl
Rbb_79_7 bitb_79_7 bitb_79_8 R_bl
Cb_79_7 bit_79_7 gnd C_bl
Cbb_79_7 bitb_79_7 gnd C_bl
Rb_79_8 bit_79_8 bit_79_9 R_bl
Rbb_79_8 bitb_79_8 bitb_79_9 R_bl
Cb_79_8 bit_79_8 gnd C_bl
Cbb_79_8 bitb_79_8 gnd C_bl
Rb_79_9 bit_79_9 bit_79_10 R_bl
Rbb_79_9 bitb_79_9 bitb_79_10 R_bl
Cb_79_9 bit_79_9 gnd C_bl
Cbb_79_9 bitb_79_9 gnd C_bl
Rb_79_10 bit_79_10 bit_79_11 R_bl
Rbb_79_10 bitb_79_10 bitb_79_11 R_bl
Cb_79_10 bit_79_10 gnd C_bl
Cbb_79_10 bitb_79_10 gnd C_bl
Rb_79_11 bit_79_11 bit_79_12 R_bl
Rbb_79_11 bitb_79_11 bitb_79_12 R_bl
Cb_79_11 bit_79_11 gnd C_bl
Cbb_79_11 bitb_79_11 gnd C_bl
Rb_79_12 bit_79_12 bit_79_13 R_bl
Rbb_79_12 bitb_79_12 bitb_79_13 R_bl
Cb_79_12 bit_79_12 gnd C_bl
Cbb_79_12 bitb_79_12 gnd C_bl
Rb_79_13 bit_79_13 bit_79_14 R_bl
Rbb_79_13 bitb_79_13 bitb_79_14 R_bl
Cb_79_13 bit_79_13 gnd C_bl
Cbb_79_13 bitb_79_13 gnd C_bl
Rb_79_14 bit_79_14 bit_79_15 R_bl
Rbb_79_14 bitb_79_14 bitb_79_15 R_bl
Cb_79_14 bit_79_14 gnd C_bl
Cbb_79_14 bitb_79_14 gnd C_bl
Rb_79_15 bit_79_15 bit_79_16 R_bl
Rbb_79_15 bitb_79_15 bitb_79_16 R_bl
Cb_79_15 bit_79_15 gnd C_bl
Cbb_79_15 bitb_79_15 gnd C_bl
Rb_79_16 bit_79_16 bit_79_17 R_bl
Rbb_79_16 bitb_79_16 bitb_79_17 R_bl
Cb_79_16 bit_79_16 gnd C_bl
Cbb_79_16 bitb_79_16 gnd C_bl
Rb_79_17 bit_79_17 bit_79_18 R_bl
Rbb_79_17 bitb_79_17 bitb_79_18 R_bl
Cb_79_17 bit_79_17 gnd C_bl
Cbb_79_17 bitb_79_17 gnd C_bl
Rb_79_18 bit_79_18 bit_79_19 R_bl
Rbb_79_18 bitb_79_18 bitb_79_19 R_bl
Cb_79_18 bit_79_18 gnd C_bl
Cbb_79_18 bitb_79_18 gnd C_bl
Rb_79_19 bit_79_19 bit_79_20 R_bl
Rbb_79_19 bitb_79_19 bitb_79_20 R_bl
Cb_79_19 bit_79_19 gnd C_bl
Cbb_79_19 bitb_79_19 gnd C_bl
Rb_79_20 bit_79_20 bit_79_21 R_bl
Rbb_79_20 bitb_79_20 bitb_79_21 R_bl
Cb_79_20 bit_79_20 gnd C_bl
Cbb_79_20 bitb_79_20 gnd C_bl
Rb_79_21 bit_79_21 bit_79_22 R_bl
Rbb_79_21 bitb_79_21 bitb_79_22 R_bl
Cb_79_21 bit_79_21 gnd C_bl
Cbb_79_21 bitb_79_21 gnd C_bl
Rb_79_22 bit_79_22 bit_79_23 R_bl
Rbb_79_22 bitb_79_22 bitb_79_23 R_bl
Cb_79_22 bit_79_22 gnd C_bl
Cbb_79_22 bitb_79_22 gnd C_bl
Rb_79_23 bit_79_23 bit_79_24 R_bl
Rbb_79_23 bitb_79_23 bitb_79_24 R_bl
Cb_79_23 bit_79_23 gnd C_bl
Cbb_79_23 bitb_79_23 gnd C_bl
Rb_79_24 bit_79_24 bit_79_25 R_bl
Rbb_79_24 bitb_79_24 bitb_79_25 R_bl
Cb_79_24 bit_79_24 gnd C_bl
Cbb_79_24 bitb_79_24 gnd C_bl
Rb_79_25 bit_79_25 bit_79_26 R_bl
Rbb_79_25 bitb_79_25 bitb_79_26 R_bl
Cb_79_25 bit_79_25 gnd C_bl
Cbb_79_25 bitb_79_25 gnd C_bl
Rb_79_26 bit_79_26 bit_79_27 R_bl
Rbb_79_26 bitb_79_26 bitb_79_27 R_bl
Cb_79_26 bit_79_26 gnd C_bl
Cbb_79_26 bitb_79_26 gnd C_bl
Rb_79_27 bit_79_27 bit_79_28 R_bl
Rbb_79_27 bitb_79_27 bitb_79_28 R_bl
Cb_79_27 bit_79_27 gnd C_bl
Cbb_79_27 bitb_79_27 gnd C_bl
Rb_79_28 bit_79_28 bit_79_29 R_bl
Rbb_79_28 bitb_79_28 bitb_79_29 R_bl
Cb_79_28 bit_79_28 gnd C_bl
Cbb_79_28 bitb_79_28 gnd C_bl
Rb_79_29 bit_79_29 bit_79_30 R_bl
Rbb_79_29 bitb_79_29 bitb_79_30 R_bl
Cb_79_29 bit_79_29 gnd C_bl
Cbb_79_29 bitb_79_29 gnd C_bl
Rb_79_30 bit_79_30 bit_79_31 R_bl
Rbb_79_30 bitb_79_30 bitb_79_31 R_bl
Cb_79_30 bit_79_30 gnd C_bl
Cbb_79_30 bitb_79_30 gnd C_bl
Rb_79_31 bit_79_31 bit_79_32 R_bl
Rbb_79_31 bitb_79_31 bitb_79_32 R_bl
Cb_79_31 bit_79_31 gnd C_bl
Cbb_79_31 bitb_79_31 gnd C_bl
Rb_79_32 bit_79_32 bit_79_33 R_bl
Rbb_79_32 bitb_79_32 bitb_79_33 R_bl
Cb_79_32 bit_79_32 gnd C_bl
Cbb_79_32 bitb_79_32 gnd C_bl
Rb_79_33 bit_79_33 bit_79_34 R_bl
Rbb_79_33 bitb_79_33 bitb_79_34 R_bl
Cb_79_33 bit_79_33 gnd C_bl
Cbb_79_33 bitb_79_33 gnd C_bl
Rb_79_34 bit_79_34 bit_79_35 R_bl
Rbb_79_34 bitb_79_34 bitb_79_35 R_bl
Cb_79_34 bit_79_34 gnd C_bl
Cbb_79_34 bitb_79_34 gnd C_bl
Rb_79_35 bit_79_35 bit_79_36 R_bl
Rbb_79_35 bitb_79_35 bitb_79_36 R_bl
Cb_79_35 bit_79_35 gnd C_bl
Cbb_79_35 bitb_79_35 gnd C_bl
Rb_79_36 bit_79_36 bit_79_37 R_bl
Rbb_79_36 bitb_79_36 bitb_79_37 R_bl
Cb_79_36 bit_79_36 gnd C_bl
Cbb_79_36 bitb_79_36 gnd C_bl
Rb_79_37 bit_79_37 bit_79_38 R_bl
Rbb_79_37 bitb_79_37 bitb_79_38 R_bl
Cb_79_37 bit_79_37 gnd C_bl
Cbb_79_37 bitb_79_37 gnd C_bl
Rb_79_38 bit_79_38 bit_79_39 R_bl
Rbb_79_38 bitb_79_38 bitb_79_39 R_bl
Cb_79_38 bit_79_38 gnd C_bl
Cbb_79_38 bitb_79_38 gnd C_bl
Rb_79_39 bit_79_39 bit_79_40 R_bl
Rbb_79_39 bitb_79_39 bitb_79_40 R_bl
Cb_79_39 bit_79_39 gnd C_bl
Cbb_79_39 bitb_79_39 gnd C_bl
Rb_79_40 bit_79_40 bit_79_41 R_bl
Rbb_79_40 bitb_79_40 bitb_79_41 R_bl
Cb_79_40 bit_79_40 gnd C_bl
Cbb_79_40 bitb_79_40 gnd C_bl
Rb_79_41 bit_79_41 bit_79_42 R_bl
Rbb_79_41 bitb_79_41 bitb_79_42 R_bl
Cb_79_41 bit_79_41 gnd C_bl
Cbb_79_41 bitb_79_41 gnd C_bl
Rb_79_42 bit_79_42 bit_79_43 R_bl
Rbb_79_42 bitb_79_42 bitb_79_43 R_bl
Cb_79_42 bit_79_42 gnd C_bl
Cbb_79_42 bitb_79_42 gnd C_bl
Rb_79_43 bit_79_43 bit_79_44 R_bl
Rbb_79_43 bitb_79_43 bitb_79_44 R_bl
Cb_79_43 bit_79_43 gnd C_bl
Cbb_79_43 bitb_79_43 gnd C_bl
Rb_79_44 bit_79_44 bit_79_45 R_bl
Rbb_79_44 bitb_79_44 bitb_79_45 R_bl
Cb_79_44 bit_79_44 gnd C_bl
Cbb_79_44 bitb_79_44 gnd C_bl
Rb_79_45 bit_79_45 bit_79_46 R_bl
Rbb_79_45 bitb_79_45 bitb_79_46 R_bl
Cb_79_45 bit_79_45 gnd C_bl
Cbb_79_45 bitb_79_45 gnd C_bl
Rb_79_46 bit_79_46 bit_79_47 R_bl
Rbb_79_46 bitb_79_46 bitb_79_47 R_bl
Cb_79_46 bit_79_46 gnd C_bl
Cbb_79_46 bitb_79_46 gnd C_bl
Rb_79_47 bit_79_47 bit_79_48 R_bl
Rbb_79_47 bitb_79_47 bitb_79_48 R_bl
Cb_79_47 bit_79_47 gnd C_bl
Cbb_79_47 bitb_79_47 gnd C_bl
Rb_79_48 bit_79_48 bit_79_49 R_bl
Rbb_79_48 bitb_79_48 bitb_79_49 R_bl
Cb_79_48 bit_79_48 gnd C_bl
Cbb_79_48 bitb_79_48 gnd C_bl
Rb_79_49 bit_79_49 bit_79_50 R_bl
Rbb_79_49 bitb_79_49 bitb_79_50 R_bl
Cb_79_49 bit_79_49 gnd C_bl
Cbb_79_49 bitb_79_49 gnd C_bl
Rb_79_50 bit_79_50 bit_79_51 R_bl
Rbb_79_50 bitb_79_50 bitb_79_51 R_bl
Cb_79_50 bit_79_50 gnd C_bl
Cbb_79_50 bitb_79_50 gnd C_bl
Rb_79_51 bit_79_51 bit_79_52 R_bl
Rbb_79_51 bitb_79_51 bitb_79_52 R_bl
Cb_79_51 bit_79_51 gnd C_bl
Cbb_79_51 bitb_79_51 gnd C_bl
Rb_79_52 bit_79_52 bit_79_53 R_bl
Rbb_79_52 bitb_79_52 bitb_79_53 R_bl
Cb_79_52 bit_79_52 gnd C_bl
Cbb_79_52 bitb_79_52 gnd C_bl
Rb_79_53 bit_79_53 bit_79_54 R_bl
Rbb_79_53 bitb_79_53 bitb_79_54 R_bl
Cb_79_53 bit_79_53 gnd C_bl
Cbb_79_53 bitb_79_53 gnd C_bl
Rb_79_54 bit_79_54 bit_79_55 R_bl
Rbb_79_54 bitb_79_54 bitb_79_55 R_bl
Cb_79_54 bit_79_54 gnd C_bl
Cbb_79_54 bitb_79_54 gnd C_bl
Rb_79_55 bit_79_55 bit_79_56 R_bl
Rbb_79_55 bitb_79_55 bitb_79_56 R_bl
Cb_79_55 bit_79_55 gnd C_bl
Cbb_79_55 bitb_79_55 gnd C_bl
Rb_79_56 bit_79_56 bit_79_57 R_bl
Rbb_79_56 bitb_79_56 bitb_79_57 R_bl
Cb_79_56 bit_79_56 gnd C_bl
Cbb_79_56 bitb_79_56 gnd C_bl
Rb_79_57 bit_79_57 bit_79_58 R_bl
Rbb_79_57 bitb_79_57 bitb_79_58 R_bl
Cb_79_57 bit_79_57 gnd C_bl
Cbb_79_57 bitb_79_57 gnd C_bl
Rb_79_58 bit_79_58 bit_79_59 R_bl
Rbb_79_58 bitb_79_58 bitb_79_59 R_bl
Cb_79_58 bit_79_58 gnd C_bl
Cbb_79_58 bitb_79_58 gnd C_bl
Rb_79_59 bit_79_59 bit_79_60 R_bl
Rbb_79_59 bitb_79_59 bitb_79_60 R_bl
Cb_79_59 bit_79_59 gnd C_bl
Cbb_79_59 bitb_79_59 gnd C_bl
Rb_79_60 bit_79_60 bit_79_61 R_bl
Rbb_79_60 bitb_79_60 bitb_79_61 R_bl
Cb_79_60 bit_79_60 gnd C_bl
Cbb_79_60 bitb_79_60 gnd C_bl
Rb_79_61 bit_79_61 bit_79_62 R_bl
Rbb_79_61 bitb_79_61 bitb_79_62 R_bl
Cb_79_61 bit_79_61 gnd C_bl
Cbb_79_61 bitb_79_61 gnd C_bl
Rb_79_62 bit_79_62 bit_79_63 R_bl
Rbb_79_62 bitb_79_62 bitb_79_63 R_bl
Cb_79_62 bit_79_62 gnd C_bl
Cbb_79_62 bitb_79_62 gnd C_bl
Rb_79_63 bit_79_63 bit_79_64 R_bl
Rbb_79_63 bitb_79_63 bitb_79_64 R_bl
Cb_79_63 bit_79_63 gnd C_bl
Cbb_79_63 bitb_79_63 gnd C_bl
Rb_79_64 bit_79_64 bit_79_65 R_bl
Rbb_79_64 bitb_79_64 bitb_79_65 R_bl
Cb_79_64 bit_79_64 gnd C_bl
Cbb_79_64 bitb_79_64 gnd C_bl
Rb_79_65 bit_79_65 bit_79_66 R_bl
Rbb_79_65 bitb_79_65 bitb_79_66 R_bl
Cb_79_65 bit_79_65 gnd C_bl
Cbb_79_65 bitb_79_65 gnd C_bl
Rb_79_66 bit_79_66 bit_79_67 R_bl
Rbb_79_66 bitb_79_66 bitb_79_67 R_bl
Cb_79_66 bit_79_66 gnd C_bl
Cbb_79_66 bitb_79_66 gnd C_bl
Rb_79_67 bit_79_67 bit_79_68 R_bl
Rbb_79_67 bitb_79_67 bitb_79_68 R_bl
Cb_79_67 bit_79_67 gnd C_bl
Cbb_79_67 bitb_79_67 gnd C_bl
Rb_79_68 bit_79_68 bit_79_69 R_bl
Rbb_79_68 bitb_79_68 bitb_79_69 R_bl
Cb_79_68 bit_79_68 gnd C_bl
Cbb_79_68 bitb_79_68 gnd C_bl
Rb_79_69 bit_79_69 bit_79_70 R_bl
Rbb_79_69 bitb_79_69 bitb_79_70 R_bl
Cb_79_69 bit_79_69 gnd C_bl
Cbb_79_69 bitb_79_69 gnd C_bl
Rb_79_70 bit_79_70 bit_79_71 R_bl
Rbb_79_70 bitb_79_70 bitb_79_71 R_bl
Cb_79_70 bit_79_70 gnd C_bl
Cbb_79_70 bitb_79_70 gnd C_bl
Rb_79_71 bit_79_71 bit_79_72 R_bl
Rbb_79_71 bitb_79_71 bitb_79_72 R_bl
Cb_79_71 bit_79_71 gnd C_bl
Cbb_79_71 bitb_79_71 gnd C_bl
Rb_79_72 bit_79_72 bit_79_73 R_bl
Rbb_79_72 bitb_79_72 bitb_79_73 R_bl
Cb_79_72 bit_79_72 gnd C_bl
Cbb_79_72 bitb_79_72 gnd C_bl
Rb_79_73 bit_79_73 bit_79_74 R_bl
Rbb_79_73 bitb_79_73 bitb_79_74 R_bl
Cb_79_73 bit_79_73 gnd C_bl
Cbb_79_73 bitb_79_73 gnd C_bl
Rb_79_74 bit_79_74 bit_79_75 R_bl
Rbb_79_74 bitb_79_74 bitb_79_75 R_bl
Cb_79_74 bit_79_74 gnd C_bl
Cbb_79_74 bitb_79_74 gnd C_bl
Rb_79_75 bit_79_75 bit_79_76 R_bl
Rbb_79_75 bitb_79_75 bitb_79_76 R_bl
Cb_79_75 bit_79_75 gnd C_bl
Cbb_79_75 bitb_79_75 gnd C_bl
Rb_79_76 bit_79_76 bit_79_77 R_bl
Rbb_79_76 bitb_79_76 bitb_79_77 R_bl
Cb_79_76 bit_79_76 gnd C_bl
Cbb_79_76 bitb_79_76 gnd C_bl
Rb_79_77 bit_79_77 bit_79_78 R_bl
Rbb_79_77 bitb_79_77 bitb_79_78 R_bl
Cb_79_77 bit_79_77 gnd C_bl
Cbb_79_77 bitb_79_77 gnd C_bl
Rb_79_78 bit_79_78 bit_79_79 R_bl
Rbb_79_78 bitb_79_78 bitb_79_79 R_bl
Cb_79_78 bit_79_78 gnd C_bl
Cbb_79_78 bitb_79_78 gnd C_bl
Rb_79_79 bit_79_79 bit_79_80 R_bl
Rbb_79_79 bitb_79_79 bitb_79_80 R_bl
Cb_79_79 bit_79_79 gnd C_bl
Cbb_79_79 bitb_79_79 gnd C_bl
Rb_79_80 bit_79_80 bit_79_81 R_bl
Rbb_79_80 bitb_79_80 bitb_79_81 R_bl
Cb_79_80 bit_79_80 gnd C_bl
Cbb_79_80 bitb_79_80 gnd C_bl
Rb_79_81 bit_79_81 bit_79_82 R_bl
Rbb_79_81 bitb_79_81 bitb_79_82 R_bl
Cb_79_81 bit_79_81 gnd C_bl
Cbb_79_81 bitb_79_81 gnd C_bl
Rb_79_82 bit_79_82 bit_79_83 R_bl
Rbb_79_82 bitb_79_82 bitb_79_83 R_bl
Cb_79_82 bit_79_82 gnd C_bl
Cbb_79_82 bitb_79_82 gnd C_bl
Rb_79_83 bit_79_83 bit_79_84 R_bl
Rbb_79_83 bitb_79_83 bitb_79_84 R_bl
Cb_79_83 bit_79_83 gnd C_bl
Cbb_79_83 bitb_79_83 gnd C_bl
Rb_79_84 bit_79_84 bit_79_85 R_bl
Rbb_79_84 bitb_79_84 bitb_79_85 R_bl
Cb_79_84 bit_79_84 gnd C_bl
Cbb_79_84 bitb_79_84 gnd C_bl
Rb_79_85 bit_79_85 bit_79_86 R_bl
Rbb_79_85 bitb_79_85 bitb_79_86 R_bl
Cb_79_85 bit_79_85 gnd C_bl
Cbb_79_85 bitb_79_85 gnd C_bl
Rb_79_86 bit_79_86 bit_79_87 R_bl
Rbb_79_86 bitb_79_86 bitb_79_87 R_bl
Cb_79_86 bit_79_86 gnd C_bl
Cbb_79_86 bitb_79_86 gnd C_bl
Rb_79_87 bit_79_87 bit_79_88 R_bl
Rbb_79_87 bitb_79_87 bitb_79_88 R_bl
Cb_79_87 bit_79_87 gnd C_bl
Cbb_79_87 bitb_79_87 gnd C_bl
Rb_79_88 bit_79_88 bit_79_89 R_bl
Rbb_79_88 bitb_79_88 bitb_79_89 R_bl
Cb_79_88 bit_79_88 gnd C_bl
Cbb_79_88 bitb_79_88 gnd C_bl
Rb_79_89 bit_79_89 bit_79_90 R_bl
Rbb_79_89 bitb_79_89 bitb_79_90 R_bl
Cb_79_89 bit_79_89 gnd C_bl
Cbb_79_89 bitb_79_89 gnd C_bl
Rb_79_90 bit_79_90 bit_79_91 R_bl
Rbb_79_90 bitb_79_90 bitb_79_91 R_bl
Cb_79_90 bit_79_90 gnd C_bl
Cbb_79_90 bitb_79_90 gnd C_bl
Rb_79_91 bit_79_91 bit_79_92 R_bl
Rbb_79_91 bitb_79_91 bitb_79_92 R_bl
Cb_79_91 bit_79_91 gnd C_bl
Cbb_79_91 bitb_79_91 gnd C_bl
Rb_79_92 bit_79_92 bit_79_93 R_bl
Rbb_79_92 bitb_79_92 bitb_79_93 R_bl
Cb_79_92 bit_79_92 gnd C_bl
Cbb_79_92 bitb_79_92 gnd C_bl
Rb_79_93 bit_79_93 bit_79_94 R_bl
Rbb_79_93 bitb_79_93 bitb_79_94 R_bl
Cb_79_93 bit_79_93 gnd C_bl
Cbb_79_93 bitb_79_93 gnd C_bl
Rb_79_94 bit_79_94 bit_79_95 R_bl
Rbb_79_94 bitb_79_94 bitb_79_95 R_bl
Cb_79_94 bit_79_94 gnd C_bl
Cbb_79_94 bitb_79_94 gnd C_bl
Rb_79_95 bit_79_95 bit_79_96 R_bl
Rbb_79_95 bitb_79_95 bitb_79_96 R_bl
Cb_79_95 bit_79_95 gnd C_bl
Cbb_79_95 bitb_79_95 gnd C_bl
Rb_79_96 bit_79_96 bit_79_97 R_bl
Rbb_79_96 bitb_79_96 bitb_79_97 R_bl
Cb_79_96 bit_79_96 gnd C_bl
Cbb_79_96 bitb_79_96 gnd C_bl
Rb_79_97 bit_79_97 bit_79_98 R_bl
Rbb_79_97 bitb_79_97 bitb_79_98 R_bl
Cb_79_97 bit_79_97 gnd C_bl
Cbb_79_97 bitb_79_97 gnd C_bl
Rb_79_98 bit_79_98 bit_79_99 R_bl
Rbb_79_98 bitb_79_98 bitb_79_99 R_bl
Cb_79_98 bit_79_98 gnd C_bl
Cbb_79_98 bitb_79_98 gnd C_bl
Rb_79_99 bit_79_99 bit_79_100 R_bl
Rbb_79_99 bitb_79_99 bitb_79_100 R_bl
Cb_79_99 bit_79_99 gnd C_bl
Cbb_79_99 bitb_79_99 gnd C_bl
Rb_80_0 bit_80_0 bit_80_1 R_bl
Rbb_80_0 bitb_80_0 bitb_80_1 R_bl
Cb_80_0 bit_80_0 gnd C_bl
Cbb_80_0 bitb_80_0 gnd C_bl
Rb_80_1 bit_80_1 bit_80_2 R_bl
Rbb_80_1 bitb_80_1 bitb_80_2 R_bl
Cb_80_1 bit_80_1 gnd C_bl
Cbb_80_1 bitb_80_1 gnd C_bl
Rb_80_2 bit_80_2 bit_80_3 R_bl
Rbb_80_2 bitb_80_2 bitb_80_3 R_bl
Cb_80_2 bit_80_2 gnd C_bl
Cbb_80_2 bitb_80_2 gnd C_bl
Rb_80_3 bit_80_3 bit_80_4 R_bl
Rbb_80_3 bitb_80_3 bitb_80_4 R_bl
Cb_80_3 bit_80_3 gnd C_bl
Cbb_80_3 bitb_80_3 gnd C_bl
Rb_80_4 bit_80_4 bit_80_5 R_bl
Rbb_80_4 bitb_80_4 bitb_80_5 R_bl
Cb_80_4 bit_80_4 gnd C_bl
Cbb_80_4 bitb_80_4 gnd C_bl
Rb_80_5 bit_80_5 bit_80_6 R_bl
Rbb_80_5 bitb_80_5 bitb_80_6 R_bl
Cb_80_5 bit_80_5 gnd C_bl
Cbb_80_5 bitb_80_5 gnd C_bl
Rb_80_6 bit_80_6 bit_80_7 R_bl
Rbb_80_6 bitb_80_6 bitb_80_7 R_bl
Cb_80_6 bit_80_6 gnd C_bl
Cbb_80_6 bitb_80_6 gnd C_bl
Rb_80_7 bit_80_7 bit_80_8 R_bl
Rbb_80_7 bitb_80_7 bitb_80_8 R_bl
Cb_80_7 bit_80_7 gnd C_bl
Cbb_80_7 bitb_80_7 gnd C_bl
Rb_80_8 bit_80_8 bit_80_9 R_bl
Rbb_80_8 bitb_80_8 bitb_80_9 R_bl
Cb_80_8 bit_80_8 gnd C_bl
Cbb_80_8 bitb_80_8 gnd C_bl
Rb_80_9 bit_80_9 bit_80_10 R_bl
Rbb_80_9 bitb_80_9 bitb_80_10 R_bl
Cb_80_9 bit_80_9 gnd C_bl
Cbb_80_9 bitb_80_9 gnd C_bl
Rb_80_10 bit_80_10 bit_80_11 R_bl
Rbb_80_10 bitb_80_10 bitb_80_11 R_bl
Cb_80_10 bit_80_10 gnd C_bl
Cbb_80_10 bitb_80_10 gnd C_bl
Rb_80_11 bit_80_11 bit_80_12 R_bl
Rbb_80_11 bitb_80_11 bitb_80_12 R_bl
Cb_80_11 bit_80_11 gnd C_bl
Cbb_80_11 bitb_80_11 gnd C_bl
Rb_80_12 bit_80_12 bit_80_13 R_bl
Rbb_80_12 bitb_80_12 bitb_80_13 R_bl
Cb_80_12 bit_80_12 gnd C_bl
Cbb_80_12 bitb_80_12 gnd C_bl
Rb_80_13 bit_80_13 bit_80_14 R_bl
Rbb_80_13 bitb_80_13 bitb_80_14 R_bl
Cb_80_13 bit_80_13 gnd C_bl
Cbb_80_13 bitb_80_13 gnd C_bl
Rb_80_14 bit_80_14 bit_80_15 R_bl
Rbb_80_14 bitb_80_14 bitb_80_15 R_bl
Cb_80_14 bit_80_14 gnd C_bl
Cbb_80_14 bitb_80_14 gnd C_bl
Rb_80_15 bit_80_15 bit_80_16 R_bl
Rbb_80_15 bitb_80_15 bitb_80_16 R_bl
Cb_80_15 bit_80_15 gnd C_bl
Cbb_80_15 bitb_80_15 gnd C_bl
Rb_80_16 bit_80_16 bit_80_17 R_bl
Rbb_80_16 bitb_80_16 bitb_80_17 R_bl
Cb_80_16 bit_80_16 gnd C_bl
Cbb_80_16 bitb_80_16 gnd C_bl
Rb_80_17 bit_80_17 bit_80_18 R_bl
Rbb_80_17 bitb_80_17 bitb_80_18 R_bl
Cb_80_17 bit_80_17 gnd C_bl
Cbb_80_17 bitb_80_17 gnd C_bl
Rb_80_18 bit_80_18 bit_80_19 R_bl
Rbb_80_18 bitb_80_18 bitb_80_19 R_bl
Cb_80_18 bit_80_18 gnd C_bl
Cbb_80_18 bitb_80_18 gnd C_bl
Rb_80_19 bit_80_19 bit_80_20 R_bl
Rbb_80_19 bitb_80_19 bitb_80_20 R_bl
Cb_80_19 bit_80_19 gnd C_bl
Cbb_80_19 bitb_80_19 gnd C_bl
Rb_80_20 bit_80_20 bit_80_21 R_bl
Rbb_80_20 bitb_80_20 bitb_80_21 R_bl
Cb_80_20 bit_80_20 gnd C_bl
Cbb_80_20 bitb_80_20 gnd C_bl
Rb_80_21 bit_80_21 bit_80_22 R_bl
Rbb_80_21 bitb_80_21 bitb_80_22 R_bl
Cb_80_21 bit_80_21 gnd C_bl
Cbb_80_21 bitb_80_21 gnd C_bl
Rb_80_22 bit_80_22 bit_80_23 R_bl
Rbb_80_22 bitb_80_22 bitb_80_23 R_bl
Cb_80_22 bit_80_22 gnd C_bl
Cbb_80_22 bitb_80_22 gnd C_bl
Rb_80_23 bit_80_23 bit_80_24 R_bl
Rbb_80_23 bitb_80_23 bitb_80_24 R_bl
Cb_80_23 bit_80_23 gnd C_bl
Cbb_80_23 bitb_80_23 gnd C_bl
Rb_80_24 bit_80_24 bit_80_25 R_bl
Rbb_80_24 bitb_80_24 bitb_80_25 R_bl
Cb_80_24 bit_80_24 gnd C_bl
Cbb_80_24 bitb_80_24 gnd C_bl
Rb_80_25 bit_80_25 bit_80_26 R_bl
Rbb_80_25 bitb_80_25 bitb_80_26 R_bl
Cb_80_25 bit_80_25 gnd C_bl
Cbb_80_25 bitb_80_25 gnd C_bl
Rb_80_26 bit_80_26 bit_80_27 R_bl
Rbb_80_26 bitb_80_26 bitb_80_27 R_bl
Cb_80_26 bit_80_26 gnd C_bl
Cbb_80_26 bitb_80_26 gnd C_bl
Rb_80_27 bit_80_27 bit_80_28 R_bl
Rbb_80_27 bitb_80_27 bitb_80_28 R_bl
Cb_80_27 bit_80_27 gnd C_bl
Cbb_80_27 bitb_80_27 gnd C_bl
Rb_80_28 bit_80_28 bit_80_29 R_bl
Rbb_80_28 bitb_80_28 bitb_80_29 R_bl
Cb_80_28 bit_80_28 gnd C_bl
Cbb_80_28 bitb_80_28 gnd C_bl
Rb_80_29 bit_80_29 bit_80_30 R_bl
Rbb_80_29 bitb_80_29 bitb_80_30 R_bl
Cb_80_29 bit_80_29 gnd C_bl
Cbb_80_29 bitb_80_29 gnd C_bl
Rb_80_30 bit_80_30 bit_80_31 R_bl
Rbb_80_30 bitb_80_30 bitb_80_31 R_bl
Cb_80_30 bit_80_30 gnd C_bl
Cbb_80_30 bitb_80_30 gnd C_bl
Rb_80_31 bit_80_31 bit_80_32 R_bl
Rbb_80_31 bitb_80_31 bitb_80_32 R_bl
Cb_80_31 bit_80_31 gnd C_bl
Cbb_80_31 bitb_80_31 gnd C_bl
Rb_80_32 bit_80_32 bit_80_33 R_bl
Rbb_80_32 bitb_80_32 bitb_80_33 R_bl
Cb_80_32 bit_80_32 gnd C_bl
Cbb_80_32 bitb_80_32 gnd C_bl
Rb_80_33 bit_80_33 bit_80_34 R_bl
Rbb_80_33 bitb_80_33 bitb_80_34 R_bl
Cb_80_33 bit_80_33 gnd C_bl
Cbb_80_33 bitb_80_33 gnd C_bl
Rb_80_34 bit_80_34 bit_80_35 R_bl
Rbb_80_34 bitb_80_34 bitb_80_35 R_bl
Cb_80_34 bit_80_34 gnd C_bl
Cbb_80_34 bitb_80_34 gnd C_bl
Rb_80_35 bit_80_35 bit_80_36 R_bl
Rbb_80_35 bitb_80_35 bitb_80_36 R_bl
Cb_80_35 bit_80_35 gnd C_bl
Cbb_80_35 bitb_80_35 gnd C_bl
Rb_80_36 bit_80_36 bit_80_37 R_bl
Rbb_80_36 bitb_80_36 bitb_80_37 R_bl
Cb_80_36 bit_80_36 gnd C_bl
Cbb_80_36 bitb_80_36 gnd C_bl
Rb_80_37 bit_80_37 bit_80_38 R_bl
Rbb_80_37 bitb_80_37 bitb_80_38 R_bl
Cb_80_37 bit_80_37 gnd C_bl
Cbb_80_37 bitb_80_37 gnd C_bl
Rb_80_38 bit_80_38 bit_80_39 R_bl
Rbb_80_38 bitb_80_38 bitb_80_39 R_bl
Cb_80_38 bit_80_38 gnd C_bl
Cbb_80_38 bitb_80_38 gnd C_bl
Rb_80_39 bit_80_39 bit_80_40 R_bl
Rbb_80_39 bitb_80_39 bitb_80_40 R_bl
Cb_80_39 bit_80_39 gnd C_bl
Cbb_80_39 bitb_80_39 gnd C_bl
Rb_80_40 bit_80_40 bit_80_41 R_bl
Rbb_80_40 bitb_80_40 bitb_80_41 R_bl
Cb_80_40 bit_80_40 gnd C_bl
Cbb_80_40 bitb_80_40 gnd C_bl
Rb_80_41 bit_80_41 bit_80_42 R_bl
Rbb_80_41 bitb_80_41 bitb_80_42 R_bl
Cb_80_41 bit_80_41 gnd C_bl
Cbb_80_41 bitb_80_41 gnd C_bl
Rb_80_42 bit_80_42 bit_80_43 R_bl
Rbb_80_42 bitb_80_42 bitb_80_43 R_bl
Cb_80_42 bit_80_42 gnd C_bl
Cbb_80_42 bitb_80_42 gnd C_bl
Rb_80_43 bit_80_43 bit_80_44 R_bl
Rbb_80_43 bitb_80_43 bitb_80_44 R_bl
Cb_80_43 bit_80_43 gnd C_bl
Cbb_80_43 bitb_80_43 gnd C_bl
Rb_80_44 bit_80_44 bit_80_45 R_bl
Rbb_80_44 bitb_80_44 bitb_80_45 R_bl
Cb_80_44 bit_80_44 gnd C_bl
Cbb_80_44 bitb_80_44 gnd C_bl
Rb_80_45 bit_80_45 bit_80_46 R_bl
Rbb_80_45 bitb_80_45 bitb_80_46 R_bl
Cb_80_45 bit_80_45 gnd C_bl
Cbb_80_45 bitb_80_45 gnd C_bl
Rb_80_46 bit_80_46 bit_80_47 R_bl
Rbb_80_46 bitb_80_46 bitb_80_47 R_bl
Cb_80_46 bit_80_46 gnd C_bl
Cbb_80_46 bitb_80_46 gnd C_bl
Rb_80_47 bit_80_47 bit_80_48 R_bl
Rbb_80_47 bitb_80_47 bitb_80_48 R_bl
Cb_80_47 bit_80_47 gnd C_bl
Cbb_80_47 bitb_80_47 gnd C_bl
Rb_80_48 bit_80_48 bit_80_49 R_bl
Rbb_80_48 bitb_80_48 bitb_80_49 R_bl
Cb_80_48 bit_80_48 gnd C_bl
Cbb_80_48 bitb_80_48 gnd C_bl
Rb_80_49 bit_80_49 bit_80_50 R_bl
Rbb_80_49 bitb_80_49 bitb_80_50 R_bl
Cb_80_49 bit_80_49 gnd C_bl
Cbb_80_49 bitb_80_49 gnd C_bl
Rb_80_50 bit_80_50 bit_80_51 R_bl
Rbb_80_50 bitb_80_50 bitb_80_51 R_bl
Cb_80_50 bit_80_50 gnd C_bl
Cbb_80_50 bitb_80_50 gnd C_bl
Rb_80_51 bit_80_51 bit_80_52 R_bl
Rbb_80_51 bitb_80_51 bitb_80_52 R_bl
Cb_80_51 bit_80_51 gnd C_bl
Cbb_80_51 bitb_80_51 gnd C_bl
Rb_80_52 bit_80_52 bit_80_53 R_bl
Rbb_80_52 bitb_80_52 bitb_80_53 R_bl
Cb_80_52 bit_80_52 gnd C_bl
Cbb_80_52 bitb_80_52 gnd C_bl
Rb_80_53 bit_80_53 bit_80_54 R_bl
Rbb_80_53 bitb_80_53 bitb_80_54 R_bl
Cb_80_53 bit_80_53 gnd C_bl
Cbb_80_53 bitb_80_53 gnd C_bl
Rb_80_54 bit_80_54 bit_80_55 R_bl
Rbb_80_54 bitb_80_54 bitb_80_55 R_bl
Cb_80_54 bit_80_54 gnd C_bl
Cbb_80_54 bitb_80_54 gnd C_bl
Rb_80_55 bit_80_55 bit_80_56 R_bl
Rbb_80_55 bitb_80_55 bitb_80_56 R_bl
Cb_80_55 bit_80_55 gnd C_bl
Cbb_80_55 bitb_80_55 gnd C_bl
Rb_80_56 bit_80_56 bit_80_57 R_bl
Rbb_80_56 bitb_80_56 bitb_80_57 R_bl
Cb_80_56 bit_80_56 gnd C_bl
Cbb_80_56 bitb_80_56 gnd C_bl
Rb_80_57 bit_80_57 bit_80_58 R_bl
Rbb_80_57 bitb_80_57 bitb_80_58 R_bl
Cb_80_57 bit_80_57 gnd C_bl
Cbb_80_57 bitb_80_57 gnd C_bl
Rb_80_58 bit_80_58 bit_80_59 R_bl
Rbb_80_58 bitb_80_58 bitb_80_59 R_bl
Cb_80_58 bit_80_58 gnd C_bl
Cbb_80_58 bitb_80_58 gnd C_bl
Rb_80_59 bit_80_59 bit_80_60 R_bl
Rbb_80_59 bitb_80_59 bitb_80_60 R_bl
Cb_80_59 bit_80_59 gnd C_bl
Cbb_80_59 bitb_80_59 gnd C_bl
Rb_80_60 bit_80_60 bit_80_61 R_bl
Rbb_80_60 bitb_80_60 bitb_80_61 R_bl
Cb_80_60 bit_80_60 gnd C_bl
Cbb_80_60 bitb_80_60 gnd C_bl
Rb_80_61 bit_80_61 bit_80_62 R_bl
Rbb_80_61 bitb_80_61 bitb_80_62 R_bl
Cb_80_61 bit_80_61 gnd C_bl
Cbb_80_61 bitb_80_61 gnd C_bl
Rb_80_62 bit_80_62 bit_80_63 R_bl
Rbb_80_62 bitb_80_62 bitb_80_63 R_bl
Cb_80_62 bit_80_62 gnd C_bl
Cbb_80_62 bitb_80_62 gnd C_bl
Rb_80_63 bit_80_63 bit_80_64 R_bl
Rbb_80_63 bitb_80_63 bitb_80_64 R_bl
Cb_80_63 bit_80_63 gnd C_bl
Cbb_80_63 bitb_80_63 gnd C_bl
Rb_80_64 bit_80_64 bit_80_65 R_bl
Rbb_80_64 bitb_80_64 bitb_80_65 R_bl
Cb_80_64 bit_80_64 gnd C_bl
Cbb_80_64 bitb_80_64 gnd C_bl
Rb_80_65 bit_80_65 bit_80_66 R_bl
Rbb_80_65 bitb_80_65 bitb_80_66 R_bl
Cb_80_65 bit_80_65 gnd C_bl
Cbb_80_65 bitb_80_65 gnd C_bl
Rb_80_66 bit_80_66 bit_80_67 R_bl
Rbb_80_66 bitb_80_66 bitb_80_67 R_bl
Cb_80_66 bit_80_66 gnd C_bl
Cbb_80_66 bitb_80_66 gnd C_bl
Rb_80_67 bit_80_67 bit_80_68 R_bl
Rbb_80_67 bitb_80_67 bitb_80_68 R_bl
Cb_80_67 bit_80_67 gnd C_bl
Cbb_80_67 bitb_80_67 gnd C_bl
Rb_80_68 bit_80_68 bit_80_69 R_bl
Rbb_80_68 bitb_80_68 bitb_80_69 R_bl
Cb_80_68 bit_80_68 gnd C_bl
Cbb_80_68 bitb_80_68 gnd C_bl
Rb_80_69 bit_80_69 bit_80_70 R_bl
Rbb_80_69 bitb_80_69 bitb_80_70 R_bl
Cb_80_69 bit_80_69 gnd C_bl
Cbb_80_69 bitb_80_69 gnd C_bl
Rb_80_70 bit_80_70 bit_80_71 R_bl
Rbb_80_70 bitb_80_70 bitb_80_71 R_bl
Cb_80_70 bit_80_70 gnd C_bl
Cbb_80_70 bitb_80_70 gnd C_bl
Rb_80_71 bit_80_71 bit_80_72 R_bl
Rbb_80_71 bitb_80_71 bitb_80_72 R_bl
Cb_80_71 bit_80_71 gnd C_bl
Cbb_80_71 bitb_80_71 gnd C_bl
Rb_80_72 bit_80_72 bit_80_73 R_bl
Rbb_80_72 bitb_80_72 bitb_80_73 R_bl
Cb_80_72 bit_80_72 gnd C_bl
Cbb_80_72 bitb_80_72 gnd C_bl
Rb_80_73 bit_80_73 bit_80_74 R_bl
Rbb_80_73 bitb_80_73 bitb_80_74 R_bl
Cb_80_73 bit_80_73 gnd C_bl
Cbb_80_73 bitb_80_73 gnd C_bl
Rb_80_74 bit_80_74 bit_80_75 R_bl
Rbb_80_74 bitb_80_74 bitb_80_75 R_bl
Cb_80_74 bit_80_74 gnd C_bl
Cbb_80_74 bitb_80_74 gnd C_bl
Rb_80_75 bit_80_75 bit_80_76 R_bl
Rbb_80_75 bitb_80_75 bitb_80_76 R_bl
Cb_80_75 bit_80_75 gnd C_bl
Cbb_80_75 bitb_80_75 gnd C_bl
Rb_80_76 bit_80_76 bit_80_77 R_bl
Rbb_80_76 bitb_80_76 bitb_80_77 R_bl
Cb_80_76 bit_80_76 gnd C_bl
Cbb_80_76 bitb_80_76 gnd C_bl
Rb_80_77 bit_80_77 bit_80_78 R_bl
Rbb_80_77 bitb_80_77 bitb_80_78 R_bl
Cb_80_77 bit_80_77 gnd C_bl
Cbb_80_77 bitb_80_77 gnd C_bl
Rb_80_78 bit_80_78 bit_80_79 R_bl
Rbb_80_78 bitb_80_78 bitb_80_79 R_bl
Cb_80_78 bit_80_78 gnd C_bl
Cbb_80_78 bitb_80_78 gnd C_bl
Rb_80_79 bit_80_79 bit_80_80 R_bl
Rbb_80_79 bitb_80_79 bitb_80_80 R_bl
Cb_80_79 bit_80_79 gnd C_bl
Cbb_80_79 bitb_80_79 gnd C_bl
Rb_80_80 bit_80_80 bit_80_81 R_bl
Rbb_80_80 bitb_80_80 bitb_80_81 R_bl
Cb_80_80 bit_80_80 gnd C_bl
Cbb_80_80 bitb_80_80 gnd C_bl
Rb_80_81 bit_80_81 bit_80_82 R_bl
Rbb_80_81 bitb_80_81 bitb_80_82 R_bl
Cb_80_81 bit_80_81 gnd C_bl
Cbb_80_81 bitb_80_81 gnd C_bl
Rb_80_82 bit_80_82 bit_80_83 R_bl
Rbb_80_82 bitb_80_82 bitb_80_83 R_bl
Cb_80_82 bit_80_82 gnd C_bl
Cbb_80_82 bitb_80_82 gnd C_bl
Rb_80_83 bit_80_83 bit_80_84 R_bl
Rbb_80_83 bitb_80_83 bitb_80_84 R_bl
Cb_80_83 bit_80_83 gnd C_bl
Cbb_80_83 bitb_80_83 gnd C_bl
Rb_80_84 bit_80_84 bit_80_85 R_bl
Rbb_80_84 bitb_80_84 bitb_80_85 R_bl
Cb_80_84 bit_80_84 gnd C_bl
Cbb_80_84 bitb_80_84 gnd C_bl
Rb_80_85 bit_80_85 bit_80_86 R_bl
Rbb_80_85 bitb_80_85 bitb_80_86 R_bl
Cb_80_85 bit_80_85 gnd C_bl
Cbb_80_85 bitb_80_85 gnd C_bl
Rb_80_86 bit_80_86 bit_80_87 R_bl
Rbb_80_86 bitb_80_86 bitb_80_87 R_bl
Cb_80_86 bit_80_86 gnd C_bl
Cbb_80_86 bitb_80_86 gnd C_bl
Rb_80_87 bit_80_87 bit_80_88 R_bl
Rbb_80_87 bitb_80_87 bitb_80_88 R_bl
Cb_80_87 bit_80_87 gnd C_bl
Cbb_80_87 bitb_80_87 gnd C_bl
Rb_80_88 bit_80_88 bit_80_89 R_bl
Rbb_80_88 bitb_80_88 bitb_80_89 R_bl
Cb_80_88 bit_80_88 gnd C_bl
Cbb_80_88 bitb_80_88 gnd C_bl
Rb_80_89 bit_80_89 bit_80_90 R_bl
Rbb_80_89 bitb_80_89 bitb_80_90 R_bl
Cb_80_89 bit_80_89 gnd C_bl
Cbb_80_89 bitb_80_89 gnd C_bl
Rb_80_90 bit_80_90 bit_80_91 R_bl
Rbb_80_90 bitb_80_90 bitb_80_91 R_bl
Cb_80_90 bit_80_90 gnd C_bl
Cbb_80_90 bitb_80_90 gnd C_bl
Rb_80_91 bit_80_91 bit_80_92 R_bl
Rbb_80_91 bitb_80_91 bitb_80_92 R_bl
Cb_80_91 bit_80_91 gnd C_bl
Cbb_80_91 bitb_80_91 gnd C_bl
Rb_80_92 bit_80_92 bit_80_93 R_bl
Rbb_80_92 bitb_80_92 bitb_80_93 R_bl
Cb_80_92 bit_80_92 gnd C_bl
Cbb_80_92 bitb_80_92 gnd C_bl
Rb_80_93 bit_80_93 bit_80_94 R_bl
Rbb_80_93 bitb_80_93 bitb_80_94 R_bl
Cb_80_93 bit_80_93 gnd C_bl
Cbb_80_93 bitb_80_93 gnd C_bl
Rb_80_94 bit_80_94 bit_80_95 R_bl
Rbb_80_94 bitb_80_94 bitb_80_95 R_bl
Cb_80_94 bit_80_94 gnd C_bl
Cbb_80_94 bitb_80_94 gnd C_bl
Rb_80_95 bit_80_95 bit_80_96 R_bl
Rbb_80_95 bitb_80_95 bitb_80_96 R_bl
Cb_80_95 bit_80_95 gnd C_bl
Cbb_80_95 bitb_80_95 gnd C_bl
Rb_80_96 bit_80_96 bit_80_97 R_bl
Rbb_80_96 bitb_80_96 bitb_80_97 R_bl
Cb_80_96 bit_80_96 gnd C_bl
Cbb_80_96 bitb_80_96 gnd C_bl
Rb_80_97 bit_80_97 bit_80_98 R_bl
Rbb_80_97 bitb_80_97 bitb_80_98 R_bl
Cb_80_97 bit_80_97 gnd C_bl
Cbb_80_97 bitb_80_97 gnd C_bl
Rb_80_98 bit_80_98 bit_80_99 R_bl
Rbb_80_98 bitb_80_98 bitb_80_99 R_bl
Cb_80_98 bit_80_98 gnd C_bl
Cbb_80_98 bitb_80_98 gnd C_bl
Rb_80_99 bit_80_99 bit_80_100 R_bl
Rbb_80_99 bitb_80_99 bitb_80_100 R_bl
Cb_80_99 bit_80_99 gnd C_bl
Cbb_80_99 bitb_80_99 gnd C_bl
Rb_81_0 bit_81_0 bit_81_1 R_bl
Rbb_81_0 bitb_81_0 bitb_81_1 R_bl
Cb_81_0 bit_81_0 gnd C_bl
Cbb_81_0 bitb_81_0 gnd C_bl
Rb_81_1 bit_81_1 bit_81_2 R_bl
Rbb_81_1 bitb_81_1 bitb_81_2 R_bl
Cb_81_1 bit_81_1 gnd C_bl
Cbb_81_1 bitb_81_1 gnd C_bl
Rb_81_2 bit_81_2 bit_81_3 R_bl
Rbb_81_2 bitb_81_2 bitb_81_3 R_bl
Cb_81_2 bit_81_2 gnd C_bl
Cbb_81_2 bitb_81_2 gnd C_bl
Rb_81_3 bit_81_3 bit_81_4 R_bl
Rbb_81_3 bitb_81_3 bitb_81_4 R_bl
Cb_81_3 bit_81_3 gnd C_bl
Cbb_81_3 bitb_81_3 gnd C_bl
Rb_81_4 bit_81_4 bit_81_5 R_bl
Rbb_81_4 bitb_81_4 bitb_81_5 R_bl
Cb_81_4 bit_81_4 gnd C_bl
Cbb_81_4 bitb_81_4 gnd C_bl
Rb_81_5 bit_81_5 bit_81_6 R_bl
Rbb_81_5 bitb_81_5 bitb_81_6 R_bl
Cb_81_5 bit_81_5 gnd C_bl
Cbb_81_5 bitb_81_5 gnd C_bl
Rb_81_6 bit_81_6 bit_81_7 R_bl
Rbb_81_6 bitb_81_6 bitb_81_7 R_bl
Cb_81_6 bit_81_6 gnd C_bl
Cbb_81_6 bitb_81_6 gnd C_bl
Rb_81_7 bit_81_7 bit_81_8 R_bl
Rbb_81_7 bitb_81_7 bitb_81_8 R_bl
Cb_81_7 bit_81_7 gnd C_bl
Cbb_81_7 bitb_81_7 gnd C_bl
Rb_81_8 bit_81_8 bit_81_9 R_bl
Rbb_81_8 bitb_81_8 bitb_81_9 R_bl
Cb_81_8 bit_81_8 gnd C_bl
Cbb_81_8 bitb_81_8 gnd C_bl
Rb_81_9 bit_81_9 bit_81_10 R_bl
Rbb_81_9 bitb_81_9 bitb_81_10 R_bl
Cb_81_9 bit_81_9 gnd C_bl
Cbb_81_9 bitb_81_9 gnd C_bl
Rb_81_10 bit_81_10 bit_81_11 R_bl
Rbb_81_10 bitb_81_10 bitb_81_11 R_bl
Cb_81_10 bit_81_10 gnd C_bl
Cbb_81_10 bitb_81_10 gnd C_bl
Rb_81_11 bit_81_11 bit_81_12 R_bl
Rbb_81_11 bitb_81_11 bitb_81_12 R_bl
Cb_81_11 bit_81_11 gnd C_bl
Cbb_81_11 bitb_81_11 gnd C_bl
Rb_81_12 bit_81_12 bit_81_13 R_bl
Rbb_81_12 bitb_81_12 bitb_81_13 R_bl
Cb_81_12 bit_81_12 gnd C_bl
Cbb_81_12 bitb_81_12 gnd C_bl
Rb_81_13 bit_81_13 bit_81_14 R_bl
Rbb_81_13 bitb_81_13 bitb_81_14 R_bl
Cb_81_13 bit_81_13 gnd C_bl
Cbb_81_13 bitb_81_13 gnd C_bl
Rb_81_14 bit_81_14 bit_81_15 R_bl
Rbb_81_14 bitb_81_14 bitb_81_15 R_bl
Cb_81_14 bit_81_14 gnd C_bl
Cbb_81_14 bitb_81_14 gnd C_bl
Rb_81_15 bit_81_15 bit_81_16 R_bl
Rbb_81_15 bitb_81_15 bitb_81_16 R_bl
Cb_81_15 bit_81_15 gnd C_bl
Cbb_81_15 bitb_81_15 gnd C_bl
Rb_81_16 bit_81_16 bit_81_17 R_bl
Rbb_81_16 bitb_81_16 bitb_81_17 R_bl
Cb_81_16 bit_81_16 gnd C_bl
Cbb_81_16 bitb_81_16 gnd C_bl
Rb_81_17 bit_81_17 bit_81_18 R_bl
Rbb_81_17 bitb_81_17 bitb_81_18 R_bl
Cb_81_17 bit_81_17 gnd C_bl
Cbb_81_17 bitb_81_17 gnd C_bl
Rb_81_18 bit_81_18 bit_81_19 R_bl
Rbb_81_18 bitb_81_18 bitb_81_19 R_bl
Cb_81_18 bit_81_18 gnd C_bl
Cbb_81_18 bitb_81_18 gnd C_bl
Rb_81_19 bit_81_19 bit_81_20 R_bl
Rbb_81_19 bitb_81_19 bitb_81_20 R_bl
Cb_81_19 bit_81_19 gnd C_bl
Cbb_81_19 bitb_81_19 gnd C_bl
Rb_81_20 bit_81_20 bit_81_21 R_bl
Rbb_81_20 bitb_81_20 bitb_81_21 R_bl
Cb_81_20 bit_81_20 gnd C_bl
Cbb_81_20 bitb_81_20 gnd C_bl
Rb_81_21 bit_81_21 bit_81_22 R_bl
Rbb_81_21 bitb_81_21 bitb_81_22 R_bl
Cb_81_21 bit_81_21 gnd C_bl
Cbb_81_21 bitb_81_21 gnd C_bl
Rb_81_22 bit_81_22 bit_81_23 R_bl
Rbb_81_22 bitb_81_22 bitb_81_23 R_bl
Cb_81_22 bit_81_22 gnd C_bl
Cbb_81_22 bitb_81_22 gnd C_bl
Rb_81_23 bit_81_23 bit_81_24 R_bl
Rbb_81_23 bitb_81_23 bitb_81_24 R_bl
Cb_81_23 bit_81_23 gnd C_bl
Cbb_81_23 bitb_81_23 gnd C_bl
Rb_81_24 bit_81_24 bit_81_25 R_bl
Rbb_81_24 bitb_81_24 bitb_81_25 R_bl
Cb_81_24 bit_81_24 gnd C_bl
Cbb_81_24 bitb_81_24 gnd C_bl
Rb_81_25 bit_81_25 bit_81_26 R_bl
Rbb_81_25 bitb_81_25 bitb_81_26 R_bl
Cb_81_25 bit_81_25 gnd C_bl
Cbb_81_25 bitb_81_25 gnd C_bl
Rb_81_26 bit_81_26 bit_81_27 R_bl
Rbb_81_26 bitb_81_26 bitb_81_27 R_bl
Cb_81_26 bit_81_26 gnd C_bl
Cbb_81_26 bitb_81_26 gnd C_bl
Rb_81_27 bit_81_27 bit_81_28 R_bl
Rbb_81_27 bitb_81_27 bitb_81_28 R_bl
Cb_81_27 bit_81_27 gnd C_bl
Cbb_81_27 bitb_81_27 gnd C_bl
Rb_81_28 bit_81_28 bit_81_29 R_bl
Rbb_81_28 bitb_81_28 bitb_81_29 R_bl
Cb_81_28 bit_81_28 gnd C_bl
Cbb_81_28 bitb_81_28 gnd C_bl
Rb_81_29 bit_81_29 bit_81_30 R_bl
Rbb_81_29 bitb_81_29 bitb_81_30 R_bl
Cb_81_29 bit_81_29 gnd C_bl
Cbb_81_29 bitb_81_29 gnd C_bl
Rb_81_30 bit_81_30 bit_81_31 R_bl
Rbb_81_30 bitb_81_30 bitb_81_31 R_bl
Cb_81_30 bit_81_30 gnd C_bl
Cbb_81_30 bitb_81_30 gnd C_bl
Rb_81_31 bit_81_31 bit_81_32 R_bl
Rbb_81_31 bitb_81_31 bitb_81_32 R_bl
Cb_81_31 bit_81_31 gnd C_bl
Cbb_81_31 bitb_81_31 gnd C_bl
Rb_81_32 bit_81_32 bit_81_33 R_bl
Rbb_81_32 bitb_81_32 bitb_81_33 R_bl
Cb_81_32 bit_81_32 gnd C_bl
Cbb_81_32 bitb_81_32 gnd C_bl
Rb_81_33 bit_81_33 bit_81_34 R_bl
Rbb_81_33 bitb_81_33 bitb_81_34 R_bl
Cb_81_33 bit_81_33 gnd C_bl
Cbb_81_33 bitb_81_33 gnd C_bl
Rb_81_34 bit_81_34 bit_81_35 R_bl
Rbb_81_34 bitb_81_34 bitb_81_35 R_bl
Cb_81_34 bit_81_34 gnd C_bl
Cbb_81_34 bitb_81_34 gnd C_bl
Rb_81_35 bit_81_35 bit_81_36 R_bl
Rbb_81_35 bitb_81_35 bitb_81_36 R_bl
Cb_81_35 bit_81_35 gnd C_bl
Cbb_81_35 bitb_81_35 gnd C_bl
Rb_81_36 bit_81_36 bit_81_37 R_bl
Rbb_81_36 bitb_81_36 bitb_81_37 R_bl
Cb_81_36 bit_81_36 gnd C_bl
Cbb_81_36 bitb_81_36 gnd C_bl
Rb_81_37 bit_81_37 bit_81_38 R_bl
Rbb_81_37 bitb_81_37 bitb_81_38 R_bl
Cb_81_37 bit_81_37 gnd C_bl
Cbb_81_37 bitb_81_37 gnd C_bl
Rb_81_38 bit_81_38 bit_81_39 R_bl
Rbb_81_38 bitb_81_38 bitb_81_39 R_bl
Cb_81_38 bit_81_38 gnd C_bl
Cbb_81_38 bitb_81_38 gnd C_bl
Rb_81_39 bit_81_39 bit_81_40 R_bl
Rbb_81_39 bitb_81_39 bitb_81_40 R_bl
Cb_81_39 bit_81_39 gnd C_bl
Cbb_81_39 bitb_81_39 gnd C_bl
Rb_81_40 bit_81_40 bit_81_41 R_bl
Rbb_81_40 bitb_81_40 bitb_81_41 R_bl
Cb_81_40 bit_81_40 gnd C_bl
Cbb_81_40 bitb_81_40 gnd C_bl
Rb_81_41 bit_81_41 bit_81_42 R_bl
Rbb_81_41 bitb_81_41 bitb_81_42 R_bl
Cb_81_41 bit_81_41 gnd C_bl
Cbb_81_41 bitb_81_41 gnd C_bl
Rb_81_42 bit_81_42 bit_81_43 R_bl
Rbb_81_42 bitb_81_42 bitb_81_43 R_bl
Cb_81_42 bit_81_42 gnd C_bl
Cbb_81_42 bitb_81_42 gnd C_bl
Rb_81_43 bit_81_43 bit_81_44 R_bl
Rbb_81_43 bitb_81_43 bitb_81_44 R_bl
Cb_81_43 bit_81_43 gnd C_bl
Cbb_81_43 bitb_81_43 gnd C_bl
Rb_81_44 bit_81_44 bit_81_45 R_bl
Rbb_81_44 bitb_81_44 bitb_81_45 R_bl
Cb_81_44 bit_81_44 gnd C_bl
Cbb_81_44 bitb_81_44 gnd C_bl
Rb_81_45 bit_81_45 bit_81_46 R_bl
Rbb_81_45 bitb_81_45 bitb_81_46 R_bl
Cb_81_45 bit_81_45 gnd C_bl
Cbb_81_45 bitb_81_45 gnd C_bl
Rb_81_46 bit_81_46 bit_81_47 R_bl
Rbb_81_46 bitb_81_46 bitb_81_47 R_bl
Cb_81_46 bit_81_46 gnd C_bl
Cbb_81_46 bitb_81_46 gnd C_bl
Rb_81_47 bit_81_47 bit_81_48 R_bl
Rbb_81_47 bitb_81_47 bitb_81_48 R_bl
Cb_81_47 bit_81_47 gnd C_bl
Cbb_81_47 bitb_81_47 gnd C_bl
Rb_81_48 bit_81_48 bit_81_49 R_bl
Rbb_81_48 bitb_81_48 bitb_81_49 R_bl
Cb_81_48 bit_81_48 gnd C_bl
Cbb_81_48 bitb_81_48 gnd C_bl
Rb_81_49 bit_81_49 bit_81_50 R_bl
Rbb_81_49 bitb_81_49 bitb_81_50 R_bl
Cb_81_49 bit_81_49 gnd C_bl
Cbb_81_49 bitb_81_49 gnd C_bl
Rb_81_50 bit_81_50 bit_81_51 R_bl
Rbb_81_50 bitb_81_50 bitb_81_51 R_bl
Cb_81_50 bit_81_50 gnd C_bl
Cbb_81_50 bitb_81_50 gnd C_bl
Rb_81_51 bit_81_51 bit_81_52 R_bl
Rbb_81_51 bitb_81_51 bitb_81_52 R_bl
Cb_81_51 bit_81_51 gnd C_bl
Cbb_81_51 bitb_81_51 gnd C_bl
Rb_81_52 bit_81_52 bit_81_53 R_bl
Rbb_81_52 bitb_81_52 bitb_81_53 R_bl
Cb_81_52 bit_81_52 gnd C_bl
Cbb_81_52 bitb_81_52 gnd C_bl
Rb_81_53 bit_81_53 bit_81_54 R_bl
Rbb_81_53 bitb_81_53 bitb_81_54 R_bl
Cb_81_53 bit_81_53 gnd C_bl
Cbb_81_53 bitb_81_53 gnd C_bl
Rb_81_54 bit_81_54 bit_81_55 R_bl
Rbb_81_54 bitb_81_54 bitb_81_55 R_bl
Cb_81_54 bit_81_54 gnd C_bl
Cbb_81_54 bitb_81_54 gnd C_bl
Rb_81_55 bit_81_55 bit_81_56 R_bl
Rbb_81_55 bitb_81_55 bitb_81_56 R_bl
Cb_81_55 bit_81_55 gnd C_bl
Cbb_81_55 bitb_81_55 gnd C_bl
Rb_81_56 bit_81_56 bit_81_57 R_bl
Rbb_81_56 bitb_81_56 bitb_81_57 R_bl
Cb_81_56 bit_81_56 gnd C_bl
Cbb_81_56 bitb_81_56 gnd C_bl
Rb_81_57 bit_81_57 bit_81_58 R_bl
Rbb_81_57 bitb_81_57 bitb_81_58 R_bl
Cb_81_57 bit_81_57 gnd C_bl
Cbb_81_57 bitb_81_57 gnd C_bl
Rb_81_58 bit_81_58 bit_81_59 R_bl
Rbb_81_58 bitb_81_58 bitb_81_59 R_bl
Cb_81_58 bit_81_58 gnd C_bl
Cbb_81_58 bitb_81_58 gnd C_bl
Rb_81_59 bit_81_59 bit_81_60 R_bl
Rbb_81_59 bitb_81_59 bitb_81_60 R_bl
Cb_81_59 bit_81_59 gnd C_bl
Cbb_81_59 bitb_81_59 gnd C_bl
Rb_81_60 bit_81_60 bit_81_61 R_bl
Rbb_81_60 bitb_81_60 bitb_81_61 R_bl
Cb_81_60 bit_81_60 gnd C_bl
Cbb_81_60 bitb_81_60 gnd C_bl
Rb_81_61 bit_81_61 bit_81_62 R_bl
Rbb_81_61 bitb_81_61 bitb_81_62 R_bl
Cb_81_61 bit_81_61 gnd C_bl
Cbb_81_61 bitb_81_61 gnd C_bl
Rb_81_62 bit_81_62 bit_81_63 R_bl
Rbb_81_62 bitb_81_62 bitb_81_63 R_bl
Cb_81_62 bit_81_62 gnd C_bl
Cbb_81_62 bitb_81_62 gnd C_bl
Rb_81_63 bit_81_63 bit_81_64 R_bl
Rbb_81_63 bitb_81_63 bitb_81_64 R_bl
Cb_81_63 bit_81_63 gnd C_bl
Cbb_81_63 bitb_81_63 gnd C_bl
Rb_81_64 bit_81_64 bit_81_65 R_bl
Rbb_81_64 bitb_81_64 bitb_81_65 R_bl
Cb_81_64 bit_81_64 gnd C_bl
Cbb_81_64 bitb_81_64 gnd C_bl
Rb_81_65 bit_81_65 bit_81_66 R_bl
Rbb_81_65 bitb_81_65 bitb_81_66 R_bl
Cb_81_65 bit_81_65 gnd C_bl
Cbb_81_65 bitb_81_65 gnd C_bl
Rb_81_66 bit_81_66 bit_81_67 R_bl
Rbb_81_66 bitb_81_66 bitb_81_67 R_bl
Cb_81_66 bit_81_66 gnd C_bl
Cbb_81_66 bitb_81_66 gnd C_bl
Rb_81_67 bit_81_67 bit_81_68 R_bl
Rbb_81_67 bitb_81_67 bitb_81_68 R_bl
Cb_81_67 bit_81_67 gnd C_bl
Cbb_81_67 bitb_81_67 gnd C_bl
Rb_81_68 bit_81_68 bit_81_69 R_bl
Rbb_81_68 bitb_81_68 bitb_81_69 R_bl
Cb_81_68 bit_81_68 gnd C_bl
Cbb_81_68 bitb_81_68 gnd C_bl
Rb_81_69 bit_81_69 bit_81_70 R_bl
Rbb_81_69 bitb_81_69 bitb_81_70 R_bl
Cb_81_69 bit_81_69 gnd C_bl
Cbb_81_69 bitb_81_69 gnd C_bl
Rb_81_70 bit_81_70 bit_81_71 R_bl
Rbb_81_70 bitb_81_70 bitb_81_71 R_bl
Cb_81_70 bit_81_70 gnd C_bl
Cbb_81_70 bitb_81_70 gnd C_bl
Rb_81_71 bit_81_71 bit_81_72 R_bl
Rbb_81_71 bitb_81_71 bitb_81_72 R_bl
Cb_81_71 bit_81_71 gnd C_bl
Cbb_81_71 bitb_81_71 gnd C_bl
Rb_81_72 bit_81_72 bit_81_73 R_bl
Rbb_81_72 bitb_81_72 bitb_81_73 R_bl
Cb_81_72 bit_81_72 gnd C_bl
Cbb_81_72 bitb_81_72 gnd C_bl
Rb_81_73 bit_81_73 bit_81_74 R_bl
Rbb_81_73 bitb_81_73 bitb_81_74 R_bl
Cb_81_73 bit_81_73 gnd C_bl
Cbb_81_73 bitb_81_73 gnd C_bl
Rb_81_74 bit_81_74 bit_81_75 R_bl
Rbb_81_74 bitb_81_74 bitb_81_75 R_bl
Cb_81_74 bit_81_74 gnd C_bl
Cbb_81_74 bitb_81_74 gnd C_bl
Rb_81_75 bit_81_75 bit_81_76 R_bl
Rbb_81_75 bitb_81_75 bitb_81_76 R_bl
Cb_81_75 bit_81_75 gnd C_bl
Cbb_81_75 bitb_81_75 gnd C_bl
Rb_81_76 bit_81_76 bit_81_77 R_bl
Rbb_81_76 bitb_81_76 bitb_81_77 R_bl
Cb_81_76 bit_81_76 gnd C_bl
Cbb_81_76 bitb_81_76 gnd C_bl
Rb_81_77 bit_81_77 bit_81_78 R_bl
Rbb_81_77 bitb_81_77 bitb_81_78 R_bl
Cb_81_77 bit_81_77 gnd C_bl
Cbb_81_77 bitb_81_77 gnd C_bl
Rb_81_78 bit_81_78 bit_81_79 R_bl
Rbb_81_78 bitb_81_78 bitb_81_79 R_bl
Cb_81_78 bit_81_78 gnd C_bl
Cbb_81_78 bitb_81_78 gnd C_bl
Rb_81_79 bit_81_79 bit_81_80 R_bl
Rbb_81_79 bitb_81_79 bitb_81_80 R_bl
Cb_81_79 bit_81_79 gnd C_bl
Cbb_81_79 bitb_81_79 gnd C_bl
Rb_81_80 bit_81_80 bit_81_81 R_bl
Rbb_81_80 bitb_81_80 bitb_81_81 R_bl
Cb_81_80 bit_81_80 gnd C_bl
Cbb_81_80 bitb_81_80 gnd C_bl
Rb_81_81 bit_81_81 bit_81_82 R_bl
Rbb_81_81 bitb_81_81 bitb_81_82 R_bl
Cb_81_81 bit_81_81 gnd C_bl
Cbb_81_81 bitb_81_81 gnd C_bl
Rb_81_82 bit_81_82 bit_81_83 R_bl
Rbb_81_82 bitb_81_82 bitb_81_83 R_bl
Cb_81_82 bit_81_82 gnd C_bl
Cbb_81_82 bitb_81_82 gnd C_bl
Rb_81_83 bit_81_83 bit_81_84 R_bl
Rbb_81_83 bitb_81_83 bitb_81_84 R_bl
Cb_81_83 bit_81_83 gnd C_bl
Cbb_81_83 bitb_81_83 gnd C_bl
Rb_81_84 bit_81_84 bit_81_85 R_bl
Rbb_81_84 bitb_81_84 bitb_81_85 R_bl
Cb_81_84 bit_81_84 gnd C_bl
Cbb_81_84 bitb_81_84 gnd C_bl
Rb_81_85 bit_81_85 bit_81_86 R_bl
Rbb_81_85 bitb_81_85 bitb_81_86 R_bl
Cb_81_85 bit_81_85 gnd C_bl
Cbb_81_85 bitb_81_85 gnd C_bl
Rb_81_86 bit_81_86 bit_81_87 R_bl
Rbb_81_86 bitb_81_86 bitb_81_87 R_bl
Cb_81_86 bit_81_86 gnd C_bl
Cbb_81_86 bitb_81_86 gnd C_bl
Rb_81_87 bit_81_87 bit_81_88 R_bl
Rbb_81_87 bitb_81_87 bitb_81_88 R_bl
Cb_81_87 bit_81_87 gnd C_bl
Cbb_81_87 bitb_81_87 gnd C_bl
Rb_81_88 bit_81_88 bit_81_89 R_bl
Rbb_81_88 bitb_81_88 bitb_81_89 R_bl
Cb_81_88 bit_81_88 gnd C_bl
Cbb_81_88 bitb_81_88 gnd C_bl
Rb_81_89 bit_81_89 bit_81_90 R_bl
Rbb_81_89 bitb_81_89 bitb_81_90 R_bl
Cb_81_89 bit_81_89 gnd C_bl
Cbb_81_89 bitb_81_89 gnd C_bl
Rb_81_90 bit_81_90 bit_81_91 R_bl
Rbb_81_90 bitb_81_90 bitb_81_91 R_bl
Cb_81_90 bit_81_90 gnd C_bl
Cbb_81_90 bitb_81_90 gnd C_bl
Rb_81_91 bit_81_91 bit_81_92 R_bl
Rbb_81_91 bitb_81_91 bitb_81_92 R_bl
Cb_81_91 bit_81_91 gnd C_bl
Cbb_81_91 bitb_81_91 gnd C_bl
Rb_81_92 bit_81_92 bit_81_93 R_bl
Rbb_81_92 bitb_81_92 bitb_81_93 R_bl
Cb_81_92 bit_81_92 gnd C_bl
Cbb_81_92 bitb_81_92 gnd C_bl
Rb_81_93 bit_81_93 bit_81_94 R_bl
Rbb_81_93 bitb_81_93 bitb_81_94 R_bl
Cb_81_93 bit_81_93 gnd C_bl
Cbb_81_93 bitb_81_93 gnd C_bl
Rb_81_94 bit_81_94 bit_81_95 R_bl
Rbb_81_94 bitb_81_94 bitb_81_95 R_bl
Cb_81_94 bit_81_94 gnd C_bl
Cbb_81_94 bitb_81_94 gnd C_bl
Rb_81_95 bit_81_95 bit_81_96 R_bl
Rbb_81_95 bitb_81_95 bitb_81_96 R_bl
Cb_81_95 bit_81_95 gnd C_bl
Cbb_81_95 bitb_81_95 gnd C_bl
Rb_81_96 bit_81_96 bit_81_97 R_bl
Rbb_81_96 bitb_81_96 bitb_81_97 R_bl
Cb_81_96 bit_81_96 gnd C_bl
Cbb_81_96 bitb_81_96 gnd C_bl
Rb_81_97 bit_81_97 bit_81_98 R_bl
Rbb_81_97 bitb_81_97 bitb_81_98 R_bl
Cb_81_97 bit_81_97 gnd C_bl
Cbb_81_97 bitb_81_97 gnd C_bl
Rb_81_98 bit_81_98 bit_81_99 R_bl
Rbb_81_98 bitb_81_98 bitb_81_99 R_bl
Cb_81_98 bit_81_98 gnd C_bl
Cbb_81_98 bitb_81_98 gnd C_bl
Rb_81_99 bit_81_99 bit_81_100 R_bl
Rbb_81_99 bitb_81_99 bitb_81_100 R_bl
Cb_81_99 bit_81_99 gnd C_bl
Cbb_81_99 bitb_81_99 gnd C_bl
Rb_82_0 bit_82_0 bit_82_1 R_bl
Rbb_82_0 bitb_82_0 bitb_82_1 R_bl
Cb_82_0 bit_82_0 gnd C_bl
Cbb_82_0 bitb_82_0 gnd C_bl
Rb_82_1 bit_82_1 bit_82_2 R_bl
Rbb_82_1 bitb_82_1 bitb_82_2 R_bl
Cb_82_1 bit_82_1 gnd C_bl
Cbb_82_1 bitb_82_1 gnd C_bl
Rb_82_2 bit_82_2 bit_82_3 R_bl
Rbb_82_2 bitb_82_2 bitb_82_3 R_bl
Cb_82_2 bit_82_2 gnd C_bl
Cbb_82_2 bitb_82_2 gnd C_bl
Rb_82_3 bit_82_3 bit_82_4 R_bl
Rbb_82_3 bitb_82_3 bitb_82_4 R_bl
Cb_82_3 bit_82_3 gnd C_bl
Cbb_82_3 bitb_82_3 gnd C_bl
Rb_82_4 bit_82_4 bit_82_5 R_bl
Rbb_82_4 bitb_82_4 bitb_82_5 R_bl
Cb_82_4 bit_82_4 gnd C_bl
Cbb_82_4 bitb_82_4 gnd C_bl
Rb_82_5 bit_82_5 bit_82_6 R_bl
Rbb_82_5 bitb_82_5 bitb_82_6 R_bl
Cb_82_5 bit_82_5 gnd C_bl
Cbb_82_5 bitb_82_5 gnd C_bl
Rb_82_6 bit_82_6 bit_82_7 R_bl
Rbb_82_6 bitb_82_6 bitb_82_7 R_bl
Cb_82_6 bit_82_6 gnd C_bl
Cbb_82_6 bitb_82_6 gnd C_bl
Rb_82_7 bit_82_7 bit_82_8 R_bl
Rbb_82_7 bitb_82_7 bitb_82_8 R_bl
Cb_82_7 bit_82_7 gnd C_bl
Cbb_82_7 bitb_82_7 gnd C_bl
Rb_82_8 bit_82_8 bit_82_9 R_bl
Rbb_82_8 bitb_82_8 bitb_82_9 R_bl
Cb_82_8 bit_82_8 gnd C_bl
Cbb_82_8 bitb_82_8 gnd C_bl
Rb_82_9 bit_82_9 bit_82_10 R_bl
Rbb_82_9 bitb_82_9 bitb_82_10 R_bl
Cb_82_9 bit_82_9 gnd C_bl
Cbb_82_9 bitb_82_9 gnd C_bl
Rb_82_10 bit_82_10 bit_82_11 R_bl
Rbb_82_10 bitb_82_10 bitb_82_11 R_bl
Cb_82_10 bit_82_10 gnd C_bl
Cbb_82_10 bitb_82_10 gnd C_bl
Rb_82_11 bit_82_11 bit_82_12 R_bl
Rbb_82_11 bitb_82_11 bitb_82_12 R_bl
Cb_82_11 bit_82_11 gnd C_bl
Cbb_82_11 bitb_82_11 gnd C_bl
Rb_82_12 bit_82_12 bit_82_13 R_bl
Rbb_82_12 bitb_82_12 bitb_82_13 R_bl
Cb_82_12 bit_82_12 gnd C_bl
Cbb_82_12 bitb_82_12 gnd C_bl
Rb_82_13 bit_82_13 bit_82_14 R_bl
Rbb_82_13 bitb_82_13 bitb_82_14 R_bl
Cb_82_13 bit_82_13 gnd C_bl
Cbb_82_13 bitb_82_13 gnd C_bl
Rb_82_14 bit_82_14 bit_82_15 R_bl
Rbb_82_14 bitb_82_14 bitb_82_15 R_bl
Cb_82_14 bit_82_14 gnd C_bl
Cbb_82_14 bitb_82_14 gnd C_bl
Rb_82_15 bit_82_15 bit_82_16 R_bl
Rbb_82_15 bitb_82_15 bitb_82_16 R_bl
Cb_82_15 bit_82_15 gnd C_bl
Cbb_82_15 bitb_82_15 gnd C_bl
Rb_82_16 bit_82_16 bit_82_17 R_bl
Rbb_82_16 bitb_82_16 bitb_82_17 R_bl
Cb_82_16 bit_82_16 gnd C_bl
Cbb_82_16 bitb_82_16 gnd C_bl
Rb_82_17 bit_82_17 bit_82_18 R_bl
Rbb_82_17 bitb_82_17 bitb_82_18 R_bl
Cb_82_17 bit_82_17 gnd C_bl
Cbb_82_17 bitb_82_17 gnd C_bl
Rb_82_18 bit_82_18 bit_82_19 R_bl
Rbb_82_18 bitb_82_18 bitb_82_19 R_bl
Cb_82_18 bit_82_18 gnd C_bl
Cbb_82_18 bitb_82_18 gnd C_bl
Rb_82_19 bit_82_19 bit_82_20 R_bl
Rbb_82_19 bitb_82_19 bitb_82_20 R_bl
Cb_82_19 bit_82_19 gnd C_bl
Cbb_82_19 bitb_82_19 gnd C_bl
Rb_82_20 bit_82_20 bit_82_21 R_bl
Rbb_82_20 bitb_82_20 bitb_82_21 R_bl
Cb_82_20 bit_82_20 gnd C_bl
Cbb_82_20 bitb_82_20 gnd C_bl
Rb_82_21 bit_82_21 bit_82_22 R_bl
Rbb_82_21 bitb_82_21 bitb_82_22 R_bl
Cb_82_21 bit_82_21 gnd C_bl
Cbb_82_21 bitb_82_21 gnd C_bl
Rb_82_22 bit_82_22 bit_82_23 R_bl
Rbb_82_22 bitb_82_22 bitb_82_23 R_bl
Cb_82_22 bit_82_22 gnd C_bl
Cbb_82_22 bitb_82_22 gnd C_bl
Rb_82_23 bit_82_23 bit_82_24 R_bl
Rbb_82_23 bitb_82_23 bitb_82_24 R_bl
Cb_82_23 bit_82_23 gnd C_bl
Cbb_82_23 bitb_82_23 gnd C_bl
Rb_82_24 bit_82_24 bit_82_25 R_bl
Rbb_82_24 bitb_82_24 bitb_82_25 R_bl
Cb_82_24 bit_82_24 gnd C_bl
Cbb_82_24 bitb_82_24 gnd C_bl
Rb_82_25 bit_82_25 bit_82_26 R_bl
Rbb_82_25 bitb_82_25 bitb_82_26 R_bl
Cb_82_25 bit_82_25 gnd C_bl
Cbb_82_25 bitb_82_25 gnd C_bl
Rb_82_26 bit_82_26 bit_82_27 R_bl
Rbb_82_26 bitb_82_26 bitb_82_27 R_bl
Cb_82_26 bit_82_26 gnd C_bl
Cbb_82_26 bitb_82_26 gnd C_bl
Rb_82_27 bit_82_27 bit_82_28 R_bl
Rbb_82_27 bitb_82_27 bitb_82_28 R_bl
Cb_82_27 bit_82_27 gnd C_bl
Cbb_82_27 bitb_82_27 gnd C_bl
Rb_82_28 bit_82_28 bit_82_29 R_bl
Rbb_82_28 bitb_82_28 bitb_82_29 R_bl
Cb_82_28 bit_82_28 gnd C_bl
Cbb_82_28 bitb_82_28 gnd C_bl
Rb_82_29 bit_82_29 bit_82_30 R_bl
Rbb_82_29 bitb_82_29 bitb_82_30 R_bl
Cb_82_29 bit_82_29 gnd C_bl
Cbb_82_29 bitb_82_29 gnd C_bl
Rb_82_30 bit_82_30 bit_82_31 R_bl
Rbb_82_30 bitb_82_30 bitb_82_31 R_bl
Cb_82_30 bit_82_30 gnd C_bl
Cbb_82_30 bitb_82_30 gnd C_bl
Rb_82_31 bit_82_31 bit_82_32 R_bl
Rbb_82_31 bitb_82_31 bitb_82_32 R_bl
Cb_82_31 bit_82_31 gnd C_bl
Cbb_82_31 bitb_82_31 gnd C_bl
Rb_82_32 bit_82_32 bit_82_33 R_bl
Rbb_82_32 bitb_82_32 bitb_82_33 R_bl
Cb_82_32 bit_82_32 gnd C_bl
Cbb_82_32 bitb_82_32 gnd C_bl
Rb_82_33 bit_82_33 bit_82_34 R_bl
Rbb_82_33 bitb_82_33 bitb_82_34 R_bl
Cb_82_33 bit_82_33 gnd C_bl
Cbb_82_33 bitb_82_33 gnd C_bl
Rb_82_34 bit_82_34 bit_82_35 R_bl
Rbb_82_34 bitb_82_34 bitb_82_35 R_bl
Cb_82_34 bit_82_34 gnd C_bl
Cbb_82_34 bitb_82_34 gnd C_bl
Rb_82_35 bit_82_35 bit_82_36 R_bl
Rbb_82_35 bitb_82_35 bitb_82_36 R_bl
Cb_82_35 bit_82_35 gnd C_bl
Cbb_82_35 bitb_82_35 gnd C_bl
Rb_82_36 bit_82_36 bit_82_37 R_bl
Rbb_82_36 bitb_82_36 bitb_82_37 R_bl
Cb_82_36 bit_82_36 gnd C_bl
Cbb_82_36 bitb_82_36 gnd C_bl
Rb_82_37 bit_82_37 bit_82_38 R_bl
Rbb_82_37 bitb_82_37 bitb_82_38 R_bl
Cb_82_37 bit_82_37 gnd C_bl
Cbb_82_37 bitb_82_37 gnd C_bl
Rb_82_38 bit_82_38 bit_82_39 R_bl
Rbb_82_38 bitb_82_38 bitb_82_39 R_bl
Cb_82_38 bit_82_38 gnd C_bl
Cbb_82_38 bitb_82_38 gnd C_bl
Rb_82_39 bit_82_39 bit_82_40 R_bl
Rbb_82_39 bitb_82_39 bitb_82_40 R_bl
Cb_82_39 bit_82_39 gnd C_bl
Cbb_82_39 bitb_82_39 gnd C_bl
Rb_82_40 bit_82_40 bit_82_41 R_bl
Rbb_82_40 bitb_82_40 bitb_82_41 R_bl
Cb_82_40 bit_82_40 gnd C_bl
Cbb_82_40 bitb_82_40 gnd C_bl
Rb_82_41 bit_82_41 bit_82_42 R_bl
Rbb_82_41 bitb_82_41 bitb_82_42 R_bl
Cb_82_41 bit_82_41 gnd C_bl
Cbb_82_41 bitb_82_41 gnd C_bl
Rb_82_42 bit_82_42 bit_82_43 R_bl
Rbb_82_42 bitb_82_42 bitb_82_43 R_bl
Cb_82_42 bit_82_42 gnd C_bl
Cbb_82_42 bitb_82_42 gnd C_bl
Rb_82_43 bit_82_43 bit_82_44 R_bl
Rbb_82_43 bitb_82_43 bitb_82_44 R_bl
Cb_82_43 bit_82_43 gnd C_bl
Cbb_82_43 bitb_82_43 gnd C_bl
Rb_82_44 bit_82_44 bit_82_45 R_bl
Rbb_82_44 bitb_82_44 bitb_82_45 R_bl
Cb_82_44 bit_82_44 gnd C_bl
Cbb_82_44 bitb_82_44 gnd C_bl
Rb_82_45 bit_82_45 bit_82_46 R_bl
Rbb_82_45 bitb_82_45 bitb_82_46 R_bl
Cb_82_45 bit_82_45 gnd C_bl
Cbb_82_45 bitb_82_45 gnd C_bl
Rb_82_46 bit_82_46 bit_82_47 R_bl
Rbb_82_46 bitb_82_46 bitb_82_47 R_bl
Cb_82_46 bit_82_46 gnd C_bl
Cbb_82_46 bitb_82_46 gnd C_bl
Rb_82_47 bit_82_47 bit_82_48 R_bl
Rbb_82_47 bitb_82_47 bitb_82_48 R_bl
Cb_82_47 bit_82_47 gnd C_bl
Cbb_82_47 bitb_82_47 gnd C_bl
Rb_82_48 bit_82_48 bit_82_49 R_bl
Rbb_82_48 bitb_82_48 bitb_82_49 R_bl
Cb_82_48 bit_82_48 gnd C_bl
Cbb_82_48 bitb_82_48 gnd C_bl
Rb_82_49 bit_82_49 bit_82_50 R_bl
Rbb_82_49 bitb_82_49 bitb_82_50 R_bl
Cb_82_49 bit_82_49 gnd C_bl
Cbb_82_49 bitb_82_49 gnd C_bl
Rb_82_50 bit_82_50 bit_82_51 R_bl
Rbb_82_50 bitb_82_50 bitb_82_51 R_bl
Cb_82_50 bit_82_50 gnd C_bl
Cbb_82_50 bitb_82_50 gnd C_bl
Rb_82_51 bit_82_51 bit_82_52 R_bl
Rbb_82_51 bitb_82_51 bitb_82_52 R_bl
Cb_82_51 bit_82_51 gnd C_bl
Cbb_82_51 bitb_82_51 gnd C_bl
Rb_82_52 bit_82_52 bit_82_53 R_bl
Rbb_82_52 bitb_82_52 bitb_82_53 R_bl
Cb_82_52 bit_82_52 gnd C_bl
Cbb_82_52 bitb_82_52 gnd C_bl
Rb_82_53 bit_82_53 bit_82_54 R_bl
Rbb_82_53 bitb_82_53 bitb_82_54 R_bl
Cb_82_53 bit_82_53 gnd C_bl
Cbb_82_53 bitb_82_53 gnd C_bl
Rb_82_54 bit_82_54 bit_82_55 R_bl
Rbb_82_54 bitb_82_54 bitb_82_55 R_bl
Cb_82_54 bit_82_54 gnd C_bl
Cbb_82_54 bitb_82_54 gnd C_bl
Rb_82_55 bit_82_55 bit_82_56 R_bl
Rbb_82_55 bitb_82_55 bitb_82_56 R_bl
Cb_82_55 bit_82_55 gnd C_bl
Cbb_82_55 bitb_82_55 gnd C_bl
Rb_82_56 bit_82_56 bit_82_57 R_bl
Rbb_82_56 bitb_82_56 bitb_82_57 R_bl
Cb_82_56 bit_82_56 gnd C_bl
Cbb_82_56 bitb_82_56 gnd C_bl
Rb_82_57 bit_82_57 bit_82_58 R_bl
Rbb_82_57 bitb_82_57 bitb_82_58 R_bl
Cb_82_57 bit_82_57 gnd C_bl
Cbb_82_57 bitb_82_57 gnd C_bl
Rb_82_58 bit_82_58 bit_82_59 R_bl
Rbb_82_58 bitb_82_58 bitb_82_59 R_bl
Cb_82_58 bit_82_58 gnd C_bl
Cbb_82_58 bitb_82_58 gnd C_bl
Rb_82_59 bit_82_59 bit_82_60 R_bl
Rbb_82_59 bitb_82_59 bitb_82_60 R_bl
Cb_82_59 bit_82_59 gnd C_bl
Cbb_82_59 bitb_82_59 gnd C_bl
Rb_82_60 bit_82_60 bit_82_61 R_bl
Rbb_82_60 bitb_82_60 bitb_82_61 R_bl
Cb_82_60 bit_82_60 gnd C_bl
Cbb_82_60 bitb_82_60 gnd C_bl
Rb_82_61 bit_82_61 bit_82_62 R_bl
Rbb_82_61 bitb_82_61 bitb_82_62 R_bl
Cb_82_61 bit_82_61 gnd C_bl
Cbb_82_61 bitb_82_61 gnd C_bl
Rb_82_62 bit_82_62 bit_82_63 R_bl
Rbb_82_62 bitb_82_62 bitb_82_63 R_bl
Cb_82_62 bit_82_62 gnd C_bl
Cbb_82_62 bitb_82_62 gnd C_bl
Rb_82_63 bit_82_63 bit_82_64 R_bl
Rbb_82_63 bitb_82_63 bitb_82_64 R_bl
Cb_82_63 bit_82_63 gnd C_bl
Cbb_82_63 bitb_82_63 gnd C_bl
Rb_82_64 bit_82_64 bit_82_65 R_bl
Rbb_82_64 bitb_82_64 bitb_82_65 R_bl
Cb_82_64 bit_82_64 gnd C_bl
Cbb_82_64 bitb_82_64 gnd C_bl
Rb_82_65 bit_82_65 bit_82_66 R_bl
Rbb_82_65 bitb_82_65 bitb_82_66 R_bl
Cb_82_65 bit_82_65 gnd C_bl
Cbb_82_65 bitb_82_65 gnd C_bl
Rb_82_66 bit_82_66 bit_82_67 R_bl
Rbb_82_66 bitb_82_66 bitb_82_67 R_bl
Cb_82_66 bit_82_66 gnd C_bl
Cbb_82_66 bitb_82_66 gnd C_bl
Rb_82_67 bit_82_67 bit_82_68 R_bl
Rbb_82_67 bitb_82_67 bitb_82_68 R_bl
Cb_82_67 bit_82_67 gnd C_bl
Cbb_82_67 bitb_82_67 gnd C_bl
Rb_82_68 bit_82_68 bit_82_69 R_bl
Rbb_82_68 bitb_82_68 bitb_82_69 R_bl
Cb_82_68 bit_82_68 gnd C_bl
Cbb_82_68 bitb_82_68 gnd C_bl
Rb_82_69 bit_82_69 bit_82_70 R_bl
Rbb_82_69 bitb_82_69 bitb_82_70 R_bl
Cb_82_69 bit_82_69 gnd C_bl
Cbb_82_69 bitb_82_69 gnd C_bl
Rb_82_70 bit_82_70 bit_82_71 R_bl
Rbb_82_70 bitb_82_70 bitb_82_71 R_bl
Cb_82_70 bit_82_70 gnd C_bl
Cbb_82_70 bitb_82_70 gnd C_bl
Rb_82_71 bit_82_71 bit_82_72 R_bl
Rbb_82_71 bitb_82_71 bitb_82_72 R_bl
Cb_82_71 bit_82_71 gnd C_bl
Cbb_82_71 bitb_82_71 gnd C_bl
Rb_82_72 bit_82_72 bit_82_73 R_bl
Rbb_82_72 bitb_82_72 bitb_82_73 R_bl
Cb_82_72 bit_82_72 gnd C_bl
Cbb_82_72 bitb_82_72 gnd C_bl
Rb_82_73 bit_82_73 bit_82_74 R_bl
Rbb_82_73 bitb_82_73 bitb_82_74 R_bl
Cb_82_73 bit_82_73 gnd C_bl
Cbb_82_73 bitb_82_73 gnd C_bl
Rb_82_74 bit_82_74 bit_82_75 R_bl
Rbb_82_74 bitb_82_74 bitb_82_75 R_bl
Cb_82_74 bit_82_74 gnd C_bl
Cbb_82_74 bitb_82_74 gnd C_bl
Rb_82_75 bit_82_75 bit_82_76 R_bl
Rbb_82_75 bitb_82_75 bitb_82_76 R_bl
Cb_82_75 bit_82_75 gnd C_bl
Cbb_82_75 bitb_82_75 gnd C_bl
Rb_82_76 bit_82_76 bit_82_77 R_bl
Rbb_82_76 bitb_82_76 bitb_82_77 R_bl
Cb_82_76 bit_82_76 gnd C_bl
Cbb_82_76 bitb_82_76 gnd C_bl
Rb_82_77 bit_82_77 bit_82_78 R_bl
Rbb_82_77 bitb_82_77 bitb_82_78 R_bl
Cb_82_77 bit_82_77 gnd C_bl
Cbb_82_77 bitb_82_77 gnd C_bl
Rb_82_78 bit_82_78 bit_82_79 R_bl
Rbb_82_78 bitb_82_78 bitb_82_79 R_bl
Cb_82_78 bit_82_78 gnd C_bl
Cbb_82_78 bitb_82_78 gnd C_bl
Rb_82_79 bit_82_79 bit_82_80 R_bl
Rbb_82_79 bitb_82_79 bitb_82_80 R_bl
Cb_82_79 bit_82_79 gnd C_bl
Cbb_82_79 bitb_82_79 gnd C_bl
Rb_82_80 bit_82_80 bit_82_81 R_bl
Rbb_82_80 bitb_82_80 bitb_82_81 R_bl
Cb_82_80 bit_82_80 gnd C_bl
Cbb_82_80 bitb_82_80 gnd C_bl
Rb_82_81 bit_82_81 bit_82_82 R_bl
Rbb_82_81 bitb_82_81 bitb_82_82 R_bl
Cb_82_81 bit_82_81 gnd C_bl
Cbb_82_81 bitb_82_81 gnd C_bl
Rb_82_82 bit_82_82 bit_82_83 R_bl
Rbb_82_82 bitb_82_82 bitb_82_83 R_bl
Cb_82_82 bit_82_82 gnd C_bl
Cbb_82_82 bitb_82_82 gnd C_bl
Rb_82_83 bit_82_83 bit_82_84 R_bl
Rbb_82_83 bitb_82_83 bitb_82_84 R_bl
Cb_82_83 bit_82_83 gnd C_bl
Cbb_82_83 bitb_82_83 gnd C_bl
Rb_82_84 bit_82_84 bit_82_85 R_bl
Rbb_82_84 bitb_82_84 bitb_82_85 R_bl
Cb_82_84 bit_82_84 gnd C_bl
Cbb_82_84 bitb_82_84 gnd C_bl
Rb_82_85 bit_82_85 bit_82_86 R_bl
Rbb_82_85 bitb_82_85 bitb_82_86 R_bl
Cb_82_85 bit_82_85 gnd C_bl
Cbb_82_85 bitb_82_85 gnd C_bl
Rb_82_86 bit_82_86 bit_82_87 R_bl
Rbb_82_86 bitb_82_86 bitb_82_87 R_bl
Cb_82_86 bit_82_86 gnd C_bl
Cbb_82_86 bitb_82_86 gnd C_bl
Rb_82_87 bit_82_87 bit_82_88 R_bl
Rbb_82_87 bitb_82_87 bitb_82_88 R_bl
Cb_82_87 bit_82_87 gnd C_bl
Cbb_82_87 bitb_82_87 gnd C_bl
Rb_82_88 bit_82_88 bit_82_89 R_bl
Rbb_82_88 bitb_82_88 bitb_82_89 R_bl
Cb_82_88 bit_82_88 gnd C_bl
Cbb_82_88 bitb_82_88 gnd C_bl
Rb_82_89 bit_82_89 bit_82_90 R_bl
Rbb_82_89 bitb_82_89 bitb_82_90 R_bl
Cb_82_89 bit_82_89 gnd C_bl
Cbb_82_89 bitb_82_89 gnd C_bl
Rb_82_90 bit_82_90 bit_82_91 R_bl
Rbb_82_90 bitb_82_90 bitb_82_91 R_bl
Cb_82_90 bit_82_90 gnd C_bl
Cbb_82_90 bitb_82_90 gnd C_bl
Rb_82_91 bit_82_91 bit_82_92 R_bl
Rbb_82_91 bitb_82_91 bitb_82_92 R_bl
Cb_82_91 bit_82_91 gnd C_bl
Cbb_82_91 bitb_82_91 gnd C_bl
Rb_82_92 bit_82_92 bit_82_93 R_bl
Rbb_82_92 bitb_82_92 bitb_82_93 R_bl
Cb_82_92 bit_82_92 gnd C_bl
Cbb_82_92 bitb_82_92 gnd C_bl
Rb_82_93 bit_82_93 bit_82_94 R_bl
Rbb_82_93 bitb_82_93 bitb_82_94 R_bl
Cb_82_93 bit_82_93 gnd C_bl
Cbb_82_93 bitb_82_93 gnd C_bl
Rb_82_94 bit_82_94 bit_82_95 R_bl
Rbb_82_94 bitb_82_94 bitb_82_95 R_bl
Cb_82_94 bit_82_94 gnd C_bl
Cbb_82_94 bitb_82_94 gnd C_bl
Rb_82_95 bit_82_95 bit_82_96 R_bl
Rbb_82_95 bitb_82_95 bitb_82_96 R_bl
Cb_82_95 bit_82_95 gnd C_bl
Cbb_82_95 bitb_82_95 gnd C_bl
Rb_82_96 bit_82_96 bit_82_97 R_bl
Rbb_82_96 bitb_82_96 bitb_82_97 R_bl
Cb_82_96 bit_82_96 gnd C_bl
Cbb_82_96 bitb_82_96 gnd C_bl
Rb_82_97 bit_82_97 bit_82_98 R_bl
Rbb_82_97 bitb_82_97 bitb_82_98 R_bl
Cb_82_97 bit_82_97 gnd C_bl
Cbb_82_97 bitb_82_97 gnd C_bl
Rb_82_98 bit_82_98 bit_82_99 R_bl
Rbb_82_98 bitb_82_98 bitb_82_99 R_bl
Cb_82_98 bit_82_98 gnd C_bl
Cbb_82_98 bitb_82_98 gnd C_bl
Rb_82_99 bit_82_99 bit_82_100 R_bl
Rbb_82_99 bitb_82_99 bitb_82_100 R_bl
Cb_82_99 bit_82_99 gnd C_bl
Cbb_82_99 bitb_82_99 gnd C_bl
Rb_83_0 bit_83_0 bit_83_1 R_bl
Rbb_83_0 bitb_83_0 bitb_83_1 R_bl
Cb_83_0 bit_83_0 gnd C_bl
Cbb_83_0 bitb_83_0 gnd C_bl
Rb_83_1 bit_83_1 bit_83_2 R_bl
Rbb_83_1 bitb_83_1 bitb_83_2 R_bl
Cb_83_1 bit_83_1 gnd C_bl
Cbb_83_1 bitb_83_1 gnd C_bl
Rb_83_2 bit_83_2 bit_83_3 R_bl
Rbb_83_2 bitb_83_2 bitb_83_3 R_bl
Cb_83_2 bit_83_2 gnd C_bl
Cbb_83_2 bitb_83_2 gnd C_bl
Rb_83_3 bit_83_3 bit_83_4 R_bl
Rbb_83_3 bitb_83_3 bitb_83_4 R_bl
Cb_83_3 bit_83_3 gnd C_bl
Cbb_83_3 bitb_83_3 gnd C_bl
Rb_83_4 bit_83_4 bit_83_5 R_bl
Rbb_83_4 bitb_83_4 bitb_83_5 R_bl
Cb_83_4 bit_83_4 gnd C_bl
Cbb_83_4 bitb_83_4 gnd C_bl
Rb_83_5 bit_83_5 bit_83_6 R_bl
Rbb_83_5 bitb_83_5 bitb_83_6 R_bl
Cb_83_5 bit_83_5 gnd C_bl
Cbb_83_5 bitb_83_5 gnd C_bl
Rb_83_6 bit_83_6 bit_83_7 R_bl
Rbb_83_6 bitb_83_6 bitb_83_7 R_bl
Cb_83_6 bit_83_6 gnd C_bl
Cbb_83_6 bitb_83_6 gnd C_bl
Rb_83_7 bit_83_7 bit_83_8 R_bl
Rbb_83_7 bitb_83_7 bitb_83_8 R_bl
Cb_83_7 bit_83_7 gnd C_bl
Cbb_83_7 bitb_83_7 gnd C_bl
Rb_83_8 bit_83_8 bit_83_9 R_bl
Rbb_83_8 bitb_83_8 bitb_83_9 R_bl
Cb_83_8 bit_83_8 gnd C_bl
Cbb_83_8 bitb_83_8 gnd C_bl
Rb_83_9 bit_83_9 bit_83_10 R_bl
Rbb_83_9 bitb_83_9 bitb_83_10 R_bl
Cb_83_9 bit_83_9 gnd C_bl
Cbb_83_9 bitb_83_9 gnd C_bl
Rb_83_10 bit_83_10 bit_83_11 R_bl
Rbb_83_10 bitb_83_10 bitb_83_11 R_bl
Cb_83_10 bit_83_10 gnd C_bl
Cbb_83_10 bitb_83_10 gnd C_bl
Rb_83_11 bit_83_11 bit_83_12 R_bl
Rbb_83_11 bitb_83_11 bitb_83_12 R_bl
Cb_83_11 bit_83_11 gnd C_bl
Cbb_83_11 bitb_83_11 gnd C_bl
Rb_83_12 bit_83_12 bit_83_13 R_bl
Rbb_83_12 bitb_83_12 bitb_83_13 R_bl
Cb_83_12 bit_83_12 gnd C_bl
Cbb_83_12 bitb_83_12 gnd C_bl
Rb_83_13 bit_83_13 bit_83_14 R_bl
Rbb_83_13 bitb_83_13 bitb_83_14 R_bl
Cb_83_13 bit_83_13 gnd C_bl
Cbb_83_13 bitb_83_13 gnd C_bl
Rb_83_14 bit_83_14 bit_83_15 R_bl
Rbb_83_14 bitb_83_14 bitb_83_15 R_bl
Cb_83_14 bit_83_14 gnd C_bl
Cbb_83_14 bitb_83_14 gnd C_bl
Rb_83_15 bit_83_15 bit_83_16 R_bl
Rbb_83_15 bitb_83_15 bitb_83_16 R_bl
Cb_83_15 bit_83_15 gnd C_bl
Cbb_83_15 bitb_83_15 gnd C_bl
Rb_83_16 bit_83_16 bit_83_17 R_bl
Rbb_83_16 bitb_83_16 bitb_83_17 R_bl
Cb_83_16 bit_83_16 gnd C_bl
Cbb_83_16 bitb_83_16 gnd C_bl
Rb_83_17 bit_83_17 bit_83_18 R_bl
Rbb_83_17 bitb_83_17 bitb_83_18 R_bl
Cb_83_17 bit_83_17 gnd C_bl
Cbb_83_17 bitb_83_17 gnd C_bl
Rb_83_18 bit_83_18 bit_83_19 R_bl
Rbb_83_18 bitb_83_18 bitb_83_19 R_bl
Cb_83_18 bit_83_18 gnd C_bl
Cbb_83_18 bitb_83_18 gnd C_bl
Rb_83_19 bit_83_19 bit_83_20 R_bl
Rbb_83_19 bitb_83_19 bitb_83_20 R_bl
Cb_83_19 bit_83_19 gnd C_bl
Cbb_83_19 bitb_83_19 gnd C_bl
Rb_83_20 bit_83_20 bit_83_21 R_bl
Rbb_83_20 bitb_83_20 bitb_83_21 R_bl
Cb_83_20 bit_83_20 gnd C_bl
Cbb_83_20 bitb_83_20 gnd C_bl
Rb_83_21 bit_83_21 bit_83_22 R_bl
Rbb_83_21 bitb_83_21 bitb_83_22 R_bl
Cb_83_21 bit_83_21 gnd C_bl
Cbb_83_21 bitb_83_21 gnd C_bl
Rb_83_22 bit_83_22 bit_83_23 R_bl
Rbb_83_22 bitb_83_22 bitb_83_23 R_bl
Cb_83_22 bit_83_22 gnd C_bl
Cbb_83_22 bitb_83_22 gnd C_bl
Rb_83_23 bit_83_23 bit_83_24 R_bl
Rbb_83_23 bitb_83_23 bitb_83_24 R_bl
Cb_83_23 bit_83_23 gnd C_bl
Cbb_83_23 bitb_83_23 gnd C_bl
Rb_83_24 bit_83_24 bit_83_25 R_bl
Rbb_83_24 bitb_83_24 bitb_83_25 R_bl
Cb_83_24 bit_83_24 gnd C_bl
Cbb_83_24 bitb_83_24 gnd C_bl
Rb_83_25 bit_83_25 bit_83_26 R_bl
Rbb_83_25 bitb_83_25 bitb_83_26 R_bl
Cb_83_25 bit_83_25 gnd C_bl
Cbb_83_25 bitb_83_25 gnd C_bl
Rb_83_26 bit_83_26 bit_83_27 R_bl
Rbb_83_26 bitb_83_26 bitb_83_27 R_bl
Cb_83_26 bit_83_26 gnd C_bl
Cbb_83_26 bitb_83_26 gnd C_bl
Rb_83_27 bit_83_27 bit_83_28 R_bl
Rbb_83_27 bitb_83_27 bitb_83_28 R_bl
Cb_83_27 bit_83_27 gnd C_bl
Cbb_83_27 bitb_83_27 gnd C_bl
Rb_83_28 bit_83_28 bit_83_29 R_bl
Rbb_83_28 bitb_83_28 bitb_83_29 R_bl
Cb_83_28 bit_83_28 gnd C_bl
Cbb_83_28 bitb_83_28 gnd C_bl
Rb_83_29 bit_83_29 bit_83_30 R_bl
Rbb_83_29 bitb_83_29 bitb_83_30 R_bl
Cb_83_29 bit_83_29 gnd C_bl
Cbb_83_29 bitb_83_29 gnd C_bl
Rb_83_30 bit_83_30 bit_83_31 R_bl
Rbb_83_30 bitb_83_30 bitb_83_31 R_bl
Cb_83_30 bit_83_30 gnd C_bl
Cbb_83_30 bitb_83_30 gnd C_bl
Rb_83_31 bit_83_31 bit_83_32 R_bl
Rbb_83_31 bitb_83_31 bitb_83_32 R_bl
Cb_83_31 bit_83_31 gnd C_bl
Cbb_83_31 bitb_83_31 gnd C_bl
Rb_83_32 bit_83_32 bit_83_33 R_bl
Rbb_83_32 bitb_83_32 bitb_83_33 R_bl
Cb_83_32 bit_83_32 gnd C_bl
Cbb_83_32 bitb_83_32 gnd C_bl
Rb_83_33 bit_83_33 bit_83_34 R_bl
Rbb_83_33 bitb_83_33 bitb_83_34 R_bl
Cb_83_33 bit_83_33 gnd C_bl
Cbb_83_33 bitb_83_33 gnd C_bl
Rb_83_34 bit_83_34 bit_83_35 R_bl
Rbb_83_34 bitb_83_34 bitb_83_35 R_bl
Cb_83_34 bit_83_34 gnd C_bl
Cbb_83_34 bitb_83_34 gnd C_bl
Rb_83_35 bit_83_35 bit_83_36 R_bl
Rbb_83_35 bitb_83_35 bitb_83_36 R_bl
Cb_83_35 bit_83_35 gnd C_bl
Cbb_83_35 bitb_83_35 gnd C_bl
Rb_83_36 bit_83_36 bit_83_37 R_bl
Rbb_83_36 bitb_83_36 bitb_83_37 R_bl
Cb_83_36 bit_83_36 gnd C_bl
Cbb_83_36 bitb_83_36 gnd C_bl
Rb_83_37 bit_83_37 bit_83_38 R_bl
Rbb_83_37 bitb_83_37 bitb_83_38 R_bl
Cb_83_37 bit_83_37 gnd C_bl
Cbb_83_37 bitb_83_37 gnd C_bl
Rb_83_38 bit_83_38 bit_83_39 R_bl
Rbb_83_38 bitb_83_38 bitb_83_39 R_bl
Cb_83_38 bit_83_38 gnd C_bl
Cbb_83_38 bitb_83_38 gnd C_bl
Rb_83_39 bit_83_39 bit_83_40 R_bl
Rbb_83_39 bitb_83_39 bitb_83_40 R_bl
Cb_83_39 bit_83_39 gnd C_bl
Cbb_83_39 bitb_83_39 gnd C_bl
Rb_83_40 bit_83_40 bit_83_41 R_bl
Rbb_83_40 bitb_83_40 bitb_83_41 R_bl
Cb_83_40 bit_83_40 gnd C_bl
Cbb_83_40 bitb_83_40 gnd C_bl
Rb_83_41 bit_83_41 bit_83_42 R_bl
Rbb_83_41 bitb_83_41 bitb_83_42 R_bl
Cb_83_41 bit_83_41 gnd C_bl
Cbb_83_41 bitb_83_41 gnd C_bl
Rb_83_42 bit_83_42 bit_83_43 R_bl
Rbb_83_42 bitb_83_42 bitb_83_43 R_bl
Cb_83_42 bit_83_42 gnd C_bl
Cbb_83_42 bitb_83_42 gnd C_bl
Rb_83_43 bit_83_43 bit_83_44 R_bl
Rbb_83_43 bitb_83_43 bitb_83_44 R_bl
Cb_83_43 bit_83_43 gnd C_bl
Cbb_83_43 bitb_83_43 gnd C_bl
Rb_83_44 bit_83_44 bit_83_45 R_bl
Rbb_83_44 bitb_83_44 bitb_83_45 R_bl
Cb_83_44 bit_83_44 gnd C_bl
Cbb_83_44 bitb_83_44 gnd C_bl
Rb_83_45 bit_83_45 bit_83_46 R_bl
Rbb_83_45 bitb_83_45 bitb_83_46 R_bl
Cb_83_45 bit_83_45 gnd C_bl
Cbb_83_45 bitb_83_45 gnd C_bl
Rb_83_46 bit_83_46 bit_83_47 R_bl
Rbb_83_46 bitb_83_46 bitb_83_47 R_bl
Cb_83_46 bit_83_46 gnd C_bl
Cbb_83_46 bitb_83_46 gnd C_bl
Rb_83_47 bit_83_47 bit_83_48 R_bl
Rbb_83_47 bitb_83_47 bitb_83_48 R_bl
Cb_83_47 bit_83_47 gnd C_bl
Cbb_83_47 bitb_83_47 gnd C_bl
Rb_83_48 bit_83_48 bit_83_49 R_bl
Rbb_83_48 bitb_83_48 bitb_83_49 R_bl
Cb_83_48 bit_83_48 gnd C_bl
Cbb_83_48 bitb_83_48 gnd C_bl
Rb_83_49 bit_83_49 bit_83_50 R_bl
Rbb_83_49 bitb_83_49 bitb_83_50 R_bl
Cb_83_49 bit_83_49 gnd C_bl
Cbb_83_49 bitb_83_49 gnd C_bl
Rb_83_50 bit_83_50 bit_83_51 R_bl
Rbb_83_50 bitb_83_50 bitb_83_51 R_bl
Cb_83_50 bit_83_50 gnd C_bl
Cbb_83_50 bitb_83_50 gnd C_bl
Rb_83_51 bit_83_51 bit_83_52 R_bl
Rbb_83_51 bitb_83_51 bitb_83_52 R_bl
Cb_83_51 bit_83_51 gnd C_bl
Cbb_83_51 bitb_83_51 gnd C_bl
Rb_83_52 bit_83_52 bit_83_53 R_bl
Rbb_83_52 bitb_83_52 bitb_83_53 R_bl
Cb_83_52 bit_83_52 gnd C_bl
Cbb_83_52 bitb_83_52 gnd C_bl
Rb_83_53 bit_83_53 bit_83_54 R_bl
Rbb_83_53 bitb_83_53 bitb_83_54 R_bl
Cb_83_53 bit_83_53 gnd C_bl
Cbb_83_53 bitb_83_53 gnd C_bl
Rb_83_54 bit_83_54 bit_83_55 R_bl
Rbb_83_54 bitb_83_54 bitb_83_55 R_bl
Cb_83_54 bit_83_54 gnd C_bl
Cbb_83_54 bitb_83_54 gnd C_bl
Rb_83_55 bit_83_55 bit_83_56 R_bl
Rbb_83_55 bitb_83_55 bitb_83_56 R_bl
Cb_83_55 bit_83_55 gnd C_bl
Cbb_83_55 bitb_83_55 gnd C_bl
Rb_83_56 bit_83_56 bit_83_57 R_bl
Rbb_83_56 bitb_83_56 bitb_83_57 R_bl
Cb_83_56 bit_83_56 gnd C_bl
Cbb_83_56 bitb_83_56 gnd C_bl
Rb_83_57 bit_83_57 bit_83_58 R_bl
Rbb_83_57 bitb_83_57 bitb_83_58 R_bl
Cb_83_57 bit_83_57 gnd C_bl
Cbb_83_57 bitb_83_57 gnd C_bl
Rb_83_58 bit_83_58 bit_83_59 R_bl
Rbb_83_58 bitb_83_58 bitb_83_59 R_bl
Cb_83_58 bit_83_58 gnd C_bl
Cbb_83_58 bitb_83_58 gnd C_bl
Rb_83_59 bit_83_59 bit_83_60 R_bl
Rbb_83_59 bitb_83_59 bitb_83_60 R_bl
Cb_83_59 bit_83_59 gnd C_bl
Cbb_83_59 bitb_83_59 gnd C_bl
Rb_83_60 bit_83_60 bit_83_61 R_bl
Rbb_83_60 bitb_83_60 bitb_83_61 R_bl
Cb_83_60 bit_83_60 gnd C_bl
Cbb_83_60 bitb_83_60 gnd C_bl
Rb_83_61 bit_83_61 bit_83_62 R_bl
Rbb_83_61 bitb_83_61 bitb_83_62 R_bl
Cb_83_61 bit_83_61 gnd C_bl
Cbb_83_61 bitb_83_61 gnd C_bl
Rb_83_62 bit_83_62 bit_83_63 R_bl
Rbb_83_62 bitb_83_62 bitb_83_63 R_bl
Cb_83_62 bit_83_62 gnd C_bl
Cbb_83_62 bitb_83_62 gnd C_bl
Rb_83_63 bit_83_63 bit_83_64 R_bl
Rbb_83_63 bitb_83_63 bitb_83_64 R_bl
Cb_83_63 bit_83_63 gnd C_bl
Cbb_83_63 bitb_83_63 gnd C_bl
Rb_83_64 bit_83_64 bit_83_65 R_bl
Rbb_83_64 bitb_83_64 bitb_83_65 R_bl
Cb_83_64 bit_83_64 gnd C_bl
Cbb_83_64 bitb_83_64 gnd C_bl
Rb_83_65 bit_83_65 bit_83_66 R_bl
Rbb_83_65 bitb_83_65 bitb_83_66 R_bl
Cb_83_65 bit_83_65 gnd C_bl
Cbb_83_65 bitb_83_65 gnd C_bl
Rb_83_66 bit_83_66 bit_83_67 R_bl
Rbb_83_66 bitb_83_66 bitb_83_67 R_bl
Cb_83_66 bit_83_66 gnd C_bl
Cbb_83_66 bitb_83_66 gnd C_bl
Rb_83_67 bit_83_67 bit_83_68 R_bl
Rbb_83_67 bitb_83_67 bitb_83_68 R_bl
Cb_83_67 bit_83_67 gnd C_bl
Cbb_83_67 bitb_83_67 gnd C_bl
Rb_83_68 bit_83_68 bit_83_69 R_bl
Rbb_83_68 bitb_83_68 bitb_83_69 R_bl
Cb_83_68 bit_83_68 gnd C_bl
Cbb_83_68 bitb_83_68 gnd C_bl
Rb_83_69 bit_83_69 bit_83_70 R_bl
Rbb_83_69 bitb_83_69 bitb_83_70 R_bl
Cb_83_69 bit_83_69 gnd C_bl
Cbb_83_69 bitb_83_69 gnd C_bl
Rb_83_70 bit_83_70 bit_83_71 R_bl
Rbb_83_70 bitb_83_70 bitb_83_71 R_bl
Cb_83_70 bit_83_70 gnd C_bl
Cbb_83_70 bitb_83_70 gnd C_bl
Rb_83_71 bit_83_71 bit_83_72 R_bl
Rbb_83_71 bitb_83_71 bitb_83_72 R_bl
Cb_83_71 bit_83_71 gnd C_bl
Cbb_83_71 bitb_83_71 gnd C_bl
Rb_83_72 bit_83_72 bit_83_73 R_bl
Rbb_83_72 bitb_83_72 bitb_83_73 R_bl
Cb_83_72 bit_83_72 gnd C_bl
Cbb_83_72 bitb_83_72 gnd C_bl
Rb_83_73 bit_83_73 bit_83_74 R_bl
Rbb_83_73 bitb_83_73 bitb_83_74 R_bl
Cb_83_73 bit_83_73 gnd C_bl
Cbb_83_73 bitb_83_73 gnd C_bl
Rb_83_74 bit_83_74 bit_83_75 R_bl
Rbb_83_74 bitb_83_74 bitb_83_75 R_bl
Cb_83_74 bit_83_74 gnd C_bl
Cbb_83_74 bitb_83_74 gnd C_bl
Rb_83_75 bit_83_75 bit_83_76 R_bl
Rbb_83_75 bitb_83_75 bitb_83_76 R_bl
Cb_83_75 bit_83_75 gnd C_bl
Cbb_83_75 bitb_83_75 gnd C_bl
Rb_83_76 bit_83_76 bit_83_77 R_bl
Rbb_83_76 bitb_83_76 bitb_83_77 R_bl
Cb_83_76 bit_83_76 gnd C_bl
Cbb_83_76 bitb_83_76 gnd C_bl
Rb_83_77 bit_83_77 bit_83_78 R_bl
Rbb_83_77 bitb_83_77 bitb_83_78 R_bl
Cb_83_77 bit_83_77 gnd C_bl
Cbb_83_77 bitb_83_77 gnd C_bl
Rb_83_78 bit_83_78 bit_83_79 R_bl
Rbb_83_78 bitb_83_78 bitb_83_79 R_bl
Cb_83_78 bit_83_78 gnd C_bl
Cbb_83_78 bitb_83_78 gnd C_bl
Rb_83_79 bit_83_79 bit_83_80 R_bl
Rbb_83_79 bitb_83_79 bitb_83_80 R_bl
Cb_83_79 bit_83_79 gnd C_bl
Cbb_83_79 bitb_83_79 gnd C_bl
Rb_83_80 bit_83_80 bit_83_81 R_bl
Rbb_83_80 bitb_83_80 bitb_83_81 R_bl
Cb_83_80 bit_83_80 gnd C_bl
Cbb_83_80 bitb_83_80 gnd C_bl
Rb_83_81 bit_83_81 bit_83_82 R_bl
Rbb_83_81 bitb_83_81 bitb_83_82 R_bl
Cb_83_81 bit_83_81 gnd C_bl
Cbb_83_81 bitb_83_81 gnd C_bl
Rb_83_82 bit_83_82 bit_83_83 R_bl
Rbb_83_82 bitb_83_82 bitb_83_83 R_bl
Cb_83_82 bit_83_82 gnd C_bl
Cbb_83_82 bitb_83_82 gnd C_bl
Rb_83_83 bit_83_83 bit_83_84 R_bl
Rbb_83_83 bitb_83_83 bitb_83_84 R_bl
Cb_83_83 bit_83_83 gnd C_bl
Cbb_83_83 bitb_83_83 gnd C_bl
Rb_83_84 bit_83_84 bit_83_85 R_bl
Rbb_83_84 bitb_83_84 bitb_83_85 R_bl
Cb_83_84 bit_83_84 gnd C_bl
Cbb_83_84 bitb_83_84 gnd C_bl
Rb_83_85 bit_83_85 bit_83_86 R_bl
Rbb_83_85 bitb_83_85 bitb_83_86 R_bl
Cb_83_85 bit_83_85 gnd C_bl
Cbb_83_85 bitb_83_85 gnd C_bl
Rb_83_86 bit_83_86 bit_83_87 R_bl
Rbb_83_86 bitb_83_86 bitb_83_87 R_bl
Cb_83_86 bit_83_86 gnd C_bl
Cbb_83_86 bitb_83_86 gnd C_bl
Rb_83_87 bit_83_87 bit_83_88 R_bl
Rbb_83_87 bitb_83_87 bitb_83_88 R_bl
Cb_83_87 bit_83_87 gnd C_bl
Cbb_83_87 bitb_83_87 gnd C_bl
Rb_83_88 bit_83_88 bit_83_89 R_bl
Rbb_83_88 bitb_83_88 bitb_83_89 R_bl
Cb_83_88 bit_83_88 gnd C_bl
Cbb_83_88 bitb_83_88 gnd C_bl
Rb_83_89 bit_83_89 bit_83_90 R_bl
Rbb_83_89 bitb_83_89 bitb_83_90 R_bl
Cb_83_89 bit_83_89 gnd C_bl
Cbb_83_89 bitb_83_89 gnd C_bl
Rb_83_90 bit_83_90 bit_83_91 R_bl
Rbb_83_90 bitb_83_90 bitb_83_91 R_bl
Cb_83_90 bit_83_90 gnd C_bl
Cbb_83_90 bitb_83_90 gnd C_bl
Rb_83_91 bit_83_91 bit_83_92 R_bl
Rbb_83_91 bitb_83_91 bitb_83_92 R_bl
Cb_83_91 bit_83_91 gnd C_bl
Cbb_83_91 bitb_83_91 gnd C_bl
Rb_83_92 bit_83_92 bit_83_93 R_bl
Rbb_83_92 bitb_83_92 bitb_83_93 R_bl
Cb_83_92 bit_83_92 gnd C_bl
Cbb_83_92 bitb_83_92 gnd C_bl
Rb_83_93 bit_83_93 bit_83_94 R_bl
Rbb_83_93 bitb_83_93 bitb_83_94 R_bl
Cb_83_93 bit_83_93 gnd C_bl
Cbb_83_93 bitb_83_93 gnd C_bl
Rb_83_94 bit_83_94 bit_83_95 R_bl
Rbb_83_94 bitb_83_94 bitb_83_95 R_bl
Cb_83_94 bit_83_94 gnd C_bl
Cbb_83_94 bitb_83_94 gnd C_bl
Rb_83_95 bit_83_95 bit_83_96 R_bl
Rbb_83_95 bitb_83_95 bitb_83_96 R_bl
Cb_83_95 bit_83_95 gnd C_bl
Cbb_83_95 bitb_83_95 gnd C_bl
Rb_83_96 bit_83_96 bit_83_97 R_bl
Rbb_83_96 bitb_83_96 bitb_83_97 R_bl
Cb_83_96 bit_83_96 gnd C_bl
Cbb_83_96 bitb_83_96 gnd C_bl
Rb_83_97 bit_83_97 bit_83_98 R_bl
Rbb_83_97 bitb_83_97 bitb_83_98 R_bl
Cb_83_97 bit_83_97 gnd C_bl
Cbb_83_97 bitb_83_97 gnd C_bl
Rb_83_98 bit_83_98 bit_83_99 R_bl
Rbb_83_98 bitb_83_98 bitb_83_99 R_bl
Cb_83_98 bit_83_98 gnd C_bl
Cbb_83_98 bitb_83_98 gnd C_bl
Rb_83_99 bit_83_99 bit_83_100 R_bl
Rbb_83_99 bitb_83_99 bitb_83_100 R_bl
Cb_83_99 bit_83_99 gnd C_bl
Cbb_83_99 bitb_83_99 gnd C_bl
Rb_84_0 bit_84_0 bit_84_1 R_bl
Rbb_84_0 bitb_84_0 bitb_84_1 R_bl
Cb_84_0 bit_84_0 gnd C_bl
Cbb_84_0 bitb_84_0 gnd C_bl
Rb_84_1 bit_84_1 bit_84_2 R_bl
Rbb_84_1 bitb_84_1 bitb_84_2 R_bl
Cb_84_1 bit_84_1 gnd C_bl
Cbb_84_1 bitb_84_1 gnd C_bl
Rb_84_2 bit_84_2 bit_84_3 R_bl
Rbb_84_2 bitb_84_2 bitb_84_3 R_bl
Cb_84_2 bit_84_2 gnd C_bl
Cbb_84_2 bitb_84_2 gnd C_bl
Rb_84_3 bit_84_3 bit_84_4 R_bl
Rbb_84_3 bitb_84_3 bitb_84_4 R_bl
Cb_84_3 bit_84_3 gnd C_bl
Cbb_84_3 bitb_84_3 gnd C_bl
Rb_84_4 bit_84_4 bit_84_5 R_bl
Rbb_84_4 bitb_84_4 bitb_84_5 R_bl
Cb_84_4 bit_84_4 gnd C_bl
Cbb_84_4 bitb_84_4 gnd C_bl
Rb_84_5 bit_84_5 bit_84_6 R_bl
Rbb_84_5 bitb_84_5 bitb_84_6 R_bl
Cb_84_5 bit_84_5 gnd C_bl
Cbb_84_5 bitb_84_5 gnd C_bl
Rb_84_6 bit_84_6 bit_84_7 R_bl
Rbb_84_6 bitb_84_6 bitb_84_7 R_bl
Cb_84_6 bit_84_6 gnd C_bl
Cbb_84_6 bitb_84_6 gnd C_bl
Rb_84_7 bit_84_7 bit_84_8 R_bl
Rbb_84_7 bitb_84_7 bitb_84_8 R_bl
Cb_84_7 bit_84_7 gnd C_bl
Cbb_84_7 bitb_84_7 gnd C_bl
Rb_84_8 bit_84_8 bit_84_9 R_bl
Rbb_84_8 bitb_84_8 bitb_84_9 R_bl
Cb_84_8 bit_84_8 gnd C_bl
Cbb_84_8 bitb_84_8 gnd C_bl
Rb_84_9 bit_84_9 bit_84_10 R_bl
Rbb_84_9 bitb_84_9 bitb_84_10 R_bl
Cb_84_9 bit_84_9 gnd C_bl
Cbb_84_9 bitb_84_9 gnd C_bl
Rb_84_10 bit_84_10 bit_84_11 R_bl
Rbb_84_10 bitb_84_10 bitb_84_11 R_bl
Cb_84_10 bit_84_10 gnd C_bl
Cbb_84_10 bitb_84_10 gnd C_bl
Rb_84_11 bit_84_11 bit_84_12 R_bl
Rbb_84_11 bitb_84_11 bitb_84_12 R_bl
Cb_84_11 bit_84_11 gnd C_bl
Cbb_84_11 bitb_84_11 gnd C_bl
Rb_84_12 bit_84_12 bit_84_13 R_bl
Rbb_84_12 bitb_84_12 bitb_84_13 R_bl
Cb_84_12 bit_84_12 gnd C_bl
Cbb_84_12 bitb_84_12 gnd C_bl
Rb_84_13 bit_84_13 bit_84_14 R_bl
Rbb_84_13 bitb_84_13 bitb_84_14 R_bl
Cb_84_13 bit_84_13 gnd C_bl
Cbb_84_13 bitb_84_13 gnd C_bl
Rb_84_14 bit_84_14 bit_84_15 R_bl
Rbb_84_14 bitb_84_14 bitb_84_15 R_bl
Cb_84_14 bit_84_14 gnd C_bl
Cbb_84_14 bitb_84_14 gnd C_bl
Rb_84_15 bit_84_15 bit_84_16 R_bl
Rbb_84_15 bitb_84_15 bitb_84_16 R_bl
Cb_84_15 bit_84_15 gnd C_bl
Cbb_84_15 bitb_84_15 gnd C_bl
Rb_84_16 bit_84_16 bit_84_17 R_bl
Rbb_84_16 bitb_84_16 bitb_84_17 R_bl
Cb_84_16 bit_84_16 gnd C_bl
Cbb_84_16 bitb_84_16 gnd C_bl
Rb_84_17 bit_84_17 bit_84_18 R_bl
Rbb_84_17 bitb_84_17 bitb_84_18 R_bl
Cb_84_17 bit_84_17 gnd C_bl
Cbb_84_17 bitb_84_17 gnd C_bl
Rb_84_18 bit_84_18 bit_84_19 R_bl
Rbb_84_18 bitb_84_18 bitb_84_19 R_bl
Cb_84_18 bit_84_18 gnd C_bl
Cbb_84_18 bitb_84_18 gnd C_bl
Rb_84_19 bit_84_19 bit_84_20 R_bl
Rbb_84_19 bitb_84_19 bitb_84_20 R_bl
Cb_84_19 bit_84_19 gnd C_bl
Cbb_84_19 bitb_84_19 gnd C_bl
Rb_84_20 bit_84_20 bit_84_21 R_bl
Rbb_84_20 bitb_84_20 bitb_84_21 R_bl
Cb_84_20 bit_84_20 gnd C_bl
Cbb_84_20 bitb_84_20 gnd C_bl
Rb_84_21 bit_84_21 bit_84_22 R_bl
Rbb_84_21 bitb_84_21 bitb_84_22 R_bl
Cb_84_21 bit_84_21 gnd C_bl
Cbb_84_21 bitb_84_21 gnd C_bl
Rb_84_22 bit_84_22 bit_84_23 R_bl
Rbb_84_22 bitb_84_22 bitb_84_23 R_bl
Cb_84_22 bit_84_22 gnd C_bl
Cbb_84_22 bitb_84_22 gnd C_bl
Rb_84_23 bit_84_23 bit_84_24 R_bl
Rbb_84_23 bitb_84_23 bitb_84_24 R_bl
Cb_84_23 bit_84_23 gnd C_bl
Cbb_84_23 bitb_84_23 gnd C_bl
Rb_84_24 bit_84_24 bit_84_25 R_bl
Rbb_84_24 bitb_84_24 bitb_84_25 R_bl
Cb_84_24 bit_84_24 gnd C_bl
Cbb_84_24 bitb_84_24 gnd C_bl
Rb_84_25 bit_84_25 bit_84_26 R_bl
Rbb_84_25 bitb_84_25 bitb_84_26 R_bl
Cb_84_25 bit_84_25 gnd C_bl
Cbb_84_25 bitb_84_25 gnd C_bl
Rb_84_26 bit_84_26 bit_84_27 R_bl
Rbb_84_26 bitb_84_26 bitb_84_27 R_bl
Cb_84_26 bit_84_26 gnd C_bl
Cbb_84_26 bitb_84_26 gnd C_bl
Rb_84_27 bit_84_27 bit_84_28 R_bl
Rbb_84_27 bitb_84_27 bitb_84_28 R_bl
Cb_84_27 bit_84_27 gnd C_bl
Cbb_84_27 bitb_84_27 gnd C_bl
Rb_84_28 bit_84_28 bit_84_29 R_bl
Rbb_84_28 bitb_84_28 bitb_84_29 R_bl
Cb_84_28 bit_84_28 gnd C_bl
Cbb_84_28 bitb_84_28 gnd C_bl
Rb_84_29 bit_84_29 bit_84_30 R_bl
Rbb_84_29 bitb_84_29 bitb_84_30 R_bl
Cb_84_29 bit_84_29 gnd C_bl
Cbb_84_29 bitb_84_29 gnd C_bl
Rb_84_30 bit_84_30 bit_84_31 R_bl
Rbb_84_30 bitb_84_30 bitb_84_31 R_bl
Cb_84_30 bit_84_30 gnd C_bl
Cbb_84_30 bitb_84_30 gnd C_bl
Rb_84_31 bit_84_31 bit_84_32 R_bl
Rbb_84_31 bitb_84_31 bitb_84_32 R_bl
Cb_84_31 bit_84_31 gnd C_bl
Cbb_84_31 bitb_84_31 gnd C_bl
Rb_84_32 bit_84_32 bit_84_33 R_bl
Rbb_84_32 bitb_84_32 bitb_84_33 R_bl
Cb_84_32 bit_84_32 gnd C_bl
Cbb_84_32 bitb_84_32 gnd C_bl
Rb_84_33 bit_84_33 bit_84_34 R_bl
Rbb_84_33 bitb_84_33 bitb_84_34 R_bl
Cb_84_33 bit_84_33 gnd C_bl
Cbb_84_33 bitb_84_33 gnd C_bl
Rb_84_34 bit_84_34 bit_84_35 R_bl
Rbb_84_34 bitb_84_34 bitb_84_35 R_bl
Cb_84_34 bit_84_34 gnd C_bl
Cbb_84_34 bitb_84_34 gnd C_bl
Rb_84_35 bit_84_35 bit_84_36 R_bl
Rbb_84_35 bitb_84_35 bitb_84_36 R_bl
Cb_84_35 bit_84_35 gnd C_bl
Cbb_84_35 bitb_84_35 gnd C_bl
Rb_84_36 bit_84_36 bit_84_37 R_bl
Rbb_84_36 bitb_84_36 bitb_84_37 R_bl
Cb_84_36 bit_84_36 gnd C_bl
Cbb_84_36 bitb_84_36 gnd C_bl
Rb_84_37 bit_84_37 bit_84_38 R_bl
Rbb_84_37 bitb_84_37 bitb_84_38 R_bl
Cb_84_37 bit_84_37 gnd C_bl
Cbb_84_37 bitb_84_37 gnd C_bl
Rb_84_38 bit_84_38 bit_84_39 R_bl
Rbb_84_38 bitb_84_38 bitb_84_39 R_bl
Cb_84_38 bit_84_38 gnd C_bl
Cbb_84_38 bitb_84_38 gnd C_bl
Rb_84_39 bit_84_39 bit_84_40 R_bl
Rbb_84_39 bitb_84_39 bitb_84_40 R_bl
Cb_84_39 bit_84_39 gnd C_bl
Cbb_84_39 bitb_84_39 gnd C_bl
Rb_84_40 bit_84_40 bit_84_41 R_bl
Rbb_84_40 bitb_84_40 bitb_84_41 R_bl
Cb_84_40 bit_84_40 gnd C_bl
Cbb_84_40 bitb_84_40 gnd C_bl
Rb_84_41 bit_84_41 bit_84_42 R_bl
Rbb_84_41 bitb_84_41 bitb_84_42 R_bl
Cb_84_41 bit_84_41 gnd C_bl
Cbb_84_41 bitb_84_41 gnd C_bl
Rb_84_42 bit_84_42 bit_84_43 R_bl
Rbb_84_42 bitb_84_42 bitb_84_43 R_bl
Cb_84_42 bit_84_42 gnd C_bl
Cbb_84_42 bitb_84_42 gnd C_bl
Rb_84_43 bit_84_43 bit_84_44 R_bl
Rbb_84_43 bitb_84_43 bitb_84_44 R_bl
Cb_84_43 bit_84_43 gnd C_bl
Cbb_84_43 bitb_84_43 gnd C_bl
Rb_84_44 bit_84_44 bit_84_45 R_bl
Rbb_84_44 bitb_84_44 bitb_84_45 R_bl
Cb_84_44 bit_84_44 gnd C_bl
Cbb_84_44 bitb_84_44 gnd C_bl
Rb_84_45 bit_84_45 bit_84_46 R_bl
Rbb_84_45 bitb_84_45 bitb_84_46 R_bl
Cb_84_45 bit_84_45 gnd C_bl
Cbb_84_45 bitb_84_45 gnd C_bl
Rb_84_46 bit_84_46 bit_84_47 R_bl
Rbb_84_46 bitb_84_46 bitb_84_47 R_bl
Cb_84_46 bit_84_46 gnd C_bl
Cbb_84_46 bitb_84_46 gnd C_bl
Rb_84_47 bit_84_47 bit_84_48 R_bl
Rbb_84_47 bitb_84_47 bitb_84_48 R_bl
Cb_84_47 bit_84_47 gnd C_bl
Cbb_84_47 bitb_84_47 gnd C_bl
Rb_84_48 bit_84_48 bit_84_49 R_bl
Rbb_84_48 bitb_84_48 bitb_84_49 R_bl
Cb_84_48 bit_84_48 gnd C_bl
Cbb_84_48 bitb_84_48 gnd C_bl
Rb_84_49 bit_84_49 bit_84_50 R_bl
Rbb_84_49 bitb_84_49 bitb_84_50 R_bl
Cb_84_49 bit_84_49 gnd C_bl
Cbb_84_49 bitb_84_49 gnd C_bl
Rb_84_50 bit_84_50 bit_84_51 R_bl
Rbb_84_50 bitb_84_50 bitb_84_51 R_bl
Cb_84_50 bit_84_50 gnd C_bl
Cbb_84_50 bitb_84_50 gnd C_bl
Rb_84_51 bit_84_51 bit_84_52 R_bl
Rbb_84_51 bitb_84_51 bitb_84_52 R_bl
Cb_84_51 bit_84_51 gnd C_bl
Cbb_84_51 bitb_84_51 gnd C_bl
Rb_84_52 bit_84_52 bit_84_53 R_bl
Rbb_84_52 bitb_84_52 bitb_84_53 R_bl
Cb_84_52 bit_84_52 gnd C_bl
Cbb_84_52 bitb_84_52 gnd C_bl
Rb_84_53 bit_84_53 bit_84_54 R_bl
Rbb_84_53 bitb_84_53 bitb_84_54 R_bl
Cb_84_53 bit_84_53 gnd C_bl
Cbb_84_53 bitb_84_53 gnd C_bl
Rb_84_54 bit_84_54 bit_84_55 R_bl
Rbb_84_54 bitb_84_54 bitb_84_55 R_bl
Cb_84_54 bit_84_54 gnd C_bl
Cbb_84_54 bitb_84_54 gnd C_bl
Rb_84_55 bit_84_55 bit_84_56 R_bl
Rbb_84_55 bitb_84_55 bitb_84_56 R_bl
Cb_84_55 bit_84_55 gnd C_bl
Cbb_84_55 bitb_84_55 gnd C_bl
Rb_84_56 bit_84_56 bit_84_57 R_bl
Rbb_84_56 bitb_84_56 bitb_84_57 R_bl
Cb_84_56 bit_84_56 gnd C_bl
Cbb_84_56 bitb_84_56 gnd C_bl
Rb_84_57 bit_84_57 bit_84_58 R_bl
Rbb_84_57 bitb_84_57 bitb_84_58 R_bl
Cb_84_57 bit_84_57 gnd C_bl
Cbb_84_57 bitb_84_57 gnd C_bl
Rb_84_58 bit_84_58 bit_84_59 R_bl
Rbb_84_58 bitb_84_58 bitb_84_59 R_bl
Cb_84_58 bit_84_58 gnd C_bl
Cbb_84_58 bitb_84_58 gnd C_bl
Rb_84_59 bit_84_59 bit_84_60 R_bl
Rbb_84_59 bitb_84_59 bitb_84_60 R_bl
Cb_84_59 bit_84_59 gnd C_bl
Cbb_84_59 bitb_84_59 gnd C_bl
Rb_84_60 bit_84_60 bit_84_61 R_bl
Rbb_84_60 bitb_84_60 bitb_84_61 R_bl
Cb_84_60 bit_84_60 gnd C_bl
Cbb_84_60 bitb_84_60 gnd C_bl
Rb_84_61 bit_84_61 bit_84_62 R_bl
Rbb_84_61 bitb_84_61 bitb_84_62 R_bl
Cb_84_61 bit_84_61 gnd C_bl
Cbb_84_61 bitb_84_61 gnd C_bl
Rb_84_62 bit_84_62 bit_84_63 R_bl
Rbb_84_62 bitb_84_62 bitb_84_63 R_bl
Cb_84_62 bit_84_62 gnd C_bl
Cbb_84_62 bitb_84_62 gnd C_bl
Rb_84_63 bit_84_63 bit_84_64 R_bl
Rbb_84_63 bitb_84_63 bitb_84_64 R_bl
Cb_84_63 bit_84_63 gnd C_bl
Cbb_84_63 bitb_84_63 gnd C_bl
Rb_84_64 bit_84_64 bit_84_65 R_bl
Rbb_84_64 bitb_84_64 bitb_84_65 R_bl
Cb_84_64 bit_84_64 gnd C_bl
Cbb_84_64 bitb_84_64 gnd C_bl
Rb_84_65 bit_84_65 bit_84_66 R_bl
Rbb_84_65 bitb_84_65 bitb_84_66 R_bl
Cb_84_65 bit_84_65 gnd C_bl
Cbb_84_65 bitb_84_65 gnd C_bl
Rb_84_66 bit_84_66 bit_84_67 R_bl
Rbb_84_66 bitb_84_66 bitb_84_67 R_bl
Cb_84_66 bit_84_66 gnd C_bl
Cbb_84_66 bitb_84_66 gnd C_bl
Rb_84_67 bit_84_67 bit_84_68 R_bl
Rbb_84_67 bitb_84_67 bitb_84_68 R_bl
Cb_84_67 bit_84_67 gnd C_bl
Cbb_84_67 bitb_84_67 gnd C_bl
Rb_84_68 bit_84_68 bit_84_69 R_bl
Rbb_84_68 bitb_84_68 bitb_84_69 R_bl
Cb_84_68 bit_84_68 gnd C_bl
Cbb_84_68 bitb_84_68 gnd C_bl
Rb_84_69 bit_84_69 bit_84_70 R_bl
Rbb_84_69 bitb_84_69 bitb_84_70 R_bl
Cb_84_69 bit_84_69 gnd C_bl
Cbb_84_69 bitb_84_69 gnd C_bl
Rb_84_70 bit_84_70 bit_84_71 R_bl
Rbb_84_70 bitb_84_70 bitb_84_71 R_bl
Cb_84_70 bit_84_70 gnd C_bl
Cbb_84_70 bitb_84_70 gnd C_bl
Rb_84_71 bit_84_71 bit_84_72 R_bl
Rbb_84_71 bitb_84_71 bitb_84_72 R_bl
Cb_84_71 bit_84_71 gnd C_bl
Cbb_84_71 bitb_84_71 gnd C_bl
Rb_84_72 bit_84_72 bit_84_73 R_bl
Rbb_84_72 bitb_84_72 bitb_84_73 R_bl
Cb_84_72 bit_84_72 gnd C_bl
Cbb_84_72 bitb_84_72 gnd C_bl
Rb_84_73 bit_84_73 bit_84_74 R_bl
Rbb_84_73 bitb_84_73 bitb_84_74 R_bl
Cb_84_73 bit_84_73 gnd C_bl
Cbb_84_73 bitb_84_73 gnd C_bl
Rb_84_74 bit_84_74 bit_84_75 R_bl
Rbb_84_74 bitb_84_74 bitb_84_75 R_bl
Cb_84_74 bit_84_74 gnd C_bl
Cbb_84_74 bitb_84_74 gnd C_bl
Rb_84_75 bit_84_75 bit_84_76 R_bl
Rbb_84_75 bitb_84_75 bitb_84_76 R_bl
Cb_84_75 bit_84_75 gnd C_bl
Cbb_84_75 bitb_84_75 gnd C_bl
Rb_84_76 bit_84_76 bit_84_77 R_bl
Rbb_84_76 bitb_84_76 bitb_84_77 R_bl
Cb_84_76 bit_84_76 gnd C_bl
Cbb_84_76 bitb_84_76 gnd C_bl
Rb_84_77 bit_84_77 bit_84_78 R_bl
Rbb_84_77 bitb_84_77 bitb_84_78 R_bl
Cb_84_77 bit_84_77 gnd C_bl
Cbb_84_77 bitb_84_77 gnd C_bl
Rb_84_78 bit_84_78 bit_84_79 R_bl
Rbb_84_78 bitb_84_78 bitb_84_79 R_bl
Cb_84_78 bit_84_78 gnd C_bl
Cbb_84_78 bitb_84_78 gnd C_bl
Rb_84_79 bit_84_79 bit_84_80 R_bl
Rbb_84_79 bitb_84_79 bitb_84_80 R_bl
Cb_84_79 bit_84_79 gnd C_bl
Cbb_84_79 bitb_84_79 gnd C_bl
Rb_84_80 bit_84_80 bit_84_81 R_bl
Rbb_84_80 bitb_84_80 bitb_84_81 R_bl
Cb_84_80 bit_84_80 gnd C_bl
Cbb_84_80 bitb_84_80 gnd C_bl
Rb_84_81 bit_84_81 bit_84_82 R_bl
Rbb_84_81 bitb_84_81 bitb_84_82 R_bl
Cb_84_81 bit_84_81 gnd C_bl
Cbb_84_81 bitb_84_81 gnd C_bl
Rb_84_82 bit_84_82 bit_84_83 R_bl
Rbb_84_82 bitb_84_82 bitb_84_83 R_bl
Cb_84_82 bit_84_82 gnd C_bl
Cbb_84_82 bitb_84_82 gnd C_bl
Rb_84_83 bit_84_83 bit_84_84 R_bl
Rbb_84_83 bitb_84_83 bitb_84_84 R_bl
Cb_84_83 bit_84_83 gnd C_bl
Cbb_84_83 bitb_84_83 gnd C_bl
Rb_84_84 bit_84_84 bit_84_85 R_bl
Rbb_84_84 bitb_84_84 bitb_84_85 R_bl
Cb_84_84 bit_84_84 gnd C_bl
Cbb_84_84 bitb_84_84 gnd C_bl
Rb_84_85 bit_84_85 bit_84_86 R_bl
Rbb_84_85 bitb_84_85 bitb_84_86 R_bl
Cb_84_85 bit_84_85 gnd C_bl
Cbb_84_85 bitb_84_85 gnd C_bl
Rb_84_86 bit_84_86 bit_84_87 R_bl
Rbb_84_86 bitb_84_86 bitb_84_87 R_bl
Cb_84_86 bit_84_86 gnd C_bl
Cbb_84_86 bitb_84_86 gnd C_bl
Rb_84_87 bit_84_87 bit_84_88 R_bl
Rbb_84_87 bitb_84_87 bitb_84_88 R_bl
Cb_84_87 bit_84_87 gnd C_bl
Cbb_84_87 bitb_84_87 gnd C_bl
Rb_84_88 bit_84_88 bit_84_89 R_bl
Rbb_84_88 bitb_84_88 bitb_84_89 R_bl
Cb_84_88 bit_84_88 gnd C_bl
Cbb_84_88 bitb_84_88 gnd C_bl
Rb_84_89 bit_84_89 bit_84_90 R_bl
Rbb_84_89 bitb_84_89 bitb_84_90 R_bl
Cb_84_89 bit_84_89 gnd C_bl
Cbb_84_89 bitb_84_89 gnd C_bl
Rb_84_90 bit_84_90 bit_84_91 R_bl
Rbb_84_90 bitb_84_90 bitb_84_91 R_bl
Cb_84_90 bit_84_90 gnd C_bl
Cbb_84_90 bitb_84_90 gnd C_bl
Rb_84_91 bit_84_91 bit_84_92 R_bl
Rbb_84_91 bitb_84_91 bitb_84_92 R_bl
Cb_84_91 bit_84_91 gnd C_bl
Cbb_84_91 bitb_84_91 gnd C_bl
Rb_84_92 bit_84_92 bit_84_93 R_bl
Rbb_84_92 bitb_84_92 bitb_84_93 R_bl
Cb_84_92 bit_84_92 gnd C_bl
Cbb_84_92 bitb_84_92 gnd C_bl
Rb_84_93 bit_84_93 bit_84_94 R_bl
Rbb_84_93 bitb_84_93 bitb_84_94 R_bl
Cb_84_93 bit_84_93 gnd C_bl
Cbb_84_93 bitb_84_93 gnd C_bl
Rb_84_94 bit_84_94 bit_84_95 R_bl
Rbb_84_94 bitb_84_94 bitb_84_95 R_bl
Cb_84_94 bit_84_94 gnd C_bl
Cbb_84_94 bitb_84_94 gnd C_bl
Rb_84_95 bit_84_95 bit_84_96 R_bl
Rbb_84_95 bitb_84_95 bitb_84_96 R_bl
Cb_84_95 bit_84_95 gnd C_bl
Cbb_84_95 bitb_84_95 gnd C_bl
Rb_84_96 bit_84_96 bit_84_97 R_bl
Rbb_84_96 bitb_84_96 bitb_84_97 R_bl
Cb_84_96 bit_84_96 gnd C_bl
Cbb_84_96 bitb_84_96 gnd C_bl
Rb_84_97 bit_84_97 bit_84_98 R_bl
Rbb_84_97 bitb_84_97 bitb_84_98 R_bl
Cb_84_97 bit_84_97 gnd C_bl
Cbb_84_97 bitb_84_97 gnd C_bl
Rb_84_98 bit_84_98 bit_84_99 R_bl
Rbb_84_98 bitb_84_98 bitb_84_99 R_bl
Cb_84_98 bit_84_98 gnd C_bl
Cbb_84_98 bitb_84_98 gnd C_bl
Rb_84_99 bit_84_99 bit_84_100 R_bl
Rbb_84_99 bitb_84_99 bitb_84_100 R_bl
Cb_84_99 bit_84_99 gnd C_bl
Cbb_84_99 bitb_84_99 gnd C_bl
Rb_85_0 bit_85_0 bit_85_1 R_bl
Rbb_85_0 bitb_85_0 bitb_85_1 R_bl
Cb_85_0 bit_85_0 gnd C_bl
Cbb_85_0 bitb_85_0 gnd C_bl
Rb_85_1 bit_85_1 bit_85_2 R_bl
Rbb_85_1 bitb_85_1 bitb_85_2 R_bl
Cb_85_1 bit_85_1 gnd C_bl
Cbb_85_1 bitb_85_1 gnd C_bl
Rb_85_2 bit_85_2 bit_85_3 R_bl
Rbb_85_2 bitb_85_2 bitb_85_3 R_bl
Cb_85_2 bit_85_2 gnd C_bl
Cbb_85_2 bitb_85_2 gnd C_bl
Rb_85_3 bit_85_3 bit_85_4 R_bl
Rbb_85_3 bitb_85_3 bitb_85_4 R_bl
Cb_85_3 bit_85_3 gnd C_bl
Cbb_85_3 bitb_85_3 gnd C_bl
Rb_85_4 bit_85_4 bit_85_5 R_bl
Rbb_85_4 bitb_85_4 bitb_85_5 R_bl
Cb_85_4 bit_85_4 gnd C_bl
Cbb_85_4 bitb_85_4 gnd C_bl
Rb_85_5 bit_85_5 bit_85_6 R_bl
Rbb_85_5 bitb_85_5 bitb_85_6 R_bl
Cb_85_5 bit_85_5 gnd C_bl
Cbb_85_5 bitb_85_5 gnd C_bl
Rb_85_6 bit_85_6 bit_85_7 R_bl
Rbb_85_6 bitb_85_6 bitb_85_7 R_bl
Cb_85_6 bit_85_6 gnd C_bl
Cbb_85_6 bitb_85_6 gnd C_bl
Rb_85_7 bit_85_7 bit_85_8 R_bl
Rbb_85_7 bitb_85_7 bitb_85_8 R_bl
Cb_85_7 bit_85_7 gnd C_bl
Cbb_85_7 bitb_85_7 gnd C_bl
Rb_85_8 bit_85_8 bit_85_9 R_bl
Rbb_85_8 bitb_85_8 bitb_85_9 R_bl
Cb_85_8 bit_85_8 gnd C_bl
Cbb_85_8 bitb_85_8 gnd C_bl
Rb_85_9 bit_85_9 bit_85_10 R_bl
Rbb_85_9 bitb_85_9 bitb_85_10 R_bl
Cb_85_9 bit_85_9 gnd C_bl
Cbb_85_9 bitb_85_9 gnd C_bl
Rb_85_10 bit_85_10 bit_85_11 R_bl
Rbb_85_10 bitb_85_10 bitb_85_11 R_bl
Cb_85_10 bit_85_10 gnd C_bl
Cbb_85_10 bitb_85_10 gnd C_bl
Rb_85_11 bit_85_11 bit_85_12 R_bl
Rbb_85_11 bitb_85_11 bitb_85_12 R_bl
Cb_85_11 bit_85_11 gnd C_bl
Cbb_85_11 bitb_85_11 gnd C_bl
Rb_85_12 bit_85_12 bit_85_13 R_bl
Rbb_85_12 bitb_85_12 bitb_85_13 R_bl
Cb_85_12 bit_85_12 gnd C_bl
Cbb_85_12 bitb_85_12 gnd C_bl
Rb_85_13 bit_85_13 bit_85_14 R_bl
Rbb_85_13 bitb_85_13 bitb_85_14 R_bl
Cb_85_13 bit_85_13 gnd C_bl
Cbb_85_13 bitb_85_13 gnd C_bl
Rb_85_14 bit_85_14 bit_85_15 R_bl
Rbb_85_14 bitb_85_14 bitb_85_15 R_bl
Cb_85_14 bit_85_14 gnd C_bl
Cbb_85_14 bitb_85_14 gnd C_bl
Rb_85_15 bit_85_15 bit_85_16 R_bl
Rbb_85_15 bitb_85_15 bitb_85_16 R_bl
Cb_85_15 bit_85_15 gnd C_bl
Cbb_85_15 bitb_85_15 gnd C_bl
Rb_85_16 bit_85_16 bit_85_17 R_bl
Rbb_85_16 bitb_85_16 bitb_85_17 R_bl
Cb_85_16 bit_85_16 gnd C_bl
Cbb_85_16 bitb_85_16 gnd C_bl
Rb_85_17 bit_85_17 bit_85_18 R_bl
Rbb_85_17 bitb_85_17 bitb_85_18 R_bl
Cb_85_17 bit_85_17 gnd C_bl
Cbb_85_17 bitb_85_17 gnd C_bl
Rb_85_18 bit_85_18 bit_85_19 R_bl
Rbb_85_18 bitb_85_18 bitb_85_19 R_bl
Cb_85_18 bit_85_18 gnd C_bl
Cbb_85_18 bitb_85_18 gnd C_bl
Rb_85_19 bit_85_19 bit_85_20 R_bl
Rbb_85_19 bitb_85_19 bitb_85_20 R_bl
Cb_85_19 bit_85_19 gnd C_bl
Cbb_85_19 bitb_85_19 gnd C_bl
Rb_85_20 bit_85_20 bit_85_21 R_bl
Rbb_85_20 bitb_85_20 bitb_85_21 R_bl
Cb_85_20 bit_85_20 gnd C_bl
Cbb_85_20 bitb_85_20 gnd C_bl
Rb_85_21 bit_85_21 bit_85_22 R_bl
Rbb_85_21 bitb_85_21 bitb_85_22 R_bl
Cb_85_21 bit_85_21 gnd C_bl
Cbb_85_21 bitb_85_21 gnd C_bl
Rb_85_22 bit_85_22 bit_85_23 R_bl
Rbb_85_22 bitb_85_22 bitb_85_23 R_bl
Cb_85_22 bit_85_22 gnd C_bl
Cbb_85_22 bitb_85_22 gnd C_bl
Rb_85_23 bit_85_23 bit_85_24 R_bl
Rbb_85_23 bitb_85_23 bitb_85_24 R_bl
Cb_85_23 bit_85_23 gnd C_bl
Cbb_85_23 bitb_85_23 gnd C_bl
Rb_85_24 bit_85_24 bit_85_25 R_bl
Rbb_85_24 bitb_85_24 bitb_85_25 R_bl
Cb_85_24 bit_85_24 gnd C_bl
Cbb_85_24 bitb_85_24 gnd C_bl
Rb_85_25 bit_85_25 bit_85_26 R_bl
Rbb_85_25 bitb_85_25 bitb_85_26 R_bl
Cb_85_25 bit_85_25 gnd C_bl
Cbb_85_25 bitb_85_25 gnd C_bl
Rb_85_26 bit_85_26 bit_85_27 R_bl
Rbb_85_26 bitb_85_26 bitb_85_27 R_bl
Cb_85_26 bit_85_26 gnd C_bl
Cbb_85_26 bitb_85_26 gnd C_bl
Rb_85_27 bit_85_27 bit_85_28 R_bl
Rbb_85_27 bitb_85_27 bitb_85_28 R_bl
Cb_85_27 bit_85_27 gnd C_bl
Cbb_85_27 bitb_85_27 gnd C_bl
Rb_85_28 bit_85_28 bit_85_29 R_bl
Rbb_85_28 bitb_85_28 bitb_85_29 R_bl
Cb_85_28 bit_85_28 gnd C_bl
Cbb_85_28 bitb_85_28 gnd C_bl
Rb_85_29 bit_85_29 bit_85_30 R_bl
Rbb_85_29 bitb_85_29 bitb_85_30 R_bl
Cb_85_29 bit_85_29 gnd C_bl
Cbb_85_29 bitb_85_29 gnd C_bl
Rb_85_30 bit_85_30 bit_85_31 R_bl
Rbb_85_30 bitb_85_30 bitb_85_31 R_bl
Cb_85_30 bit_85_30 gnd C_bl
Cbb_85_30 bitb_85_30 gnd C_bl
Rb_85_31 bit_85_31 bit_85_32 R_bl
Rbb_85_31 bitb_85_31 bitb_85_32 R_bl
Cb_85_31 bit_85_31 gnd C_bl
Cbb_85_31 bitb_85_31 gnd C_bl
Rb_85_32 bit_85_32 bit_85_33 R_bl
Rbb_85_32 bitb_85_32 bitb_85_33 R_bl
Cb_85_32 bit_85_32 gnd C_bl
Cbb_85_32 bitb_85_32 gnd C_bl
Rb_85_33 bit_85_33 bit_85_34 R_bl
Rbb_85_33 bitb_85_33 bitb_85_34 R_bl
Cb_85_33 bit_85_33 gnd C_bl
Cbb_85_33 bitb_85_33 gnd C_bl
Rb_85_34 bit_85_34 bit_85_35 R_bl
Rbb_85_34 bitb_85_34 bitb_85_35 R_bl
Cb_85_34 bit_85_34 gnd C_bl
Cbb_85_34 bitb_85_34 gnd C_bl
Rb_85_35 bit_85_35 bit_85_36 R_bl
Rbb_85_35 bitb_85_35 bitb_85_36 R_bl
Cb_85_35 bit_85_35 gnd C_bl
Cbb_85_35 bitb_85_35 gnd C_bl
Rb_85_36 bit_85_36 bit_85_37 R_bl
Rbb_85_36 bitb_85_36 bitb_85_37 R_bl
Cb_85_36 bit_85_36 gnd C_bl
Cbb_85_36 bitb_85_36 gnd C_bl
Rb_85_37 bit_85_37 bit_85_38 R_bl
Rbb_85_37 bitb_85_37 bitb_85_38 R_bl
Cb_85_37 bit_85_37 gnd C_bl
Cbb_85_37 bitb_85_37 gnd C_bl
Rb_85_38 bit_85_38 bit_85_39 R_bl
Rbb_85_38 bitb_85_38 bitb_85_39 R_bl
Cb_85_38 bit_85_38 gnd C_bl
Cbb_85_38 bitb_85_38 gnd C_bl
Rb_85_39 bit_85_39 bit_85_40 R_bl
Rbb_85_39 bitb_85_39 bitb_85_40 R_bl
Cb_85_39 bit_85_39 gnd C_bl
Cbb_85_39 bitb_85_39 gnd C_bl
Rb_85_40 bit_85_40 bit_85_41 R_bl
Rbb_85_40 bitb_85_40 bitb_85_41 R_bl
Cb_85_40 bit_85_40 gnd C_bl
Cbb_85_40 bitb_85_40 gnd C_bl
Rb_85_41 bit_85_41 bit_85_42 R_bl
Rbb_85_41 bitb_85_41 bitb_85_42 R_bl
Cb_85_41 bit_85_41 gnd C_bl
Cbb_85_41 bitb_85_41 gnd C_bl
Rb_85_42 bit_85_42 bit_85_43 R_bl
Rbb_85_42 bitb_85_42 bitb_85_43 R_bl
Cb_85_42 bit_85_42 gnd C_bl
Cbb_85_42 bitb_85_42 gnd C_bl
Rb_85_43 bit_85_43 bit_85_44 R_bl
Rbb_85_43 bitb_85_43 bitb_85_44 R_bl
Cb_85_43 bit_85_43 gnd C_bl
Cbb_85_43 bitb_85_43 gnd C_bl
Rb_85_44 bit_85_44 bit_85_45 R_bl
Rbb_85_44 bitb_85_44 bitb_85_45 R_bl
Cb_85_44 bit_85_44 gnd C_bl
Cbb_85_44 bitb_85_44 gnd C_bl
Rb_85_45 bit_85_45 bit_85_46 R_bl
Rbb_85_45 bitb_85_45 bitb_85_46 R_bl
Cb_85_45 bit_85_45 gnd C_bl
Cbb_85_45 bitb_85_45 gnd C_bl
Rb_85_46 bit_85_46 bit_85_47 R_bl
Rbb_85_46 bitb_85_46 bitb_85_47 R_bl
Cb_85_46 bit_85_46 gnd C_bl
Cbb_85_46 bitb_85_46 gnd C_bl
Rb_85_47 bit_85_47 bit_85_48 R_bl
Rbb_85_47 bitb_85_47 bitb_85_48 R_bl
Cb_85_47 bit_85_47 gnd C_bl
Cbb_85_47 bitb_85_47 gnd C_bl
Rb_85_48 bit_85_48 bit_85_49 R_bl
Rbb_85_48 bitb_85_48 bitb_85_49 R_bl
Cb_85_48 bit_85_48 gnd C_bl
Cbb_85_48 bitb_85_48 gnd C_bl
Rb_85_49 bit_85_49 bit_85_50 R_bl
Rbb_85_49 bitb_85_49 bitb_85_50 R_bl
Cb_85_49 bit_85_49 gnd C_bl
Cbb_85_49 bitb_85_49 gnd C_bl
Rb_85_50 bit_85_50 bit_85_51 R_bl
Rbb_85_50 bitb_85_50 bitb_85_51 R_bl
Cb_85_50 bit_85_50 gnd C_bl
Cbb_85_50 bitb_85_50 gnd C_bl
Rb_85_51 bit_85_51 bit_85_52 R_bl
Rbb_85_51 bitb_85_51 bitb_85_52 R_bl
Cb_85_51 bit_85_51 gnd C_bl
Cbb_85_51 bitb_85_51 gnd C_bl
Rb_85_52 bit_85_52 bit_85_53 R_bl
Rbb_85_52 bitb_85_52 bitb_85_53 R_bl
Cb_85_52 bit_85_52 gnd C_bl
Cbb_85_52 bitb_85_52 gnd C_bl
Rb_85_53 bit_85_53 bit_85_54 R_bl
Rbb_85_53 bitb_85_53 bitb_85_54 R_bl
Cb_85_53 bit_85_53 gnd C_bl
Cbb_85_53 bitb_85_53 gnd C_bl
Rb_85_54 bit_85_54 bit_85_55 R_bl
Rbb_85_54 bitb_85_54 bitb_85_55 R_bl
Cb_85_54 bit_85_54 gnd C_bl
Cbb_85_54 bitb_85_54 gnd C_bl
Rb_85_55 bit_85_55 bit_85_56 R_bl
Rbb_85_55 bitb_85_55 bitb_85_56 R_bl
Cb_85_55 bit_85_55 gnd C_bl
Cbb_85_55 bitb_85_55 gnd C_bl
Rb_85_56 bit_85_56 bit_85_57 R_bl
Rbb_85_56 bitb_85_56 bitb_85_57 R_bl
Cb_85_56 bit_85_56 gnd C_bl
Cbb_85_56 bitb_85_56 gnd C_bl
Rb_85_57 bit_85_57 bit_85_58 R_bl
Rbb_85_57 bitb_85_57 bitb_85_58 R_bl
Cb_85_57 bit_85_57 gnd C_bl
Cbb_85_57 bitb_85_57 gnd C_bl
Rb_85_58 bit_85_58 bit_85_59 R_bl
Rbb_85_58 bitb_85_58 bitb_85_59 R_bl
Cb_85_58 bit_85_58 gnd C_bl
Cbb_85_58 bitb_85_58 gnd C_bl
Rb_85_59 bit_85_59 bit_85_60 R_bl
Rbb_85_59 bitb_85_59 bitb_85_60 R_bl
Cb_85_59 bit_85_59 gnd C_bl
Cbb_85_59 bitb_85_59 gnd C_bl
Rb_85_60 bit_85_60 bit_85_61 R_bl
Rbb_85_60 bitb_85_60 bitb_85_61 R_bl
Cb_85_60 bit_85_60 gnd C_bl
Cbb_85_60 bitb_85_60 gnd C_bl
Rb_85_61 bit_85_61 bit_85_62 R_bl
Rbb_85_61 bitb_85_61 bitb_85_62 R_bl
Cb_85_61 bit_85_61 gnd C_bl
Cbb_85_61 bitb_85_61 gnd C_bl
Rb_85_62 bit_85_62 bit_85_63 R_bl
Rbb_85_62 bitb_85_62 bitb_85_63 R_bl
Cb_85_62 bit_85_62 gnd C_bl
Cbb_85_62 bitb_85_62 gnd C_bl
Rb_85_63 bit_85_63 bit_85_64 R_bl
Rbb_85_63 bitb_85_63 bitb_85_64 R_bl
Cb_85_63 bit_85_63 gnd C_bl
Cbb_85_63 bitb_85_63 gnd C_bl
Rb_85_64 bit_85_64 bit_85_65 R_bl
Rbb_85_64 bitb_85_64 bitb_85_65 R_bl
Cb_85_64 bit_85_64 gnd C_bl
Cbb_85_64 bitb_85_64 gnd C_bl
Rb_85_65 bit_85_65 bit_85_66 R_bl
Rbb_85_65 bitb_85_65 bitb_85_66 R_bl
Cb_85_65 bit_85_65 gnd C_bl
Cbb_85_65 bitb_85_65 gnd C_bl
Rb_85_66 bit_85_66 bit_85_67 R_bl
Rbb_85_66 bitb_85_66 bitb_85_67 R_bl
Cb_85_66 bit_85_66 gnd C_bl
Cbb_85_66 bitb_85_66 gnd C_bl
Rb_85_67 bit_85_67 bit_85_68 R_bl
Rbb_85_67 bitb_85_67 bitb_85_68 R_bl
Cb_85_67 bit_85_67 gnd C_bl
Cbb_85_67 bitb_85_67 gnd C_bl
Rb_85_68 bit_85_68 bit_85_69 R_bl
Rbb_85_68 bitb_85_68 bitb_85_69 R_bl
Cb_85_68 bit_85_68 gnd C_bl
Cbb_85_68 bitb_85_68 gnd C_bl
Rb_85_69 bit_85_69 bit_85_70 R_bl
Rbb_85_69 bitb_85_69 bitb_85_70 R_bl
Cb_85_69 bit_85_69 gnd C_bl
Cbb_85_69 bitb_85_69 gnd C_bl
Rb_85_70 bit_85_70 bit_85_71 R_bl
Rbb_85_70 bitb_85_70 bitb_85_71 R_bl
Cb_85_70 bit_85_70 gnd C_bl
Cbb_85_70 bitb_85_70 gnd C_bl
Rb_85_71 bit_85_71 bit_85_72 R_bl
Rbb_85_71 bitb_85_71 bitb_85_72 R_bl
Cb_85_71 bit_85_71 gnd C_bl
Cbb_85_71 bitb_85_71 gnd C_bl
Rb_85_72 bit_85_72 bit_85_73 R_bl
Rbb_85_72 bitb_85_72 bitb_85_73 R_bl
Cb_85_72 bit_85_72 gnd C_bl
Cbb_85_72 bitb_85_72 gnd C_bl
Rb_85_73 bit_85_73 bit_85_74 R_bl
Rbb_85_73 bitb_85_73 bitb_85_74 R_bl
Cb_85_73 bit_85_73 gnd C_bl
Cbb_85_73 bitb_85_73 gnd C_bl
Rb_85_74 bit_85_74 bit_85_75 R_bl
Rbb_85_74 bitb_85_74 bitb_85_75 R_bl
Cb_85_74 bit_85_74 gnd C_bl
Cbb_85_74 bitb_85_74 gnd C_bl
Rb_85_75 bit_85_75 bit_85_76 R_bl
Rbb_85_75 bitb_85_75 bitb_85_76 R_bl
Cb_85_75 bit_85_75 gnd C_bl
Cbb_85_75 bitb_85_75 gnd C_bl
Rb_85_76 bit_85_76 bit_85_77 R_bl
Rbb_85_76 bitb_85_76 bitb_85_77 R_bl
Cb_85_76 bit_85_76 gnd C_bl
Cbb_85_76 bitb_85_76 gnd C_bl
Rb_85_77 bit_85_77 bit_85_78 R_bl
Rbb_85_77 bitb_85_77 bitb_85_78 R_bl
Cb_85_77 bit_85_77 gnd C_bl
Cbb_85_77 bitb_85_77 gnd C_bl
Rb_85_78 bit_85_78 bit_85_79 R_bl
Rbb_85_78 bitb_85_78 bitb_85_79 R_bl
Cb_85_78 bit_85_78 gnd C_bl
Cbb_85_78 bitb_85_78 gnd C_bl
Rb_85_79 bit_85_79 bit_85_80 R_bl
Rbb_85_79 bitb_85_79 bitb_85_80 R_bl
Cb_85_79 bit_85_79 gnd C_bl
Cbb_85_79 bitb_85_79 gnd C_bl
Rb_85_80 bit_85_80 bit_85_81 R_bl
Rbb_85_80 bitb_85_80 bitb_85_81 R_bl
Cb_85_80 bit_85_80 gnd C_bl
Cbb_85_80 bitb_85_80 gnd C_bl
Rb_85_81 bit_85_81 bit_85_82 R_bl
Rbb_85_81 bitb_85_81 bitb_85_82 R_bl
Cb_85_81 bit_85_81 gnd C_bl
Cbb_85_81 bitb_85_81 gnd C_bl
Rb_85_82 bit_85_82 bit_85_83 R_bl
Rbb_85_82 bitb_85_82 bitb_85_83 R_bl
Cb_85_82 bit_85_82 gnd C_bl
Cbb_85_82 bitb_85_82 gnd C_bl
Rb_85_83 bit_85_83 bit_85_84 R_bl
Rbb_85_83 bitb_85_83 bitb_85_84 R_bl
Cb_85_83 bit_85_83 gnd C_bl
Cbb_85_83 bitb_85_83 gnd C_bl
Rb_85_84 bit_85_84 bit_85_85 R_bl
Rbb_85_84 bitb_85_84 bitb_85_85 R_bl
Cb_85_84 bit_85_84 gnd C_bl
Cbb_85_84 bitb_85_84 gnd C_bl
Rb_85_85 bit_85_85 bit_85_86 R_bl
Rbb_85_85 bitb_85_85 bitb_85_86 R_bl
Cb_85_85 bit_85_85 gnd C_bl
Cbb_85_85 bitb_85_85 gnd C_bl
Rb_85_86 bit_85_86 bit_85_87 R_bl
Rbb_85_86 bitb_85_86 bitb_85_87 R_bl
Cb_85_86 bit_85_86 gnd C_bl
Cbb_85_86 bitb_85_86 gnd C_bl
Rb_85_87 bit_85_87 bit_85_88 R_bl
Rbb_85_87 bitb_85_87 bitb_85_88 R_bl
Cb_85_87 bit_85_87 gnd C_bl
Cbb_85_87 bitb_85_87 gnd C_bl
Rb_85_88 bit_85_88 bit_85_89 R_bl
Rbb_85_88 bitb_85_88 bitb_85_89 R_bl
Cb_85_88 bit_85_88 gnd C_bl
Cbb_85_88 bitb_85_88 gnd C_bl
Rb_85_89 bit_85_89 bit_85_90 R_bl
Rbb_85_89 bitb_85_89 bitb_85_90 R_bl
Cb_85_89 bit_85_89 gnd C_bl
Cbb_85_89 bitb_85_89 gnd C_bl
Rb_85_90 bit_85_90 bit_85_91 R_bl
Rbb_85_90 bitb_85_90 bitb_85_91 R_bl
Cb_85_90 bit_85_90 gnd C_bl
Cbb_85_90 bitb_85_90 gnd C_bl
Rb_85_91 bit_85_91 bit_85_92 R_bl
Rbb_85_91 bitb_85_91 bitb_85_92 R_bl
Cb_85_91 bit_85_91 gnd C_bl
Cbb_85_91 bitb_85_91 gnd C_bl
Rb_85_92 bit_85_92 bit_85_93 R_bl
Rbb_85_92 bitb_85_92 bitb_85_93 R_bl
Cb_85_92 bit_85_92 gnd C_bl
Cbb_85_92 bitb_85_92 gnd C_bl
Rb_85_93 bit_85_93 bit_85_94 R_bl
Rbb_85_93 bitb_85_93 bitb_85_94 R_bl
Cb_85_93 bit_85_93 gnd C_bl
Cbb_85_93 bitb_85_93 gnd C_bl
Rb_85_94 bit_85_94 bit_85_95 R_bl
Rbb_85_94 bitb_85_94 bitb_85_95 R_bl
Cb_85_94 bit_85_94 gnd C_bl
Cbb_85_94 bitb_85_94 gnd C_bl
Rb_85_95 bit_85_95 bit_85_96 R_bl
Rbb_85_95 bitb_85_95 bitb_85_96 R_bl
Cb_85_95 bit_85_95 gnd C_bl
Cbb_85_95 bitb_85_95 gnd C_bl
Rb_85_96 bit_85_96 bit_85_97 R_bl
Rbb_85_96 bitb_85_96 bitb_85_97 R_bl
Cb_85_96 bit_85_96 gnd C_bl
Cbb_85_96 bitb_85_96 gnd C_bl
Rb_85_97 bit_85_97 bit_85_98 R_bl
Rbb_85_97 bitb_85_97 bitb_85_98 R_bl
Cb_85_97 bit_85_97 gnd C_bl
Cbb_85_97 bitb_85_97 gnd C_bl
Rb_85_98 bit_85_98 bit_85_99 R_bl
Rbb_85_98 bitb_85_98 bitb_85_99 R_bl
Cb_85_98 bit_85_98 gnd C_bl
Cbb_85_98 bitb_85_98 gnd C_bl
Rb_85_99 bit_85_99 bit_85_100 R_bl
Rbb_85_99 bitb_85_99 bitb_85_100 R_bl
Cb_85_99 bit_85_99 gnd C_bl
Cbb_85_99 bitb_85_99 gnd C_bl
Rb_86_0 bit_86_0 bit_86_1 R_bl
Rbb_86_0 bitb_86_0 bitb_86_1 R_bl
Cb_86_0 bit_86_0 gnd C_bl
Cbb_86_0 bitb_86_0 gnd C_bl
Rb_86_1 bit_86_1 bit_86_2 R_bl
Rbb_86_1 bitb_86_1 bitb_86_2 R_bl
Cb_86_1 bit_86_1 gnd C_bl
Cbb_86_1 bitb_86_1 gnd C_bl
Rb_86_2 bit_86_2 bit_86_3 R_bl
Rbb_86_2 bitb_86_2 bitb_86_3 R_bl
Cb_86_2 bit_86_2 gnd C_bl
Cbb_86_2 bitb_86_2 gnd C_bl
Rb_86_3 bit_86_3 bit_86_4 R_bl
Rbb_86_3 bitb_86_3 bitb_86_4 R_bl
Cb_86_3 bit_86_3 gnd C_bl
Cbb_86_3 bitb_86_3 gnd C_bl
Rb_86_4 bit_86_4 bit_86_5 R_bl
Rbb_86_4 bitb_86_4 bitb_86_5 R_bl
Cb_86_4 bit_86_4 gnd C_bl
Cbb_86_4 bitb_86_4 gnd C_bl
Rb_86_5 bit_86_5 bit_86_6 R_bl
Rbb_86_5 bitb_86_5 bitb_86_6 R_bl
Cb_86_5 bit_86_5 gnd C_bl
Cbb_86_5 bitb_86_5 gnd C_bl
Rb_86_6 bit_86_6 bit_86_7 R_bl
Rbb_86_6 bitb_86_6 bitb_86_7 R_bl
Cb_86_6 bit_86_6 gnd C_bl
Cbb_86_6 bitb_86_6 gnd C_bl
Rb_86_7 bit_86_7 bit_86_8 R_bl
Rbb_86_7 bitb_86_7 bitb_86_8 R_bl
Cb_86_7 bit_86_7 gnd C_bl
Cbb_86_7 bitb_86_7 gnd C_bl
Rb_86_8 bit_86_8 bit_86_9 R_bl
Rbb_86_8 bitb_86_8 bitb_86_9 R_bl
Cb_86_8 bit_86_8 gnd C_bl
Cbb_86_8 bitb_86_8 gnd C_bl
Rb_86_9 bit_86_9 bit_86_10 R_bl
Rbb_86_9 bitb_86_9 bitb_86_10 R_bl
Cb_86_9 bit_86_9 gnd C_bl
Cbb_86_9 bitb_86_9 gnd C_bl
Rb_86_10 bit_86_10 bit_86_11 R_bl
Rbb_86_10 bitb_86_10 bitb_86_11 R_bl
Cb_86_10 bit_86_10 gnd C_bl
Cbb_86_10 bitb_86_10 gnd C_bl
Rb_86_11 bit_86_11 bit_86_12 R_bl
Rbb_86_11 bitb_86_11 bitb_86_12 R_bl
Cb_86_11 bit_86_11 gnd C_bl
Cbb_86_11 bitb_86_11 gnd C_bl
Rb_86_12 bit_86_12 bit_86_13 R_bl
Rbb_86_12 bitb_86_12 bitb_86_13 R_bl
Cb_86_12 bit_86_12 gnd C_bl
Cbb_86_12 bitb_86_12 gnd C_bl
Rb_86_13 bit_86_13 bit_86_14 R_bl
Rbb_86_13 bitb_86_13 bitb_86_14 R_bl
Cb_86_13 bit_86_13 gnd C_bl
Cbb_86_13 bitb_86_13 gnd C_bl
Rb_86_14 bit_86_14 bit_86_15 R_bl
Rbb_86_14 bitb_86_14 bitb_86_15 R_bl
Cb_86_14 bit_86_14 gnd C_bl
Cbb_86_14 bitb_86_14 gnd C_bl
Rb_86_15 bit_86_15 bit_86_16 R_bl
Rbb_86_15 bitb_86_15 bitb_86_16 R_bl
Cb_86_15 bit_86_15 gnd C_bl
Cbb_86_15 bitb_86_15 gnd C_bl
Rb_86_16 bit_86_16 bit_86_17 R_bl
Rbb_86_16 bitb_86_16 bitb_86_17 R_bl
Cb_86_16 bit_86_16 gnd C_bl
Cbb_86_16 bitb_86_16 gnd C_bl
Rb_86_17 bit_86_17 bit_86_18 R_bl
Rbb_86_17 bitb_86_17 bitb_86_18 R_bl
Cb_86_17 bit_86_17 gnd C_bl
Cbb_86_17 bitb_86_17 gnd C_bl
Rb_86_18 bit_86_18 bit_86_19 R_bl
Rbb_86_18 bitb_86_18 bitb_86_19 R_bl
Cb_86_18 bit_86_18 gnd C_bl
Cbb_86_18 bitb_86_18 gnd C_bl
Rb_86_19 bit_86_19 bit_86_20 R_bl
Rbb_86_19 bitb_86_19 bitb_86_20 R_bl
Cb_86_19 bit_86_19 gnd C_bl
Cbb_86_19 bitb_86_19 gnd C_bl
Rb_86_20 bit_86_20 bit_86_21 R_bl
Rbb_86_20 bitb_86_20 bitb_86_21 R_bl
Cb_86_20 bit_86_20 gnd C_bl
Cbb_86_20 bitb_86_20 gnd C_bl
Rb_86_21 bit_86_21 bit_86_22 R_bl
Rbb_86_21 bitb_86_21 bitb_86_22 R_bl
Cb_86_21 bit_86_21 gnd C_bl
Cbb_86_21 bitb_86_21 gnd C_bl
Rb_86_22 bit_86_22 bit_86_23 R_bl
Rbb_86_22 bitb_86_22 bitb_86_23 R_bl
Cb_86_22 bit_86_22 gnd C_bl
Cbb_86_22 bitb_86_22 gnd C_bl
Rb_86_23 bit_86_23 bit_86_24 R_bl
Rbb_86_23 bitb_86_23 bitb_86_24 R_bl
Cb_86_23 bit_86_23 gnd C_bl
Cbb_86_23 bitb_86_23 gnd C_bl
Rb_86_24 bit_86_24 bit_86_25 R_bl
Rbb_86_24 bitb_86_24 bitb_86_25 R_bl
Cb_86_24 bit_86_24 gnd C_bl
Cbb_86_24 bitb_86_24 gnd C_bl
Rb_86_25 bit_86_25 bit_86_26 R_bl
Rbb_86_25 bitb_86_25 bitb_86_26 R_bl
Cb_86_25 bit_86_25 gnd C_bl
Cbb_86_25 bitb_86_25 gnd C_bl
Rb_86_26 bit_86_26 bit_86_27 R_bl
Rbb_86_26 bitb_86_26 bitb_86_27 R_bl
Cb_86_26 bit_86_26 gnd C_bl
Cbb_86_26 bitb_86_26 gnd C_bl
Rb_86_27 bit_86_27 bit_86_28 R_bl
Rbb_86_27 bitb_86_27 bitb_86_28 R_bl
Cb_86_27 bit_86_27 gnd C_bl
Cbb_86_27 bitb_86_27 gnd C_bl
Rb_86_28 bit_86_28 bit_86_29 R_bl
Rbb_86_28 bitb_86_28 bitb_86_29 R_bl
Cb_86_28 bit_86_28 gnd C_bl
Cbb_86_28 bitb_86_28 gnd C_bl
Rb_86_29 bit_86_29 bit_86_30 R_bl
Rbb_86_29 bitb_86_29 bitb_86_30 R_bl
Cb_86_29 bit_86_29 gnd C_bl
Cbb_86_29 bitb_86_29 gnd C_bl
Rb_86_30 bit_86_30 bit_86_31 R_bl
Rbb_86_30 bitb_86_30 bitb_86_31 R_bl
Cb_86_30 bit_86_30 gnd C_bl
Cbb_86_30 bitb_86_30 gnd C_bl
Rb_86_31 bit_86_31 bit_86_32 R_bl
Rbb_86_31 bitb_86_31 bitb_86_32 R_bl
Cb_86_31 bit_86_31 gnd C_bl
Cbb_86_31 bitb_86_31 gnd C_bl
Rb_86_32 bit_86_32 bit_86_33 R_bl
Rbb_86_32 bitb_86_32 bitb_86_33 R_bl
Cb_86_32 bit_86_32 gnd C_bl
Cbb_86_32 bitb_86_32 gnd C_bl
Rb_86_33 bit_86_33 bit_86_34 R_bl
Rbb_86_33 bitb_86_33 bitb_86_34 R_bl
Cb_86_33 bit_86_33 gnd C_bl
Cbb_86_33 bitb_86_33 gnd C_bl
Rb_86_34 bit_86_34 bit_86_35 R_bl
Rbb_86_34 bitb_86_34 bitb_86_35 R_bl
Cb_86_34 bit_86_34 gnd C_bl
Cbb_86_34 bitb_86_34 gnd C_bl
Rb_86_35 bit_86_35 bit_86_36 R_bl
Rbb_86_35 bitb_86_35 bitb_86_36 R_bl
Cb_86_35 bit_86_35 gnd C_bl
Cbb_86_35 bitb_86_35 gnd C_bl
Rb_86_36 bit_86_36 bit_86_37 R_bl
Rbb_86_36 bitb_86_36 bitb_86_37 R_bl
Cb_86_36 bit_86_36 gnd C_bl
Cbb_86_36 bitb_86_36 gnd C_bl
Rb_86_37 bit_86_37 bit_86_38 R_bl
Rbb_86_37 bitb_86_37 bitb_86_38 R_bl
Cb_86_37 bit_86_37 gnd C_bl
Cbb_86_37 bitb_86_37 gnd C_bl
Rb_86_38 bit_86_38 bit_86_39 R_bl
Rbb_86_38 bitb_86_38 bitb_86_39 R_bl
Cb_86_38 bit_86_38 gnd C_bl
Cbb_86_38 bitb_86_38 gnd C_bl
Rb_86_39 bit_86_39 bit_86_40 R_bl
Rbb_86_39 bitb_86_39 bitb_86_40 R_bl
Cb_86_39 bit_86_39 gnd C_bl
Cbb_86_39 bitb_86_39 gnd C_bl
Rb_86_40 bit_86_40 bit_86_41 R_bl
Rbb_86_40 bitb_86_40 bitb_86_41 R_bl
Cb_86_40 bit_86_40 gnd C_bl
Cbb_86_40 bitb_86_40 gnd C_bl
Rb_86_41 bit_86_41 bit_86_42 R_bl
Rbb_86_41 bitb_86_41 bitb_86_42 R_bl
Cb_86_41 bit_86_41 gnd C_bl
Cbb_86_41 bitb_86_41 gnd C_bl
Rb_86_42 bit_86_42 bit_86_43 R_bl
Rbb_86_42 bitb_86_42 bitb_86_43 R_bl
Cb_86_42 bit_86_42 gnd C_bl
Cbb_86_42 bitb_86_42 gnd C_bl
Rb_86_43 bit_86_43 bit_86_44 R_bl
Rbb_86_43 bitb_86_43 bitb_86_44 R_bl
Cb_86_43 bit_86_43 gnd C_bl
Cbb_86_43 bitb_86_43 gnd C_bl
Rb_86_44 bit_86_44 bit_86_45 R_bl
Rbb_86_44 bitb_86_44 bitb_86_45 R_bl
Cb_86_44 bit_86_44 gnd C_bl
Cbb_86_44 bitb_86_44 gnd C_bl
Rb_86_45 bit_86_45 bit_86_46 R_bl
Rbb_86_45 bitb_86_45 bitb_86_46 R_bl
Cb_86_45 bit_86_45 gnd C_bl
Cbb_86_45 bitb_86_45 gnd C_bl
Rb_86_46 bit_86_46 bit_86_47 R_bl
Rbb_86_46 bitb_86_46 bitb_86_47 R_bl
Cb_86_46 bit_86_46 gnd C_bl
Cbb_86_46 bitb_86_46 gnd C_bl
Rb_86_47 bit_86_47 bit_86_48 R_bl
Rbb_86_47 bitb_86_47 bitb_86_48 R_bl
Cb_86_47 bit_86_47 gnd C_bl
Cbb_86_47 bitb_86_47 gnd C_bl
Rb_86_48 bit_86_48 bit_86_49 R_bl
Rbb_86_48 bitb_86_48 bitb_86_49 R_bl
Cb_86_48 bit_86_48 gnd C_bl
Cbb_86_48 bitb_86_48 gnd C_bl
Rb_86_49 bit_86_49 bit_86_50 R_bl
Rbb_86_49 bitb_86_49 bitb_86_50 R_bl
Cb_86_49 bit_86_49 gnd C_bl
Cbb_86_49 bitb_86_49 gnd C_bl
Rb_86_50 bit_86_50 bit_86_51 R_bl
Rbb_86_50 bitb_86_50 bitb_86_51 R_bl
Cb_86_50 bit_86_50 gnd C_bl
Cbb_86_50 bitb_86_50 gnd C_bl
Rb_86_51 bit_86_51 bit_86_52 R_bl
Rbb_86_51 bitb_86_51 bitb_86_52 R_bl
Cb_86_51 bit_86_51 gnd C_bl
Cbb_86_51 bitb_86_51 gnd C_bl
Rb_86_52 bit_86_52 bit_86_53 R_bl
Rbb_86_52 bitb_86_52 bitb_86_53 R_bl
Cb_86_52 bit_86_52 gnd C_bl
Cbb_86_52 bitb_86_52 gnd C_bl
Rb_86_53 bit_86_53 bit_86_54 R_bl
Rbb_86_53 bitb_86_53 bitb_86_54 R_bl
Cb_86_53 bit_86_53 gnd C_bl
Cbb_86_53 bitb_86_53 gnd C_bl
Rb_86_54 bit_86_54 bit_86_55 R_bl
Rbb_86_54 bitb_86_54 bitb_86_55 R_bl
Cb_86_54 bit_86_54 gnd C_bl
Cbb_86_54 bitb_86_54 gnd C_bl
Rb_86_55 bit_86_55 bit_86_56 R_bl
Rbb_86_55 bitb_86_55 bitb_86_56 R_bl
Cb_86_55 bit_86_55 gnd C_bl
Cbb_86_55 bitb_86_55 gnd C_bl
Rb_86_56 bit_86_56 bit_86_57 R_bl
Rbb_86_56 bitb_86_56 bitb_86_57 R_bl
Cb_86_56 bit_86_56 gnd C_bl
Cbb_86_56 bitb_86_56 gnd C_bl
Rb_86_57 bit_86_57 bit_86_58 R_bl
Rbb_86_57 bitb_86_57 bitb_86_58 R_bl
Cb_86_57 bit_86_57 gnd C_bl
Cbb_86_57 bitb_86_57 gnd C_bl
Rb_86_58 bit_86_58 bit_86_59 R_bl
Rbb_86_58 bitb_86_58 bitb_86_59 R_bl
Cb_86_58 bit_86_58 gnd C_bl
Cbb_86_58 bitb_86_58 gnd C_bl
Rb_86_59 bit_86_59 bit_86_60 R_bl
Rbb_86_59 bitb_86_59 bitb_86_60 R_bl
Cb_86_59 bit_86_59 gnd C_bl
Cbb_86_59 bitb_86_59 gnd C_bl
Rb_86_60 bit_86_60 bit_86_61 R_bl
Rbb_86_60 bitb_86_60 bitb_86_61 R_bl
Cb_86_60 bit_86_60 gnd C_bl
Cbb_86_60 bitb_86_60 gnd C_bl
Rb_86_61 bit_86_61 bit_86_62 R_bl
Rbb_86_61 bitb_86_61 bitb_86_62 R_bl
Cb_86_61 bit_86_61 gnd C_bl
Cbb_86_61 bitb_86_61 gnd C_bl
Rb_86_62 bit_86_62 bit_86_63 R_bl
Rbb_86_62 bitb_86_62 bitb_86_63 R_bl
Cb_86_62 bit_86_62 gnd C_bl
Cbb_86_62 bitb_86_62 gnd C_bl
Rb_86_63 bit_86_63 bit_86_64 R_bl
Rbb_86_63 bitb_86_63 bitb_86_64 R_bl
Cb_86_63 bit_86_63 gnd C_bl
Cbb_86_63 bitb_86_63 gnd C_bl
Rb_86_64 bit_86_64 bit_86_65 R_bl
Rbb_86_64 bitb_86_64 bitb_86_65 R_bl
Cb_86_64 bit_86_64 gnd C_bl
Cbb_86_64 bitb_86_64 gnd C_bl
Rb_86_65 bit_86_65 bit_86_66 R_bl
Rbb_86_65 bitb_86_65 bitb_86_66 R_bl
Cb_86_65 bit_86_65 gnd C_bl
Cbb_86_65 bitb_86_65 gnd C_bl
Rb_86_66 bit_86_66 bit_86_67 R_bl
Rbb_86_66 bitb_86_66 bitb_86_67 R_bl
Cb_86_66 bit_86_66 gnd C_bl
Cbb_86_66 bitb_86_66 gnd C_bl
Rb_86_67 bit_86_67 bit_86_68 R_bl
Rbb_86_67 bitb_86_67 bitb_86_68 R_bl
Cb_86_67 bit_86_67 gnd C_bl
Cbb_86_67 bitb_86_67 gnd C_bl
Rb_86_68 bit_86_68 bit_86_69 R_bl
Rbb_86_68 bitb_86_68 bitb_86_69 R_bl
Cb_86_68 bit_86_68 gnd C_bl
Cbb_86_68 bitb_86_68 gnd C_bl
Rb_86_69 bit_86_69 bit_86_70 R_bl
Rbb_86_69 bitb_86_69 bitb_86_70 R_bl
Cb_86_69 bit_86_69 gnd C_bl
Cbb_86_69 bitb_86_69 gnd C_bl
Rb_86_70 bit_86_70 bit_86_71 R_bl
Rbb_86_70 bitb_86_70 bitb_86_71 R_bl
Cb_86_70 bit_86_70 gnd C_bl
Cbb_86_70 bitb_86_70 gnd C_bl
Rb_86_71 bit_86_71 bit_86_72 R_bl
Rbb_86_71 bitb_86_71 bitb_86_72 R_bl
Cb_86_71 bit_86_71 gnd C_bl
Cbb_86_71 bitb_86_71 gnd C_bl
Rb_86_72 bit_86_72 bit_86_73 R_bl
Rbb_86_72 bitb_86_72 bitb_86_73 R_bl
Cb_86_72 bit_86_72 gnd C_bl
Cbb_86_72 bitb_86_72 gnd C_bl
Rb_86_73 bit_86_73 bit_86_74 R_bl
Rbb_86_73 bitb_86_73 bitb_86_74 R_bl
Cb_86_73 bit_86_73 gnd C_bl
Cbb_86_73 bitb_86_73 gnd C_bl
Rb_86_74 bit_86_74 bit_86_75 R_bl
Rbb_86_74 bitb_86_74 bitb_86_75 R_bl
Cb_86_74 bit_86_74 gnd C_bl
Cbb_86_74 bitb_86_74 gnd C_bl
Rb_86_75 bit_86_75 bit_86_76 R_bl
Rbb_86_75 bitb_86_75 bitb_86_76 R_bl
Cb_86_75 bit_86_75 gnd C_bl
Cbb_86_75 bitb_86_75 gnd C_bl
Rb_86_76 bit_86_76 bit_86_77 R_bl
Rbb_86_76 bitb_86_76 bitb_86_77 R_bl
Cb_86_76 bit_86_76 gnd C_bl
Cbb_86_76 bitb_86_76 gnd C_bl
Rb_86_77 bit_86_77 bit_86_78 R_bl
Rbb_86_77 bitb_86_77 bitb_86_78 R_bl
Cb_86_77 bit_86_77 gnd C_bl
Cbb_86_77 bitb_86_77 gnd C_bl
Rb_86_78 bit_86_78 bit_86_79 R_bl
Rbb_86_78 bitb_86_78 bitb_86_79 R_bl
Cb_86_78 bit_86_78 gnd C_bl
Cbb_86_78 bitb_86_78 gnd C_bl
Rb_86_79 bit_86_79 bit_86_80 R_bl
Rbb_86_79 bitb_86_79 bitb_86_80 R_bl
Cb_86_79 bit_86_79 gnd C_bl
Cbb_86_79 bitb_86_79 gnd C_bl
Rb_86_80 bit_86_80 bit_86_81 R_bl
Rbb_86_80 bitb_86_80 bitb_86_81 R_bl
Cb_86_80 bit_86_80 gnd C_bl
Cbb_86_80 bitb_86_80 gnd C_bl
Rb_86_81 bit_86_81 bit_86_82 R_bl
Rbb_86_81 bitb_86_81 bitb_86_82 R_bl
Cb_86_81 bit_86_81 gnd C_bl
Cbb_86_81 bitb_86_81 gnd C_bl
Rb_86_82 bit_86_82 bit_86_83 R_bl
Rbb_86_82 bitb_86_82 bitb_86_83 R_bl
Cb_86_82 bit_86_82 gnd C_bl
Cbb_86_82 bitb_86_82 gnd C_bl
Rb_86_83 bit_86_83 bit_86_84 R_bl
Rbb_86_83 bitb_86_83 bitb_86_84 R_bl
Cb_86_83 bit_86_83 gnd C_bl
Cbb_86_83 bitb_86_83 gnd C_bl
Rb_86_84 bit_86_84 bit_86_85 R_bl
Rbb_86_84 bitb_86_84 bitb_86_85 R_bl
Cb_86_84 bit_86_84 gnd C_bl
Cbb_86_84 bitb_86_84 gnd C_bl
Rb_86_85 bit_86_85 bit_86_86 R_bl
Rbb_86_85 bitb_86_85 bitb_86_86 R_bl
Cb_86_85 bit_86_85 gnd C_bl
Cbb_86_85 bitb_86_85 gnd C_bl
Rb_86_86 bit_86_86 bit_86_87 R_bl
Rbb_86_86 bitb_86_86 bitb_86_87 R_bl
Cb_86_86 bit_86_86 gnd C_bl
Cbb_86_86 bitb_86_86 gnd C_bl
Rb_86_87 bit_86_87 bit_86_88 R_bl
Rbb_86_87 bitb_86_87 bitb_86_88 R_bl
Cb_86_87 bit_86_87 gnd C_bl
Cbb_86_87 bitb_86_87 gnd C_bl
Rb_86_88 bit_86_88 bit_86_89 R_bl
Rbb_86_88 bitb_86_88 bitb_86_89 R_bl
Cb_86_88 bit_86_88 gnd C_bl
Cbb_86_88 bitb_86_88 gnd C_bl
Rb_86_89 bit_86_89 bit_86_90 R_bl
Rbb_86_89 bitb_86_89 bitb_86_90 R_bl
Cb_86_89 bit_86_89 gnd C_bl
Cbb_86_89 bitb_86_89 gnd C_bl
Rb_86_90 bit_86_90 bit_86_91 R_bl
Rbb_86_90 bitb_86_90 bitb_86_91 R_bl
Cb_86_90 bit_86_90 gnd C_bl
Cbb_86_90 bitb_86_90 gnd C_bl
Rb_86_91 bit_86_91 bit_86_92 R_bl
Rbb_86_91 bitb_86_91 bitb_86_92 R_bl
Cb_86_91 bit_86_91 gnd C_bl
Cbb_86_91 bitb_86_91 gnd C_bl
Rb_86_92 bit_86_92 bit_86_93 R_bl
Rbb_86_92 bitb_86_92 bitb_86_93 R_bl
Cb_86_92 bit_86_92 gnd C_bl
Cbb_86_92 bitb_86_92 gnd C_bl
Rb_86_93 bit_86_93 bit_86_94 R_bl
Rbb_86_93 bitb_86_93 bitb_86_94 R_bl
Cb_86_93 bit_86_93 gnd C_bl
Cbb_86_93 bitb_86_93 gnd C_bl
Rb_86_94 bit_86_94 bit_86_95 R_bl
Rbb_86_94 bitb_86_94 bitb_86_95 R_bl
Cb_86_94 bit_86_94 gnd C_bl
Cbb_86_94 bitb_86_94 gnd C_bl
Rb_86_95 bit_86_95 bit_86_96 R_bl
Rbb_86_95 bitb_86_95 bitb_86_96 R_bl
Cb_86_95 bit_86_95 gnd C_bl
Cbb_86_95 bitb_86_95 gnd C_bl
Rb_86_96 bit_86_96 bit_86_97 R_bl
Rbb_86_96 bitb_86_96 bitb_86_97 R_bl
Cb_86_96 bit_86_96 gnd C_bl
Cbb_86_96 bitb_86_96 gnd C_bl
Rb_86_97 bit_86_97 bit_86_98 R_bl
Rbb_86_97 bitb_86_97 bitb_86_98 R_bl
Cb_86_97 bit_86_97 gnd C_bl
Cbb_86_97 bitb_86_97 gnd C_bl
Rb_86_98 bit_86_98 bit_86_99 R_bl
Rbb_86_98 bitb_86_98 bitb_86_99 R_bl
Cb_86_98 bit_86_98 gnd C_bl
Cbb_86_98 bitb_86_98 gnd C_bl
Rb_86_99 bit_86_99 bit_86_100 R_bl
Rbb_86_99 bitb_86_99 bitb_86_100 R_bl
Cb_86_99 bit_86_99 gnd C_bl
Cbb_86_99 bitb_86_99 gnd C_bl
Rb_87_0 bit_87_0 bit_87_1 R_bl
Rbb_87_0 bitb_87_0 bitb_87_1 R_bl
Cb_87_0 bit_87_0 gnd C_bl
Cbb_87_0 bitb_87_0 gnd C_bl
Rb_87_1 bit_87_1 bit_87_2 R_bl
Rbb_87_1 bitb_87_1 bitb_87_2 R_bl
Cb_87_1 bit_87_1 gnd C_bl
Cbb_87_1 bitb_87_1 gnd C_bl
Rb_87_2 bit_87_2 bit_87_3 R_bl
Rbb_87_2 bitb_87_2 bitb_87_3 R_bl
Cb_87_2 bit_87_2 gnd C_bl
Cbb_87_2 bitb_87_2 gnd C_bl
Rb_87_3 bit_87_3 bit_87_4 R_bl
Rbb_87_3 bitb_87_3 bitb_87_4 R_bl
Cb_87_3 bit_87_3 gnd C_bl
Cbb_87_3 bitb_87_3 gnd C_bl
Rb_87_4 bit_87_4 bit_87_5 R_bl
Rbb_87_4 bitb_87_4 bitb_87_5 R_bl
Cb_87_4 bit_87_4 gnd C_bl
Cbb_87_4 bitb_87_4 gnd C_bl
Rb_87_5 bit_87_5 bit_87_6 R_bl
Rbb_87_5 bitb_87_5 bitb_87_6 R_bl
Cb_87_5 bit_87_5 gnd C_bl
Cbb_87_5 bitb_87_5 gnd C_bl
Rb_87_6 bit_87_6 bit_87_7 R_bl
Rbb_87_6 bitb_87_6 bitb_87_7 R_bl
Cb_87_6 bit_87_6 gnd C_bl
Cbb_87_6 bitb_87_6 gnd C_bl
Rb_87_7 bit_87_7 bit_87_8 R_bl
Rbb_87_7 bitb_87_7 bitb_87_8 R_bl
Cb_87_7 bit_87_7 gnd C_bl
Cbb_87_7 bitb_87_7 gnd C_bl
Rb_87_8 bit_87_8 bit_87_9 R_bl
Rbb_87_8 bitb_87_8 bitb_87_9 R_bl
Cb_87_8 bit_87_8 gnd C_bl
Cbb_87_8 bitb_87_8 gnd C_bl
Rb_87_9 bit_87_9 bit_87_10 R_bl
Rbb_87_9 bitb_87_9 bitb_87_10 R_bl
Cb_87_9 bit_87_9 gnd C_bl
Cbb_87_9 bitb_87_9 gnd C_bl
Rb_87_10 bit_87_10 bit_87_11 R_bl
Rbb_87_10 bitb_87_10 bitb_87_11 R_bl
Cb_87_10 bit_87_10 gnd C_bl
Cbb_87_10 bitb_87_10 gnd C_bl
Rb_87_11 bit_87_11 bit_87_12 R_bl
Rbb_87_11 bitb_87_11 bitb_87_12 R_bl
Cb_87_11 bit_87_11 gnd C_bl
Cbb_87_11 bitb_87_11 gnd C_bl
Rb_87_12 bit_87_12 bit_87_13 R_bl
Rbb_87_12 bitb_87_12 bitb_87_13 R_bl
Cb_87_12 bit_87_12 gnd C_bl
Cbb_87_12 bitb_87_12 gnd C_bl
Rb_87_13 bit_87_13 bit_87_14 R_bl
Rbb_87_13 bitb_87_13 bitb_87_14 R_bl
Cb_87_13 bit_87_13 gnd C_bl
Cbb_87_13 bitb_87_13 gnd C_bl
Rb_87_14 bit_87_14 bit_87_15 R_bl
Rbb_87_14 bitb_87_14 bitb_87_15 R_bl
Cb_87_14 bit_87_14 gnd C_bl
Cbb_87_14 bitb_87_14 gnd C_bl
Rb_87_15 bit_87_15 bit_87_16 R_bl
Rbb_87_15 bitb_87_15 bitb_87_16 R_bl
Cb_87_15 bit_87_15 gnd C_bl
Cbb_87_15 bitb_87_15 gnd C_bl
Rb_87_16 bit_87_16 bit_87_17 R_bl
Rbb_87_16 bitb_87_16 bitb_87_17 R_bl
Cb_87_16 bit_87_16 gnd C_bl
Cbb_87_16 bitb_87_16 gnd C_bl
Rb_87_17 bit_87_17 bit_87_18 R_bl
Rbb_87_17 bitb_87_17 bitb_87_18 R_bl
Cb_87_17 bit_87_17 gnd C_bl
Cbb_87_17 bitb_87_17 gnd C_bl
Rb_87_18 bit_87_18 bit_87_19 R_bl
Rbb_87_18 bitb_87_18 bitb_87_19 R_bl
Cb_87_18 bit_87_18 gnd C_bl
Cbb_87_18 bitb_87_18 gnd C_bl
Rb_87_19 bit_87_19 bit_87_20 R_bl
Rbb_87_19 bitb_87_19 bitb_87_20 R_bl
Cb_87_19 bit_87_19 gnd C_bl
Cbb_87_19 bitb_87_19 gnd C_bl
Rb_87_20 bit_87_20 bit_87_21 R_bl
Rbb_87_20 bitb_87_20 bitb_87_21 R_bl
Cb_87_20 bit_87_20 gnd C_bl
Cbb_87_20 bitb_87_20 gnd C_bl
Rb_87_21 bit_87_21 bit_87_22 R_bl
Rbb_87_21 bitb_87_21 bitb_87_22 R_bl
Cb_87_21 bit_87_21 gnd C_bl
Cbb_87_21 bitb_87_21 gnd C_bl
Rb_87_22 bit_87_22 bit_87_23 R_bl
Rbb_87_22 bitb_87_22 bitb_87_23 R_bl
Cb_87_22 bit_87_22 gnd C_bl
Cbb_87_22 bitb_87_22 gnd C_bl
Rb_87_23 bit_87_23 bit_87_24 R_bl
Rbb_87_23 bitb_87_23 bitb_87_24 R_bl
Cb_87_23 bit_87_23 gnd C_bl
Cbb_87_23 bitb_87_23 gnd C_bl
Rb_87_24 bit_87_24 bit_87_25 R_bl
Rbb_87_24 bitb_87_24 bitb_87_25 R_bl
Cb_87_24 bit_87_24 gnd C_bl
Cbb_87_24 bitb_87_24 gnd C_bl
Rb_87_25 bit_87_25 bit_87_26 R_bl
Rbb_87_25 bitb_87_25 bitb_87_26 R_bl
Cb_87_25 bit_87_25 gnd C_bl
Cbb_87_25 bitb_87_25 gnd C_bl
Rb_87_26 bit_87_26 bit_87_27 R_bl
Rbb_87_26 bitb_87_26 bitb_87_27 R_bl
Cb_87_26 bit_87_26 gnd C_bl
Cbb_87_26 bitb_87_26 gnd C_bl
Rb_87_27 bit_87_27 bit_87_28 R_bl
Rbb_87_27 bitb_87_27 bitb_87_28 R_bl
Cb_87_27 bit_87_27 gnd C_bl
Cbb_87_27 bitb_87_27 gnd C_bl
Rb_87_28 bit_87_28 bit_87_29 R_bl
Rbb_87_28 bitb_87_28 bitb_87_29 R_bl
Cb_87_28 bit_87_28 gnd C_bl
Cbb_87_28 bitb_87_28 gnd C_bl
Rb_87_29 bit_87_29 bit_87_30 R_bl
Rbb_87_29 bitb_87_29 bitb_87_30 R_bl
Cb_87_29 bit_87_29 gnd C_bl
Cbb_87_29 bitb_87_29 gnd C_bl
Rb_87_30 bit_87_30 bit_87_31 R_bl
Rbb_87_30 bitb_87_30 bitb_87_31 R_bl
Cb_87_30 bit_87_30 gnd C_bl
Cbb_87_30 bitb_87_30 gnd C_bl
Rb_87_31 bit_87_31 bit_87_32 R_bl
Rbb_87_31 bitb_87_31 bitb_87_32 R_bl
Cb_87_31 bit_87_31 gnd C_bl
Cbb_87_31 bitb_87_31 gnd C_bl
Rb_87_32 bit_87_32 bit_87_33 R_bl
Rbb_87_32 bitb_87_32 bitb_87_33 R_bl
Cb_87_32 bit_87_32 gnd C_bl
Cbb_87_32 bitb_87_32 gnd C_bl
Rb_87_33 bit_87_33 bit_87_34 R_bl
Rbb_87_33 bitb_87_33 bitb_87_34 R_bl
Cb_87_33 bit_87_33 gnd C_bl
Cbb_87_33 bitb_87_33 gnd C_bl
Rb_87_34 bit_87_34 bit_87_35 R_bl
Rbb_87_34 bitb_87_34 bitb_87_35 R_bl
Cb_87_34 bit_87_34 gnd C_bl
Cbb_87_34 bitb_87_34 gnd C_bl
Rb_87_35 bit_87_35 bit_87_36 R_bl
Rbb_87_35 bitb_87_35 bitb_87_36 R_bl
Cb_87_35 bit_87_35 gnd C_bl
Cbb_87_35 bitb_87_35 gnd C_bl
Rb_87_36 bit_87_36 bit_87_37 R_bl
Rbb_87_36 bitb_87_36 bitb_87_37 R_bl
Cb_87_36 bit_87_36 gnd C_bl
Cbb_87_36 bitb_87_36 gnd C_bl
Rb_87_37 bit_87_37 bit_87_38 R_bl
Rbb_87_37 bitb_87_37 bitb_87_38 R_bl
Cb_87_37 bit_87_37 gnd C_bl
Cbb_87_37 bitb_87_37 gnd C_bl
Rb_87_38 bit_87_38 bit_87_39 R_bl
Rbb_87_38 bitb_87_38 bitb_87_39 R_bl
Cb_87_38 bit_87_38 gnd C_bl
Cbb_87_38 bitb_87_38 gnd C_bl
Rb_87_39 bit_87_39 bit_87_40 R_bl
Rbb_87_39 bitb_87_39 bitb_87_40 R_bl
Cb_87_39 bit_87_39 gnd C_bl
Cbb_87_39 bitb_87_39 gnd C_bl
Rb_87_40 bit_87_40 bit_87_41 R_bl
Rbb_87_40 bitb_87_40 bitb_87_41 R_bl
Cb_87_40 bit_87_40 gnd C_bl
Cbb_87_40 bitb_87_40 gnd C_bl
Rb_87_41 bit_87_41 bit_87_42 R_bl
Rbb_87_41 bitb_87_41 bitb_87_42 R_bl
Cb_87_41 bit_87_41 gnd C_bl
Cbb_87_41 bitb_87_41 gnd C_bl
Rb_87_42 bit_87_42 bit_87_43 R_bl
Rbb_87_42 bitb_87_42 bitb_87_43 R_bl
Cb_87_42 bit_87_42 gnd C_bl
Cbb_87_42 bitb_87_42 gnd C_bl
Rb_87_43 bit_87_43 bit_87_44 R_bl
Rbb_87_43 bitb_87_43 bitb_87_44 R_bl
Cb_87_43 bit_87_43 gnd C_bl
Cbb_87_43 bitb_87_43 gnd C_bl
Rb_87_44 bit_87_44 bit_87_45 R_bl
Rbb_87_44 bitb_87_44 bitb_87_45 R_bl
Cb_87_44 bit_87_44 gnd C_bl
Cbb_87_44 bitb_87_44 gnd C_bl
Rb_87_45 bit_87_45 bit_87_46 R_bl
Rbb_87_45 bitb_87_45 bitb_87_46 R_bl
Cb_87_45 bit_87_45 gnd C_bl
Cbb_87_45 bitb_87_45 gnd C_bl
Rb_87_46 bit_87_46 bit_87_47 R_bl
Rbb_87_46 bitb_87_46 bitb_87_47 R_bl
Cb_87_46 bit_87_46 gnd C_bl
Cbb_87_46 bitb_87_46 gnd C_bl
Rb_87_47 bit_87_47 bit_87_48 R_bl
Rbb_87_47 bitb_87_47 bitb_87_48 R_bl
Cb_87_47 bit_87_47 gnd C_bl
Cbb_87_47 bitb_87_47 gnd C_bl
Rb_87_48 bit_87_48 bit_87_49 R_bl
Rbb_87_48 bitb_87_48 bitb_87_49 R_bl
Cb_87_48 bit_87_48 gnd C_bl
Cbb_87_48 bitb_87_48 gnd C_bl
Rb_87_49 bit_87_49 bit_87_50 R_bl
Rbb_87_49 bitb_87_49 bitb_87_50 R_bl
Cb_87_49 bit_87_49 gnd C_bl
Cbb_87_49 bitb_87_49 gnd C_bl
Rb_87_50 bit_87_50 bit_87_51 R_bl
Rbb_87_50 bitb_87_50 bitb_87_51 R_bl
Cb_87_50 bit_87_50 gnd C_bl
Cbb_87_50 bitb_87_50 gnd C_bl
Rb_87_51 bit_87_51 bit_87_52 R_bl
Rbb_87_51 bitb_87_51 bitb_87_52 R_bl
Cb_87_51 bit_87_51 gnd C_bl
Cbb_87_51 bitb_87_51 gnd C_bl
Rb_87_52 bit_87_52 bit_87_53 R_bl
Rbb_87_52 bitb_87_52 bitb_87_53 R_bl
Cb_87_52 bit_87_52 gnd C_bl
Cbb_87_52 bitb_87_52 gnd C_bl
Rb_87_53 bit_87_53 bit_87_54 R_bl
Rbb_87_53 bitb_87_53 bitb_87_54 R_bl
Cb_87_53 bit_87_53 gnd C_bl
Cbb_87_53 bitb_87_53 gnd C_bl
Rb_87_54 bit_87_54 bit_87_55 R_bl
Rbb_87_54 bitb_87_54 bitb_87_55 R_bl
Cb_87_54 bit_87_54 gnd C_bl
Cbb_87_54 bitb_87_54 gnd C_bl
Rb_87_55 bit_87_55 bit_87_56 R_bl
Rbb_87_55 bitb_87_55 bitb_87_56 R_bl
Cb_87_55 bit_87_55 gnd C_bl
Cbb_87_55 bitb_87_55 gnd C_bl
Rb_87_56 bit_87_56 bit_87_57 R_bl
Rbb_87_56 bitb_87_56 bitb_87_57 R_bl
Cb_87_56 bit_87_56 gnd C_bl
Cbb_87_56 bitb_87_56 gnd C_bl
Rb_87_57 bit_87_57 bit_87_58 R_bl
Rbb_87_57 bitb_87_57 bitb_87_58 R_bl
Cb_87_57 bit_87_57 gnd C_bl
Cbb_87_57 bitb_87_57 gnd C_bl
Rb_87_58 bit_87_58 bit_87_59 R_bl
Rbb_87_58 bitb_87_58 bitb_87_59 R_bl
Cb_87_58 bit_87_58 gnd C_bl
Cbb_87_58 bitb_87_58 gnd C_bl
Rb_87_59 bit_87_59 bit_87_60 R_bl
Rbb_87_59 bitb_87_59 bitb_87_60 R_bl
Cb_87_59 bit_87_59 gnd C_bl
Cbb_87_59 bitb_87_59 gnd C_bl
Rb_87_60 bit_87_60 bit_87_61 R_bl
Rbb_87_60 bitb_87_60 bitb_87_61 R_bl
Cb_87_60 bit_87_60 gnd C_bl
Cbb_87_60 bitb_87_60 gnd C_bl
Rb_87_61 bit_87_61 bit_87_62 R_bl
Rbb_87_61 bitb_87_61 bitb_87_62 R_bl
Cb_87_61 bit_87_61 gnd C_bl
Cbb_87_61 bitb_87_61 gnd C_bl
Rb_87_62 bit_87_62 bit_87_63 R_bl
Rbb_87_62 bitb_87_62 bitb_87_63 R_bl
Cb_87_62 bit_87_62 gnd C_bl
Cbb_87_62 bitb_87_62 gnd C_bl
Rb_87_63 bit_87_63 bit_87_64 R_bl
Rbb_87_63 bitb_87_63 bitb_87_64 R_bl
Cb_87_63 bit_87_63 gnd C_bl
Cbb_87_63 bitb_87_63 gnd C_bl
Rb_87_64 bit_87_64 bit_87_65 R_bl
Rbb_87_64 bitb_87_64 bitb_87_65 R_bl
Cb_87_64 bit_87_64 gnd C_bl
Cbb_87_64 bitb_87_64 gnd C_bl
Rb_87_65 bit_87_65 bit_87_66 R_bl
Rbb_87_65 bitb_87_65 bitb_87_66 R_bl
Cb_87_65 bit_87_65 gnd C_bl
Cbb_87_65 bitb_87_65 gnd C_bl
Rb_87_66 bit_87_66 bit_87_67 R_bl
Rbb_87_66 bitb_87_66 bitb_87_67 R_bl
Cb_87_66 bit_87_66 gnd C_bl
Cbb_87_66 bitb_87_66 gnd C_bl
Rb_87_67 bit_87_67 bit_87_68 R_bl
Rbb_87_67 bitb_87_67 bitb_87_68 R_bl
Cb_87_67 bit_87_67 gnd C_bl
Cbb_87_67 bitb_87_67 gnd C_bl
Rb_87_68 bit_87_68 bit_87_69 R_bl
Rbb_87_68 bitb_87_68 bitb_87_69 R_bl
Cb_87_68 bit_87_68 gnd C_bl
Cbb_87_68 bitb_87_68 gnd C_bl
Rb_87_69 bit_87_69 bit_87_70 R_bl
Rbb_87_69 bitb_87_69 bitb_87_70 R_bl
Cb_87_69 bit_87_69 gnd C_bl
Cbb_87_69 bitb_87_69 gnd C_bl
Rb_87_70 bit_87_70 bit_87_71 R_bl
Rbb_87_70 bitb_87_70 bitb_87_71 R_bl
Cb_87_70 bit_87_70 gnd C_bl
Cbb_87_70 bitb_87_70 gnd C_bl
Rb_87_71 bit_87_71 bit_87_72 R_bl
Rbb_87_71 bitb_87_71 bitb_87_72 R_bl
Cb_87_71 bit_87_71 gnd C_bl
Cbb_87_71 bitb_87_71 gnd C_bl
Rb_87_72 bit_87_72 bit_87_73 R_bl
Rbb_87_72 bitb_87_72 bitb_87_73 R_bl
Cb_87_72 bit_87_72 gnd C_bl
Cbb_87_72 bitb_87_72 gnd C_bl
Rb_87_73 bit_87_73 bit_87_74 R_bl
Rbb_87_73 bitb_87_73 bitb_87_74 R_bl
Cb_87_73 bit_87_73 gnd C_bl
Cbb_87_73 bitb_87_73 gnd C_bl
Rb_87_74 bit_87_74 bit_87_75 R_bl
Rbb_87_74 bitb_87_74 bitb_87_75 R_bl
Cb_87_74 bit_87_74 gnd C_bl
Cbb_87_74 bitb_87_74 gnd C_bl
Rb_87_75 bit_87_75 bit_87_76 R_bl
Rbb_87_75 bitb_87_75 bitb_87_76 R_bl
Cb_87_75 bit_87_75 gnd C_bl
Cbb_87_75 bitb_87_75 gnd C_bl
Rb_87_76 bit_87_76 bit_87_77 R_bl
Rbb_87_76 bitb_87_76 bitb_87_77 R_bl
Cb_87_76 bit_87_76 gnd C_bl
Cbb_87_76 bitb_87_76 gnd C_bl
Rb_87_77 bit_87_77 bit_87_78 R_bl
Rbb_87_77 bitb_87_77 bitb_87_78 R_bl
Cb_87_77 bit_87_77 gnd C_bl
Cbb_87_77 bitb_87_77 gnd C_bl
Rb_87_78 bit_87_78 bit_87_79 R_bl
Rbb_87_78 bitb_87_78 bitb_87_79 R_bl
Cb_87_78 bit_87_78 gnd C_bl
Cbb_87_78 bitb_87_78 gnd C_bl
Rb_87_79 bit_87_79 bit_87_80 R_bl
Rbb_87_79 bitb_87_79 bitb_87_80 R_bl
Cb_87_79 bit_87_79 gnd C_bl
Cbb_87_79 bitb_87_79 gnd C_bl
Rb_87_80 bit_87_80 bit_87_81 R_bl
Rbb_87_80 bitb_87_80 bitb_87_81 R_bl
Cb_87_80 bit_87_80 gnd C_bl
Cbb_87_80 bitb_87_80 gnd C_bl
Rb_87_81 bit_87_81 bit_87_82 R_bl
Rbb_87_81 bitb_87_81 bitb_87_82 R_bl
Cb_87_81 bit_87_81 gnd C_bl
Cbb_87_81 bitb_87_81 gnd C_bl
Rb_87_82 bit_87_82 bit_87_83 R_bl
Rbb_87_82 bitb_87_82 bitb_87_83 R_bl
Cb_87_82 bit_87_82 gnd C_bl
Cbb_87_82 bitb_87_82 gnd C_bl
Rb_87_83 bit_87_83 bit_87_84 R_bl
Rbb_87_83 bitb_87_83 bitb_87_84 R_bl
Cb_87_83 bit_87_83 gnd C_bl
Cbb_87_83 bitb_87_83 gnd C_bl
Rb_87_84 bit_87_84 bit_87_85 R_bl
Rbb_87_84 bitb_87_84 bitb_87_85 R_bl
Cb_87_84 bit_87_84 gnd C_bl
Cbb_87_84 bitb_87_84 gnd C_bl
Rb_87_85 bit_87_85 bit_87_86 R_bl
Rbb_87_85 bitb_87_85 bitb_87_86 R_bl
Cb_87_85 bit_87_85 gnd C_bl
Cbb_87_85 bitb_87_85 gnd C_bl
Rb_87_86 bit_87_86 bit_87_87 R_bl
Rbb_87_86 bitb_87_86 bitb_87_87 R_bl
Cb_87_86 bit_87_86 gnd C_bl
Cbb_87_86 bitb_87_86 gnd C_bl
Rb_87_87 bit_87_87 bit_87_88 R_bl
Rbb_87_87 bitb_87_87 bitb_87_88 R_bl
Cb_87_87 bit_87_87 gnd C_bl
Cbb_87_87 bitb_87_87 gnd C_bl
Rb_87_88 bit_87_88 bit_87_89 R_bl
Rbb_87_88 bitb_87_88 bitb_87_89 R_bl
Cb_87_88 bit_87_88 gnd C_bl
Cbb_87_88 bitb_87_88 gnd C_bl
Rb_87_89 bit_87_89 bit_87_90 R_bl
Rbb_87_89 bitb_87_89 bitb_87_90 R_bl
Cb_87_89 bit_87_89 gnd C_bl
Cbb_87_89 bitb_87_89 gnd C_bl
Rb_87_90 bit_87_90 bit_87_91 R_bl
Rbb_87_90 bitb_87_90 bitb_87_91 R_bl
Cb_87_90 bit_87_90 gnd C_bl
Cbb_87_90 bitb_87_90 gnd C_bl
Rb_87_91 bit_87_91 bit_87_92 R_bl
Rbb_87_91 bitb_87_91 bitb_87_92 R_bl
Cb_87_91 bit_87_91 gnd C_bl
Cbb_87_91 bitb_87_91 gnd C_bl
Rb_87_92 bit_87_92 bit_87_93 R_bl
Rbb_87_92 bitb_87_92 bitb_87_93 R_bl
Cb_87_92 bit_87_92 gnd C_bl
Cbb_87_92 bitb_87_92 gnd C_bl
Rb_87_93 bit_87_93 bit_87_94 R_bl
Rbb_87_93 bitb_87_93 bitb_87_94 R_bl
Cb_87_93 bit_87_93 gnd C_bl
Cbb_87_93 bitb_87_93 gnd C_bl
Rb_87_94 bit_87_94 bit_87_95 R_bl
Rbb_87_94 bitb_87_94 bitb_87_95 R_bl
Cb_87_94 bit_87_94 gnd C_bl
Cbb_87_94 bitb_87_94 gnd C_bl
Rb_87_95 bit_87_95 bit_87_96 R_bl
Rbb_87_95 bitb_87_95 bitb_87_96 R_bl
Cb_87_95 bit_87_95 gnd C_bl
Cbb_87_95 bitb_87_95 gnd C_bl
Rb_87_96 bit_87_96 bit_87_97 R_bl
Rbb_87_96 bitb_87_96 bitb_87_97 R_bl
Cb_87_96 bit_87_96 gnd C_bl
Cbb_87_96 bitb_87_96 gnd C_bl
Rb_87_97 bit_87_97 bit_87_98 R_bl
Rbb_87_97 bitb_87_97 bitb_87_98 R_bl
Cb_87_97 bit_87_97 gnd C_bl
Cbb_87_97 bitb_87_97 gnd C_bl
Rb_87_98 bit_87_98 bit_87_99 R_bl
Rbb_87_98 bitb_87_98 bitb_87_99 R_bl
Cb_87_98 bit_87_98 gnd C_bl
Cbb_87_98 bitb_87_98 gnd C_bl
Rb_87_99 bit_87_99 bit_87_100 R_bl
Rbb_87_99 bitb_87_99 bitb_87_100 R_bl
Cb_87_99 bit_87_99 gnd C_bl
Cbb_87_99 bitb_87_99 gnd C_bl
Rb_88_0 bit_88_0 bit_88_1 R_bl
Rbb_88_0 bitb_88_0 bitb_88_1 R_bl
Cb_88_0 bit_88_0 gnd C_bl
Cbb_88_0 bitb_88_0 gnd C_bl
Rb_88_1 bit_88_1 bit_88_2 R_bl
Rbb_88_1 bitb_88_1 bitb_88_2 R_bl
Cb_88_1 bit_88_1 gnd C_bl
Cbb_88_1 bitb_88_1 gnd C_bl
Rb_88_2 bit_88_2 bit_88_3 R_bl
Rbb_88_2 bitb_88_2 bitb_88_3 R_bl
Cb_88_2 bit_88_2 gnd C_bl
Cbb_88_2 bitb_88_2 gnd C_bl
Rb_88_3 bit_88_3 bit_88_4 R_bl
Rbb_88_3 bitb_88_3 bitb_88_4 R_bl
Cb_88_3 bit_88_3 gnd C_bl
Cbb_88_3 bitb_88_3 gnd C_bl
Rb_88_4 bit_88_4 bit_88_5 R_bl
Rbb_88_4 bitb_88_4 bitb_88_5 R_bl
Cb_88_4 bit_88_4 gnd C_bl
Cbb_88_4 bitb_88_4 gnd C_bl
Rb_88_5 bit_88_5 bit_88_6 R_bl
Rbb_88_5 bitb_88_5 bitb_88_6 R_bl
Cb_88_5 bit_88_5 gnd C_bl
Cbb_88_5 bitb_88_5 gnd C_bl
Rb_88_6 bit_88_6 bit_88_7 R_bl
Rbb_88_6 bitb_88_6 bitb_88_7 R_bl
Cb_88_6 bit_88_6 gnd C_bl
Cbb_88_6 bitb_88_6 gnd C_bl
Rb_88_7 bit_88_7 bit_88_8 R_bl
Rbb_88_7 bitb_88_7 bitb_88_8 R_bl
Cb_88_7 bit_88_7 gnd C_bl
Cbb_88_7 bitb_88_7 gnd C_bl
Rb_88_8 bit_88_8 bit_88_9 R_bl
Rbb_88_8 bitb_88_8 bitb_88_9 R_bl
Cb_88_8 bit_88_8 gnd C_bl
Cbb_88_8 bitb_88_8 gnd C_bl
Rb_88_9 bit_88_9 bit_88_10 R_bl
Rbb_88_9 bitb_88_9 bitb_88_10 R_bl
Cb_88_9 bit_88_9 gnd C_bl
Cbb_88_9 bitb_88_9 gnd C_bl
Rb_88_10 bit_88_10 bit_88_11 R_bl
Rbb_88_10 bitb_88_10 bitb_88_11 R_bl
Cb_88_10 bit_88_10 gnd C_bl
Cbb_88_10 bitb_88_10 gnd C_bl
Rb_88_11 bit_88_11 bit_88_12 R_bl
Rbb_88_11 bitb_88_11 bitb_88_12 R_bl
Cb_88_11 bit_88_11 gnd C_bl
Cbb_88_11 bitb_88_11 gnd C_bl
Rb_88_12 bit_88_12 bit_88_13 R_bl
Rbb_88_12 bitb_88_12 bitb_88_13 R_bl
Cb_88_12 bit_88_12 gnd C_bl
Cbb_88_12 bitb_88_12 gnd C_bl
Rb_88_13 bit_88_13 bit_88_14 R_bl
Rbb_88_13 bitb_88_13 bitb_88_14 R_bl
Cb_88_13 bit_88_13 gnd C_bl
Cbb_88_13 bitb_88_13 gnd C_bl
Rb_88_14 bit_88_14 bit_88_15 R_bl
Rbb_88_14 bitb_88_14 bitb_88_15 R_bl
Cb_88_14 bit_88_14 gnd C_bl
Cbb_88_14 bitb_88_14 gnd C_bl
Rb_88_15 bit_88_15 bit_88_16 R_bl
Rbb_88_15 bitb_88_15 bitb_88_16 R_bl
Cb_88_15 bit_88_15 gnd C_bl
Cbb_88_15 bitb_88_15 gnd C_bl
Rb_88_16 bit_88_16 bit_88_17 R_bl
Rbb_88_16 bitb_88_16 bitb_88_17 R_bl
Cb_88_16 bit_88_16 gnd C_bl
Cbb_88_16 bitb_88_16 gnd C_bl
Rb_88_17 bit_88_17 bit_88_18 R_bl
Rbb_88_17 bitb_88_17 bitb_88_18 R_bl
Cb_88_17 bit_88_17 gnd C_bl
Cbb_88_17 bitb_88_17 gnd C_bl
Rb_88_18 bit_88_18 bit_88_19 R_bl
Rbb_88_18 bitb_88_18 bitb_88_19 R_bl
Cb_88_18 bit_88_18 gnd C_bl
Cbb_88_18 bitb_88_18 gnd C_bl
Rb_88_19 bit_88_19 bit_88_20 R_bl
Rbb_88_19 bitb_88_19 bitb_88_20 R_bl
Cb_88_19 bit_88_19 gnd C_bl
Cbb_88_19 bitb_88_19 gnd C_bl
Rb_88_20 bit_88_20 bit_88_21 R_bl
Rbb_88_20 bitb_88_20 bitb_88_21 R_bl
Cb_88_20 bit_88_20 gnd C_bl
Cbb_88_20 bitb_88_20 gnd C_bl
Rb_88_21 bit_88_21 bit_88_22 R_bl
Rbb_88_21 bitb_88_21 bitb_88_22 R_bl
Cb_88_21 bit_88_21 gnd C_bl
Cbb_88_21 bitb_88_21 gnd C_bl
Rb_88_22 bit_88_22 bit_88_23 R_bl
Rbb_88_22 bitb_88_22 bitb_88_23 R_bl
Cb_88_22 bit_88_22 gnd C_bl
Cbb_88_22 bitb_88_22 gnd C_bl
Rb_88_23 bit_88_23 bit_88_24 R_bl
Rbb_88_23 bitb_88_23 bitb_88_24 R_bl
Cb_88_23 bit_88_23 gnd C_bl
Cbb_88_23 bitb_88_23 gnd C_bl
Rb_88_24 bit_88_24 bit_88_25 R_bl
Rbb_88_24 bitb_88_24 bitb_88_25 R_bl
Cb_88_24 bit_88_24 gnd C_bl
Cbb_88_24 bitb_88_24 gnd C_bl
Rb_88_25 bit_88_25 bit_88_26 R_bl
Rbb_88_25 bitb_88_25 bitb_88_26 R_bl
Cb_88_25 bit_88_25 gnd C_bl
Cbb_88_25 bitb_88_25 gnd C_bl
Rb_88_26 bit_88_26 bit_88_27 R_bl
Rbb_88_26 bitb_88_26 bitb_88_27 R_bl
Cb_88_26 bit_88_26 gnd C_bl
Cbb_88_26 bitb_88_26 gnd C_bl
Rb_88_27 bit_88_27 bit_88_28 R_bl
Rbb_88_27 bitb_88_27 bitb_88_28 R_bl
Cb_88_27 bit_88_27 gnd C_bl
Cbb_88_27 bitb_88_27 gnd C_bl
Rb_88_28 bit_88_28 bit_88_29 R_bl
Rbb_88_28 bitb_88_28 bitb_88_29 R_bl
Cb_88_28 bit_88_28 gnd C_bl
Cbb_88_28 bitb_88_28 gnd C_bl
Rb_88_29 bit_88_29 bit_88_30 R_bl
Rbb_88_29 bitb_88_29 bitb_88_30 R_bl
Cb_88_29 bit_88_29 gnd C_bl
Cbb_88_29 bitb_88_29 gnd C_bl
Rb_88_30 bit_88_30 bit_88_31 R_bl
Rbb_88_30 bitb_88_30 bitb_88_31 R_bl
Cb_88_30 bit_88_30 gnd C_bl
Cbb_88_30 bitb_88_30 gnd C_bl
Rb_88_31 bit_88_31 bit_88_32 R_bl
Rbb_88_31 bitb_88_31 bitb_88_32 R_bl
Cb_88_31 bit_88_31 gnd C_bl
Cbb_88_31 bitb_88_31 gnd C_bl
Rb_88_32 bit_88_32 bit_88_33 R_bl
Rbb_88_32 bitb_88_32 bitb_88_33 R_bl
Cb_88_32 bit_88_32 gnd C_bl
Cbb_88_32 bitb_88_32 gnd C_bl
Rb_88_33 bit_88_33 bit_88_34 R_bl
Rbb_88_33 bitb_88_33 bitb_88_34 R_bl
Cb_88_33 bit_88_33 gnd C_bl
Cbb_88_33 bitb_88_33 gnd C_bl
Rb_88_34 bit_88_34 bit_88_35 R_bl
Rbb_88_34 bitb_88_34 bitb_88_35 R_bl
Cb_88_34 bit_88_34 gnd C_bl
Cbb_88_34 bitb_88_34 gnd C_bl
Rb_88_35 bit_88_35 bit_88_36 R_bl
Rbb_88_35 bitb_88_35 bitb_88_36 R_bl
Cb_88_35 bit_88_35 gnd C_bl
Cbb_88_35 bitb_88_35 gnd C_bl
Rb_88_36 bit_88_36 bit_88_37 R_bl
Rbb_88_36 bitb_88_36 bitb_88_37 R_bl
Cb_88_36 bit_88_36 gnd C_bl
Cbb_88_36 bitb_88_36 gnd C_bl
Rb_88_37 bit_88_37 bit_88_38 R_bl
Rbb_88_37 bitb_88_37 bitb_88_38 R_bl
Cb_88_37 bit_88_37 gnd C_bl
Cbb_88_37 bitb_88_37 gnd C_bl
Rb_88_38 bit_88_38 bit_88_39 R_bl
Rbb_88_38 bitb_88_38 bitb_88_39 R_bl
Cb_88_38 bit_88_38 gnd C_bl
Cbb_88_38 bitb_88_38 gnd C_bl
Rb_88_39 bit_88_39 bit_88_40 R_bl
Rbb_88_39 bitb_88_39 bitb_88_40 R_bl
Cb_88_39 bit_88_39 gnd C_bl
Cbb_88_39 bitb_88_39 gnd C_bl
Rb_88_40 bit_88_40 bit_88_41 R_bl
Rbb_88_40 bitb_88_40 bitb_88_41 R_bl
Cb_88_40 bit_88_40 gnd C_bl
Cbb_88_40 bitb_88_40 gnd C_bl
Rb_88_41 bit_88_41 bit_88_42 R_bl
Rbb_88_41 bitb_88_41 bitb_88_42 R_bl
Cb_88_41 bit_88_41 gnd C_bl
Cbb_88_41 bitb_88_41 gnd C_bl
Rb_88_42 bit_88_42 bit_88_43 R_bl
Rbb_88_42 bitb_88_42 bitb_88_43 R_bl
Cb_88_42 bit_88_42 gnd C_bl
Cbb_88_42 bitb_88_42 gnd C_bl
Rb_88_43 bit_88_43 bit_88_44 R_bl
Rbb_88_43 bitb_88_43 bitb_88_44 R_bl
Cb_88_43 bit_88_43 gnd C_bl
Cbb_88_43 bitb_88_43 gnd C_bl
Rb_88_44 bit_88_44 bit_88_45 R_bl
Rbb_88_44 bitb_88_44 bitb_88_45 R_bl
Cb_88_44 bit_88_44 gnd C_bl
Cbb_88_44 bitb_88_44 gnd C_bl
Rb_88_45 bit_88_45 bit_88_46 R_bl
Rbb_88_45 bitb_88_45 bitb_88_46 R_bl
Cb_88_45 bit_88_45 gnd C_bl
Cbb_88_45 bitb_88_45 gnd C_bl
Rb_88_46 bit_88_46 bit_88_47 R_bl
Rbb_88_46 bitb_88_46 bitb_88_47 R_bl
Cb_88_46 bit_88_46 gnd C_bl
Cbb_88_46 bitb_88_46 gnd C_bl
Rb_88_47 bit_88_47 bit_88_48 R_bl
Rbb_88_47 bitb_88_47 bitb_88_48 R_bl
Cb_88_47 bit_88_47 gnd C_bl
Cbb_88_47 bitb_88_47 gnd C_bl
Rb_88_48 bit_88_48 bit_88_49 R_bl
Rbb_88_48 bitb_88_48 bitb_88_49 R_bl
Cb_88_48 bit_88_48 gnd C_bl
Cbb_88_48 bitb_88_48 gnd C_bl
Rb_88_49 bit_88_49 bit_88_50 R_bl
Rbb_88_49 bitb_88_49 bitb_88_50 R_bl
Cb_88_49 bit_88_49 gnd C_bl
Cbb_88_49 bitb_88_49 gnd C_bl
Rb_88_50 bit_88_50 bit_88_51 R_bl
Rbb_88_50 bitb_88_50 bitb_88_51 R_bl
Cb_88_50 bit_88_50 gnd C_bl
Cbb_88_50 bitb_88_50 gnd C_bl
Rb_88_51 bit_88_51 bit_88_52 R_bl
Rbb_88_51 bitb_88_51 bitb_88_52 R_bl
Cb_88_51 bit_88_51 gnd C_bl
Cbb_88_51 bitb_88_51 gnd C_bl
Rb_88_52 bit_88_52 bit_88_53 R_bl
Rbb_88_52 bitb_88_52 bitb_88_53 R_bl
Cb_88_52 bit_88_52 gnd C_bl
Cbb_88_52 bitb_88_52 gnd C_bl
Rb_88_53 bit_88_53 bit_88_54 R_bl
Rbb_88_53 bitb_88_53 bitb_88_54 R_bl
Cb_88_53 bit_88_53 gnd C_bl
Cbb_88_53 bitb_88_53 gnd C_bl
Rb_88_54 bit_88_54 bit_88_55 R_bl
Rbb_88_54 bitb_88_54 bitb_88_55 R_bl
Cb_88_54 bit_88_54 gnd C_bl
Cbb_88_54 bitb_88_54 gnd C_bl
Rb_88_55 bit_88_55 bit_88_56 R_bl
Rbb_88_55 bitb_88_55 bitb_88_56 R_bl
Cb_88_55 bit_88_55 gnd C_bl
Cbb_88_55 bitb_88_55 gnd C_bl
Rb_88_56 bit_88_56 bit_88_57 R_bl
Rbb_88_56 bitb_88_56 bitb_88_57 R_bl
Cb_88_56 bit_88_56 gnd C_bl
Cbb_88_56 bitb_88_56 gnd C_bl
Rb_88_57 bit_88_57 bit_88_58 R_bl
Rbb_88_57 bitb_88_57 bitb_88_58 R_bl
Cb_88_57 bit_88_57 gnd C_bl
Cbb_88_57 bitb_88_57 gnd C_bl
Rb_88_58 bit_88_58 bit_88_59 R_bl
Rbb_88_58 bitb_88_58 bitb_88_59 R_bl
Cb_88_58 bit_88_58 gnd C_bl
Cbb_88_58 bitb_88_58 gnd C_bl
Rb_88_59 bit_88_59 bit_88_60 R_bl
Rbb_88_59 bitb_88_59 bitb_88_60 R_bl
Cb_88_59 bit_88_59 gnd C_bl
Cbb_88_59 bitb_88_59 gnd C_bl
Rb_88_60 bit_88_60 bit_88_61 R_bl
Rbb_88_60 bitb_88_60 bitb_88_61 R_bl
Cb_88_60 bit_88_60 gnd C_bl
Cbb_88_60 bitb_88_60 gnd C_bl
Rb_88_61 bit_88_61 bit_88_62 R_bl
Rbb_88_61 bitb_88_61 bitb_88_62 R_bl
Cb_88_61 bit_88_61 gnd C_bl
Cbb_88_61 bitb_88_61 gnd C_bl
Rb_88_62 bit_88_62 bit_88_63 R_bl
Rbb_88_62 bitb_88_62 bitb_88_63 R_bl
Cb_88_62 bit_88_62 gnd C_bl
Cbb_88_62 bitb_88_62 gnd C_bl
Rb_88_63 bit_88_63 bit_88_64 R_bl
Rbb_88_63 bitb_88_63 bitb_88_64 R_bl
Cb_88_63 bit_88_63 gnd C_bl
Cbb_88_63 bitb_88_63 gnd C_bl
Rb_88_64 bit_88_64 bit_88_65 R_bl
Rbb_88_64 bitb_88_64 bitb_88_65 R_bl
Cb_88_64 bit_88_64 gnd C_bl
Cbb_88_64 bitb_88_64 gnd C_bl
Rb_88_65 bit_88_65 bit_88_66 R_bl
Rbb_88_65 bitb_88_65 bitb_88_66 R_bl
Cb_88_65 bit_88_65 gnd C_bl
Cbb_88_65 bitb_88_65 gnd C_bl
Rb_88_66 bit_88_66 bit_88_67 R_bl
Rbb_88_66 bitb_88_66 bitb_88_67 R_bl
Cb_88_66 bit_88_66 gnd C_bl
Cbb_88_66 bitb_88_66 gnd C_bl
Rb_88_67 bit_88_67 bit_88_68 R_bl
Rbb_88_67 bitb_88_67 bitb_88_68 R_bl
Cb_88_67 bit_88_67 gnd C_bl
Cbb_88_67 bitb_88_67 gnd C_bl
Rb_88_68 bit_88_68 bit_88_69 R_bl
Rbb_88_68 bitb_88_68 bitb_88_69 R_bl
Cb_88_68 bit_88_68 gnd C_bl
Cbb_88_68 bitb_88_68 gnd C_bl
Rb_88_69 bit_88_69 bit_88_70 R_bl
Rbb_88_69 bitb_88_69 bitb_88_70 R_bl
Cb_88_69 bit_88_69 gnd C_bl
Cbb_88_69 bitb_88_69 gnd C_bl
Rb_88_70 bit_88_70 bit_88_71 R_bl
Rbb_88_70 bitb_88_70 bitb_88_71 R_bl
Cb_88_70 bit_88_70 gnd C_bl
Cbb_88_70 bitb_88_70 gnd C_bl
Rb_88_71 bit_88_71 bit_88_72 R_bl
Rbb_88_71 bitb_88_71 bitb_88_72 R_bl
Cb_88_71 bit_88_71 gnd C_bl
Cbb_88_71 bitb_88_71 gnd C_bl
Rb_88_72 bit_88_72 bit_88_73 R_bl
Rbb_88_72 bitb_88_72 bitb_88_73 R_bl
Cb_88_72 bit_88_72 gnd C_bl
Cbb_88_72 bitb_88_72 gnd C_bl
Rb_88_73 bit_88_73 bit_88_74 R_bl
Rbb_88_73 bitb_88_73 bitb_88_74 R_bl
Cb_88_73 bit_88_73 gnd C_bl
Cbb_88_73 bitb_88_73 gnd C_bl
Rb_88_74 bit_88_74 bit_88_75 R_bl
Rbb_88_74 bitb_88_74 bitb_88_75 R_bl
Cb_88_74 bit_88_74 gnd C_bl
Cbb_88_74 bitb_88_74 gnd C_bl
Rb_88_75 bit_88_75 bit_88_76 R_bl
Rbb_88_75 bitb_88_75 bitb_88_76 R_bl
Cb_88_75 bit_88_75 gnd C_bl
Cbb_88_75 bitb_88_75 gnd C_bl
Rb_88_76 bit_88_76 bit_88_77 R_bl
Rbb_88_76 bitb_88_76 bitb_88_77 R_bl
Cb_88_76 bit_88_76 gnd C_bl
Cbb_88_76 bitb_88_76 gnd C_bl
Rb_88_77 bit_88_77 bit_88_78 R_bl
Rbb_88_77 bitb_88_77 bitb_88_78 R_bl
Cb_88_77 bit_88_77 gnd C_bl
Cbb_88_77 bitb_88_77 gnd C_bl
Rb_88_78 bit_88_78 bit_88_79 R_bl
Rbb_88_78 bitb_88_78 bitb_88_79 R_bl
Cb_88_78 bit_88_78 gnd C_bl
Cbb_88_78 bitb_88_78 gnd C_bl
Rb_88_79 bit_88_79 bit_88_80 R_bl
Rbb_88_79 bitb_88_79 bitb_88_80 R_bl
Cb_88_79 bit_88_79 gnd C_bl
Cbb_88_79 bitb_88_79 gnd C_bl
Rb_88_80 bit_88_80 bit_88_81 R_bl
Rbb_88_80 bitb_88_80 bitb_88_81 R_bl
Cb_88_80 bit_88_80 gnd C_bl
Cbb_88_80 bitb_88_80 gnd C_bl
Rb_88_81 bit_88_81 bit_88_82 R_bl
Rbb_88_81 bitb_88_81 bitb_88_82 R_bl
Cb_88_81 bit_88_81 gnd C_bl
Cbb_88_81 bitb_88_81 gnd C_bl
Rb_88_82 bit_88_82 bit_88_83 R_bl
Rbb_88_82 bitb_88_82 bitb_88_83 R_bl
Cb_88_82 bit_88_82 gnd C_bl
Cbb_88_82 bitb_88_82 gnd C_bl
Rb_88_83 bit_88_83 bit_88_84 R_bl
Rbb_88_83 bitb_88_83 bitb_88_84 R_bl
Cb_88_83 bit_88_83 gnd C_bl
Cbb_88_83 bitb_88_83 gnd C_bl
Rb_88_84 bit_88_84 bit_88_85 R_bl
Rbb_88_84 bitb_88_84 bitb_88_85 R_bl
Cb_88_84 bit_88_84 gnd C_bl
Cbb_88_84 bitb_88_84 gnd C_bl
Rb_88_85 bit_88_85 bit_88_86 R_bl
Rbb_88_85 bitb_88_85 bitb_88_86 R_bl
Cb_88_85 bit_88_85 gnd C_bl
Cbb_88_85 bitb_88_85 gnd C_bl
Rb_88_86 bit_88_86 bit_88_87 R_bl
Rbb_88_86 bitb_88_86 bitb_88_87 R_bl
Cb_88_86 bit_88_86 gnd C_bl
Cbb_88_86 bitb_88_86 gnd C_bl
Rb_88_87 bit_88_87 bit_88_88 R_bl
Rbb_88_87 bitb_88_87 bitb_88_88 R_bl
Cb_88_87 bit_88_87 gnd C_bl
Cbb_88_87 bitb_88_87 gnd C_bl
Rb_88_88 bit_88_88 bit_88_89 R_bl
Rbb_88_88 bitb_88_88 bitb_88_89 R_bl
Cb_88_88 bit_88_88 gnd C_bl
Cbb_88_88 bitb_88_88 gnd C_bl
Rb_88_89 bit_88_89 bit_88_90 R_bl
Rbb_88_89 bitb_88_89 bitb_88_90 R_bl
Cb_88_89 bit_88_89 gnd C_bl
Cbb_88_89 bitb_88_89 gnd C_bl
Rb_88_90 bit_88_90 bit_88_91 R_bl
Rbb_88_90 bitb_88_90 bitb_88_91 R_bl
Cb_88_90 bit_88_90 gnd C_bl
Cbb_88_90 bitb_88_90 gnd C_bl
Rb_88_91 bit_88_91 bit_88_92 R_bl
Rbb_88_91 bitb_88_91 bitb_88_92 R_bl
Cb_88_91 bit_88_91 gnd C_bl
Cbb_88_91 bitb_88_91 gnd C_bl
Rb_88_92 bit_88_92 bit_88_93 R_bl
Rbb_88_92 bitb_88_92 bitb_88_93 R_bl
Cb_88_92 bit_88_92 gnd C_bl
Cbb_88_92 bitb_88_92 gnd C_bl
Rb_88_93 bit_88_93 bit_88_94 R_bl
Rbb_88_93 bitb_88_93 bitb_88_94 R_bl
Cb_88_93 bit_88_93 gnd C_bl
Cbb_88_93 bitb_88_93 gnd C_bl
Rb_88_94 bit_88_94 bit_88_95 R_bl
Rbb_88_94 bitb_88_94 bitb_88_95 R_bl
Cb_88_94 bit_88_94 gnd C_bl
Cbb_88_94 bitb_88_94 gnd C_bl
Rb_88_95 bit_88_95 bit_88_96 R_bl
Rbb_88_95 bitb_88_95 bitb_88_96 R_bl
Cb_88_95 bit_88_95 gnd C_bl
Cbb_88_95 bitb_88_95 gnd C_bl
Rb_88_96 bit_88_96 bit_88_97 R_bl
Rbb_88_96 bitb_88_96 bitb_88_97 R_bl
Cb_88_96 bit_88_96 gnd C_bl
Cbb_88_96 bitb_88_96 gnd C_bl
Rb_88_97 bit_88_97 bit_88_98 R_bl
Rbb_88_97 bitb_88_97 bitb_88_98 R_bl
Cb_88_97 bit_88_97 gnd C_bl
Cbb_88_97 bitb_88_97 gnd C_bl
Rb_88_98 bit_88_98 bit_88_99 R_bl
Rbb_88_98 bitb_88_98 bitb_88_99 R_bl
Cb_88_98 bit_88_98 gnd C_bl
Cbb_88_98 bitb_88_98 gnd C_bl
Rb_88_99 bit_88_99 bit_88_100 R_bl
Rbb_88_99 bitb_88_99 bitb_88_100 R_bl
Cb_88_99 bit_88_99 gnd C_bl
Cbb_88_99 bitb_88_99 gnd C_bl
Rb_89_0 bit_89_0 bit_89_1 R_bl
Rbb_89_0 bitb_89_0 bitb_89_1 R_bl
Cb_89_0 bit_89_0 gnd C_bl
Cbb_89_0 bitb_89_0 gnd C_bl
Rb_89_1 bit_89_1 bit_89_2 R_bl
Rbb_89_1 bitb_89_1 bitb_89_2 R_bl
Cb_89_1 bit_89_1 gnd C_bl
Cbb_89_1 bitb_89_1 gnd C_bl
Rb_89_2 bit_89_2 bit_89_3 R_bl
Rbb_89_2 bitb_89_2 bitb_89_3 R_bl
Cb_89_2 bit_89_2 gnd C_bl
Cbb_89_2 bitb_89_2 gnd C_bl
Rb_89_3 bit_89_3 bit_89_4 R_bl
Rbb_89_3 bitb_89_3 bitb_89_4 R_bl
Cb_89_3 bit_89_3 gnd C_bl
Cbb_89_3 bitb_89_3 gnd C_bl
Rb_89_4 bit_89_4 bit_89_5 R_bl
Rbb_89_4 bitb_89_4 bitb_89_5 R_bl
Cb_89_4 bit_89_4 gnd C_bl
Cbb_89_4 bitb_89_4 gnd C_bl
Rb_89_5 bit_89_5 bit_89_6 R_bl
Rbb_89_5 bitb_89_5 bitb_89_6 R_bl
Cb_89_5 bit_89_5 gnd C_bl
Cbb_89_5 bitb_89_5 gnd C_bl
Rb_89_6 bit_89_6 bit_89_7 R_bl
Rbb_89_6 bitb_89_6 bitb_89_7 R_bl
Cb_89_6 bit_89_6 gnd C_bl
Cbb_89_6 bitb_89_6 gnd C_bl
Rb_89_7 bit_89_7 bit_89_8 R_bl
Rbb_89_7 bitb_89_7 bitb_89_8 R_bl
Cb_89_7 bit_89_7 gnd C_bl
Cbb_89_7 bitb_89_7 gnd C_bl
Rb_89_8 bit_89_8 bit_89_9 R_bl
Rbb_89_8 bitb_89_8 bitb_89_9 R_bl
Cb_89_8 bit_89_8 gnd C_bl
Cbb_89_8 bitb_89_8 gnd C_bl
Rb_89_9 bit_89_9 bit_89_10 R_bl
Rbb_89_9 bitb_89_9 bitb_89_10 R_bl
Cb_89_9 bit_89_9 gnd C_bl
Cbb_89_9 bitb_89_9 gnd C_bl
Rb_89_10 bit_89_10 bit_89_11 R_bl
Rbb_89_10 bitb_89_10 bitb_89_11 R_bl
Cb_89_10 bit_89_10 gnd C_bl
Cbb_89_10 bitb_89_10 gnd C_bl
Rb_89_11 bit_89_11 bit_89_12 R_bl
Rbb_89_11 bitb_89_11 bitb_89_12 R_bl
Cb_89_11 bit_89_11 gnd C_bl
Cbb_89_11 bitb_89_11 gnd C_bl
Rb_89_12 bit_89_12 bit_89_13 R_bl
Rbb_89_12 bitb_89_12 bitb_89_13 R_bl
Cb_89_12 bit_89_12 gnd C_bl
Cbb_89_12 bitb_89_12 gnd C_bl
Rb_89_13 bit_89_13 bit_89_14 R_bl
Rbb_89_13 bitb_89_13 bitb_89_14 R_bl
Cb_89_13 bit_89_13 gnd C_bl
Cbb_89_13 bitb_89_13 gnd C_bl
Rb_89_14 bit_89_14 bit_89_15 R_bl
Rbb_89_14 bitb_89_14 bitb_89_15 R_bl
Cb_89_14 bit_89_14 gnd C_bl
Cbb_89_14 bitb_89_14 gnd C_bl
Rb_89_15 bit_89_15 bit_89_16 R_bl
Rbb_89_15 bitb_89_15 bitb_89_16 R_bl
Cb_89_15 bit_89_15 gnd C_bl
Cbb_89_15 bitb_89_15 gnd C_bl
Rb_89_16 bit_89_16 bit_89_17 R_bl
Rbb_89_16 bitb_89_16 bitb_89_17 R_bl
Cb_89_16 bit_89_16 gnd C_bl
Cbb_89_16 bitb_89_16 gnd C_bl
Rb_89_17 bit_89_17 bit_89_18 R_bl
Rbb_89_17 bitb_89_17 bitb_89_18 R_bl
Cb_89_17 bit_89_17 gnd C_bl
Cbb_89_17 bitb_89_17 gnd C_bl
Rb_89_18 bit_89_18 bit_89_19 R_bl
Rbb_89_18 bitb_89_18 bitb_89_19 R_bl
Cb_89_18 bit_89_18 gnd C_bl
Cbb_89_18 bitb_89_18 gnd C_bl
Rb_89_19 bit_89_19 bit_89_20 R_bl
Rbb_89_19 bitb_89_19 bitb_89_20 R_bl
Cb_89_19 bit_89_19 gnd C_bl
Cbb_89_19 bitb_89_19 gnd C_bl
Rb_89_20 bit_89_20 bit_89_21 R_bl
Rbb_89_20 bitb_89_20 bitb_89_21 R_bl
Cb_89_20 bit_89_20 gnd C_bl
Cbb_89_20 bitb_89_20 gnd C_bl
Rb_89_21 bit_89_21 bit_89_22 R_bl
Rbb_89_21 bitb_89_21 bitb_89_22 R_bl
Cb_89_21 bit_89_21 gnd C_bl
Cbb_89_21 bitb_89_21 gnd C_bl
Rb_89_22 bit_89_22 bit_89_23 R_bl
Rbb_89_22 bitb_89_22 bitb_89_23 R_bl
Cb_89_22 bit_89_22 gnd C_bl
Cbb_89_22 bitb_89_22 gnd C_bl
Rb_89_23 bit_89_23 bit_89_24 R_bl
Rbb_89_23 bitb_89_23 bitb_89_24 R_bl
Cb_89_23 bit_89_23 gnd C_bl
Cbb_89_23 bitb_89_23 gnd C_bl
Rb_89_24 bit_89_24 bit_89_25 R_bl
Rbb_89_24 bitb_89_24 bitb_89_25 R_bl
Cb_89_24 bit_89_24 gnd C_bl
Cbb_89_24 bitb_89_24 gnd C_bl
Rb_89_25 bit_89_25 bit_89_26 R_bl
Rbb_89_25 bitb_89_25 bitb_89_26 R_bl
Cb_89_25 bit_89_25 gnd C_bl
Cbb_89_25 bitb_89_25 gnd C_bl
Rb_89_26 bit_89_26 bit_89_27 R_bl
Rbb_89_26 bitb_89_26 bitb_89_27 R_bl
Cb_89_26 bit_89_26 gnd C_bl
Cbb_89_26 bitb_89_26 gnd C_bl
Rb_89_27 bit_89_27 bit_89_28 R_bl
Rbb_89_27 bitb_89_27 bitb_89_28 R_bl
Cb_89_27 bit_89_27 gnd C_bl
Cbb_89_27 bitb_89_27 gnd C_bl
Rb_89_28 bit_89_28 bit_89_29 R_bl
Rbb_89_28 bitb_89_28 bitb_89_29 R_bl
Cb_89_28 bit_89_28 gnd C_bl
Cbb_89_28 bitb_89_28 gnd C_bl
Rb_89_29 bit_89_29 bit_89_30 R_bl
Rbb_89_29 bitb_89_29 bitb_89_30 R_bl
Cb_89_29 bit_89_29 gnd C_bl
Cbb_89_29 bitb_89_29 gnd C_bl
Rb_89_30 bit_89_30 bit_89_31 R_bl
Rbb_89_30 bitb_89_30 bitb_89_31 R_bl
Cb_89_30 bit_89_30 gnd C_bl
Cbb_89_30 bitb_89_30 gnd C_bl
Rb_89_31 bit_89_31 bit_89_32 R_bl
Rbb_89_31 bitb_89_31 bitb_89_32 R_bl
Cb_89_31 bit_89_31 gnd C_bl
Cbb_89_31 bitb_89_31 gnd C_bl
Rb_89_32 bit_89_32 bit_89_33 R_bl
Rbb_89_32 bitb_89_32 bitb_89_33 R_bl
Cb_89_32 bit_89_32 gnd C_bl
Cbb_89_32 bitb_89_32 gnd C_bl
Rb_89_33 bit_89_33 bit_89_34 R_bl
Rbb_89_33 bitb_89_33 bitb_89_34 R_bl
Cb_89_33 bit_89_33 gnd C_bl
Cbb_89_33 bitb_89_33 gnd C_bl
Rb_89_34 bit_89_34 bit_89_35 R_bl
Rbb_89_34 bitb_89_34 bitb_89_35 R_bl
Cb_89_34 bit_89_34 gnd C_bl
Cbb_89_34 bitb_89_34 gnd C_bl
Rb_89_35 bit_89_35 bit_89_36 R_bl
Rbb_89_35 bitb_89_35 bitb_89_36 R_bl
Cb_89_35 bit_89_35 gnd C_bl
Cbb_89_35 bitb_89_35 gnd C_bl
Rb_89_36 bit_89_36 bit_89_37 R_bl
Rbb_89_36 bitb_89_36 bitb_89_37 R_bl
Cb_89_36 bit_89_36 gnd C_bl
Cbb_89_36 bitb_89_36 gnd C_bl
Rb_89_37 bit_89_37 bit_89_38 R_bl
Rbb_89_37 bitb_89_37 bitb_89_38 R_bl
Cb_89_37 bit_89_37 gnd C_bl
Cbb_89_37 bitb_89_37 gnd C_bl
Rb_89_38 bit_89_38 bit_89_39 R_bl
Rbb_89_38 bitb_89_38 bitb_89_39 R_bl
Cb_89_38 bit_89_38 gnd C_bl
Cbb_89_38 bitb_89_38 gnd C_bl
Rb_89_39 bit_89_39 bit_89_40 R_bl
Rbb_89_39 bitb_89_39 bitb_89_40 R_bl
Cb_89_39 bit_89_39 gnd C_bl
Cbb_89_39 bitb_89_39 gnd C_bl
Rb_89_40 bit_89_40 bit_89_41 R_bl
Rbb_89_40 bitb_89_40 bitb_89_41 R_bl
Cb_89_40 bit_89_40 gnd C_bl
Cbb_89_40 bitb_89_40 gnd C_bl
Rb_89_41 bit_89_41 bit_89_42 R_bl
Rbb_89_41 bitb_89_41 bitb_89_42 R_bl
Cb_89_41 bit_89_41 gnd C_bl
Cbb_89_41 bitb_89_41 gnd C_bl
Rb_89_42 bit_89_42 bit_89_43 R_bl
Rbb_89_42 bitb_89_42 bitb_89_43 R_bl
Cb_89_42 bit_89_42 gnd C_bl
Cbb_89_42 bitb_89_42 gnd C_bl
Rb_89_43 bit_89_43 bit_89_44 R_bl
Rbb_89_43 bitb_89_43 bitb_89_44 R_bl
Cb_89_43 bit_89_43 gnd C_bl
Cbb_89_43 bitb_89_43 gnd C_bl
Rb_89_44 bit_89_44 bit_89_45 R_bl
Rbb_89_44 bitb_89_44 bitb_89_45 R_bl
Cb_89_44 bit_89_44 gnd C_bl
Cbb_89_44 bitb_89_44 gnd C_bl
Rb_89_45 bit_89_45 bit_89_46 R_bl
Rbb_89_45 bitb_89_45 bitb_89_46 R_bl
Cb_89_45 bit_89_45 gnd C_bl
Cbb_89_45 bitb_89_45 gnd C_bl
Rb_89_46 bit_89_46 bit_89_47 R_bl
Rbb_89_46 bitb_89_46 bitb_89_47 R_bl
Cb_89_46 bit_89_46 gnd C_bl
Cbb_89_46 bitb_89_46 gnd C_bl
Rb_89_47 bit_89_47 bit_89_48 R_bl
Rbb_89_47 bitb_89_47 bitb_89_48 R_bl
Cb_89_47 bit_89_47 gnd C_bl
Cbb_89_47 bitb_89_47 gnd C_bl
Rb_89_48 bit_89_48 bit_89_49 R_bl
Rbb_89_48 bitb_89_48 bitb_89_49 R_bl
Cb_89_48 bit_89_48 gnd C_bl
Cbb_89_48 bitb_89_48 gnd C_bl
Rb_89_49 bit_89_49 bit_89_50 R_bl
Rbb_89_49 bitb_89_49 bitb_89_50 R_bl
Cb_89_49 bit_89_49 gnd C_bl
Cbb_89_49 bitb_89_49 gnd C_bl
Rb_89_50 bit_89_50 bit_89_51 R_bl
Rbb_89_50 bitb_89_50 bitb_89_51 R_bl
Cb_89_50 bit_89_50 gnd C_bl
Cbb_89_50 bitb_89_50 gnd C_bl
Rb_89_51 bit_89_51 bit_89_52 R_bl
Rbb_89_51 bitb_89_51 bitb_89_52 R_bl
Cb_89_51 bit_89_51 gnd C_bl
Cbb_89_51 bitb_89_51 gnd C_bl
Rb_89_52 bit_89_52 bit_89_53 R_bl
Rbb_89_52 bitb_89_52 bitb_89_53 R_bl
Cb_89_52 bit_89_52 gnd C_bl
Cbb_89_52 bitb_89_52 gnd C_bl
Rb_89_53 bit_89_53 bit_89_54 R_bl
Rbb_89_53 bitb_89_53 bitb_89_54 R_bl
Cb_89_53 bit_89_53 gnd C_bl
Cbb_89_53 bitb_89_53 gnd C_bl
Rb_89_54 bit_89_54 bit_89_55 R_bl
Rbb_89_54 bitb_89_54 bitb_89_55 R_bl
Cb_89_54 bit_89_54 gnd C_bl
Cbb_89_54 bitb_89_54 gnd C_bl
Rb_89_55 bit_89_55 bit_89_56 R_bl
Rbb_89_55 bitb_89_55 bitb_89_56 R_bl
Cb_89_55 bit_89_55 gnd C_bl
Cbb_89_55 bitb_89_55 gnd C_bl
Rb_89_56 bit_89_56 bit_89_57 R_bl
Rbb_89_56 bitb_89_56 bitb_89_57 R_bl
Cb_89_56 bit_89_56 gnd C_bl
Cbb_89_56 bitb_89_56 gnd C_bl
Rb_89_57 bit_89_57 bit_89_58 R_bl
Rbb_89_57 bitb_89_57 bitb_89_58 R_bl
Cb_89_57 bit_89_57 gnd C_bl
Cbb_89_57 bitb_89_57 gnd C_bl
Rb_89_58 bit_89_58 bit_89_59 R_bl
Rbb_89_58 bitb_89_58 bitb_89_59 R_bl
Cb_89_58 bit_89_58 gnd C_bl
Cbb_89_58 bitb_89_58 gnd C_bl
Rb_89_59 bit_89_59 bit_89_60 R_bl
Rbb_89_59 bitb_89_59 bitb_89_60 R_bl
Cb_89_59 bit_89_59 gnd C_bl
Cbb_89_59 bitb_89_59 gnd C_bl
Rb_89_60 bit_89_60 bit_89_61 R_bl
Rbb_89_60 bitb_89_60 bitb_89_61 R_bl
Cb_89_60 bit_89_60 gnd C_bl
Cbb_89_60 bitb_89_60 gnd C_bl
Rb_89_61 bit_89_61 bit_89_62 R_bl
Rbb_89_61 bitb_89_61 bitb_89_62 R_bl
Cb_89_61 bit_89_61 gnd C_bl
Cbb_89_61 bitb_89_61 gnd C_bl
Rb_89_62 bit_89_62 bit_89_63 R_bl
Rbb_89_62 bitb_89_62 bitb_89_63 R_bl
Cb_89_62 bit_89_62 gnd C_bl
Cbb_89_62 bitb_89_62 gnd C_bl
Rb_89_63 bit_89_63 bit_89_64 R_bl
Rbb_89_63 bitb_89_63 bitb_89_64 R_bl
Cb_89_63 bit_89_63 gnd C_bl
Cbb_89_63 bitb_89_63 gnd C_bl
Rb_89_64 bit_89_64 bit_89_65 R_bl
Rbb_89_64 bitb_89_64 bitb_89_65 R_bl
Cb_89_64 bit_89_64 gnd C_bl
Cbb_89_64 bitb_89_64 gnd C_bl
Rb_89_65 bit_89_65 bit_89_66 R_bl
Rbb_89_65 bitb_89_65 bitb_89_66 R_bl
Cb_89_65 bit_89_65 gnd C_bl
Cbb_89_65 bitb_89_65 gnd C_bl
Rb_89_66 bit_89_66 bit_89_67 R_bl
Rbb_89_66 bitb_89_66 bitb_89_67 R_bl
Cb_89_66 bit_89_66 gnd C_bl
Cbb_89_66 bitb_89_66 gnd C_bl
Rb_89_67 bit_89_67 bit_89_68 R_bl
Rbb_89_67 bitb_89_67 bitb_89_68 R_bl
Cb_89_67 bit_89_67 gnd C_bl
Cbb_89_67 bitb_89_67 gnd C_bl
Rb_89_68 bit_89_68 bit_89_69 R_bl
Rbb_89_68 bitb_89_68 bitb_89_69 R_bl
Cb_89_68 bit_89_68 gnd C_bl
Cbb_89_68 bitb_89_68 gnd C_bl
Rb_89_69 bit_89_69 bit_89_70 R_bl
Rbb_89_69 bitb_89_69 bitb_89_70 R_bl
Cb_89_69 bit_89_69 gnd C_bl
Cbb_89_69 bitb_89_69 gnd C_bl
Rb_89_70 bit_89_70 bit_89_71 R_bl
Rbb_89_70 bitb_89_70 bitb_89_71 R_bl
Cb_89_70 bit_89_70 gnd C_bl
Cbb_89_70 bitb_89_70 gnd C_bl
Rb_89_71 bit_89_71 bit_89_72 R_bl
Rbb_89_71 bitb_89_71 bitb_89_72 R_bl
Cb_89_71 bit_89_71 gnd C_bl
Cbb_89_71 bitb_89_71 gnd C_bl
Rb_89_72 bit_89_72 bit_89_73 R_bl
Rbb_89_72 bitb_89_72 bitb_89_73 R_bl
Cb_89_72 bit_89_72 gnd C_bl
Cbb_89_72 bitb_89_72 gnd C_bl
Rb_89_73 bit_89_73 bit_89_74 R_bl
Rbb_89_73 bitb_89_73 bitb_89_74 R_bl
Cb_89_73 bit_89_73 gnd C_bl
Cbb_89_73 bitb_89_73 gnd C_bl
Rb_89_74 bit_89_74 bit_89_75 R_bl
Rbb_89_74 bitb_89_74 bitb_89_75 R_bl
Cb_89_74 bit_89_74 gnd C_bl
Cbb_89_74 bitb_89_74 gnd C_bl
Rb_89_75 bit_89_75 bit_89_76 R_bl
Rbb_89_75 bitb_89_75 bitb_89_76 R_bl
Cb_89_75 bit_89_75 gnd C_bl
Cbb_89_75 bitb_89_75 gnd C_bl
Rb_89_76 bit_89_76 bit_89_77 R_bl
Rbb_89_76 bitb_89_76 bitb_89_77 R_bl
Cb_89_76 bit_89_76 gnd C_bl
Cbb_89_76 bitb_89_76 gnd C_bl
Rb_89_77 bit_89_77 bit_89_78 R_bl
Rbb_89_77 bitb_89_77 bitb_89_78 R_bl
Cb_89_77 bit_89_77 gnd C_bl
Cbb_89_77 bitb_89_77 gnd C_bl
Rb_89_78 bit_89_78 bit_89_79 R_bl
Rbb_89_78 bitb_89_78 bitb_89_79 R_bl
Cb_89_78 bit_89_78 gnd C_bl
Cbb_89_78 bitb_89_78 gnd C_bl
Rb_89_79 bit_89_79 bit_89_80 R_bl
Rbb_89_79 bitb_89_79 bitb_89_80 R_bl
Cb_89_79 bit_89_79 gnd C_bl
Cbb_89_79 bitb_89_79 gnd C_bl
Rb_89_80 bit_89_80 bit_89_81 R_bl
Rbb_89_80 bitb_89_80 bitb_89_81 R_bl
Cb_89_80 bit_89_80 gnd C_bl
Cbb_89_80 bitb_89_80 gnd C_bl
Rb_89_81 bit_89_81 bit_89_82 R_bl
Rbb_89_81 bitb_89_81 bitb_89_82 R_bl
Cb_89_81 bit_89_81 gnd C_bl
Cbb_89_81 bitb_89_81 gnd C_bl
Rb_89_82 bit_89_82 bit_89_83 R_bl
Rbb_89_82 bitb_89_82 bitb_89_83 R_bl
Cb_89_82 bit_89_82 gnd C_bl
Cbb_89_82 bitb_89_82 gnd C_bl
Rb_89_83 bit_89_83 bit_89_84 R_bl
Rbb_89_83 bitb_89_83 bitb_89_84 R_bl
Cb_89_83 bit_89_83 gnd C_bl
Cbb_89_83 bitb_89_83 gnd C_bl
Rb_89_84 bit_89_84 bit_89_85 R_bl
Rbb_89_84 bitb_89_84 bitb_89_85 R_bl
Cb_89_84 bit_89_84 gnd C_bl
Cbb_89_84 bitb_89_84 gnd C_bl
Rb_89_85 bit_89_85 bit_89_86 R_bl
Rbb_89_85 bitb_89_85 bitb_89_86 R_bl
Cb_89_85 bit_89_85 gnd C_bl
Cbb_89_85 bitb_89_85 gnd C_bl
Rb_89_86 bit_89_86 bit_89_87 R_bl
Rbb_89_86 bitb_89_86 bitb_89_87 R_bl
Cb_89_86 bit_89_86 gnd C_bl
Cbb_89_86 bitb_89_86 gnd C_bl
Rb_89_87 bit_89_87 bit_89_88 R_bl
Rbb_89_87 bitb_89_87 bitb_89_88 R_bl
Cb_89_87 bit_89_87 gnd C_bl
Cbb_89_87 bitb_89_87 gnd C_bl
Rb_89_88 bit_89_88 bit_89_89 R_bl
Rbb_89_88 bitb_89_88 bitb_89_89 R_bl
Cb_89_88 bit_89_88 gnd C_bl
Cbb_89_88 bitb_89_88 gnd C_bl
Rb_89_89 bit_89_89 bit_89_90 R_bl
Rbb_89_89 bitb_89_89 bitb_89_90 R_bl
Cb_89_89 bit_89_89 gnd C_bl
Cbb_89_89 bitb_89_89 gnd C_bl
Rb_89_90 bit_89_90 bit_89_91 R_bl
Rbb_89_90 bitb_89_90 bitb_89_91 R_bl
Cb_89_90 bit_89_90 gnd C_bl
Cbb_89_90 bitb_89_90 gnd C_bl
Rb_89_91 bit_89_91 bit_89_92 R_bl
Rbb_89_91 bitb_89_91 bitb_89_92 R_bl
Cb_89_91 bit_89_91 gnd C_bl
Cbb_89_91 bitb_89_91 gnd C_bl
Rb_89_92 bit_89_92 bit_89_93 R_bl
Rbb_89_92 bitb_89_92 bitb_89_93 R_bl
Cb_89_92 bit_89_92 gnd C_bl
Cbb_89_92 bitb_89_92 gnd C_bl
Rb_89_93 bit_89_93 bit_89_94 R_bl
Rbb_89_93 bitb_89_93 bitb_89_94 R_bl
Cb_89_93 bit_89_93 gnd C_bl
Cbb_89_93 bitb_89_93 gnd C_bl
Rb_89_94 bit_89_94 bit_89_95 R_bl
Rbb_89_94 bitb_89_94 bitb_89_95 R_bl
Cb_89_94 bit_89_94 gnd C_bl
Cbb_89_94 bitb_89_94 gnd C_bl
Rb_89_95 bit_89_95 bit_89_96 R_bl
Rbb_89_95 bitb_89_95 bitb_89_96 R_bl
Cb_89_95 bit_89_95 gnd C_bl
Cbb_89_95 bitb_89_95 gnd C_bl
Rb_89_96 bit_89_96 bit_89_97 R_bl
Rbb_89_96 bitb_89_96 bitb_89_97 R_bl
Cb_89_96 bit_89_96 gnd C_bl
Cbb_89_96 bitb_89_96 gnd C_bl
Rb_89_97 bit_89_97 bit_89_98 R_bl
Rbb_89_97 bitb_89_97 bitb_89_98 R_bl
Cb_89_97 bit_89_97 gnd C_bl
Cbb_89_97 bitb_89_97 gnd C_bl
Rb_89_98 bit_89_98 bit_89_99 R_bl
Rbb_89_98 bitb_89_98 bitb_89_99 R_bl
Cb_89_98 bit_89_98 gnd C_bl
Cbb_89_98 bitb_89_98 gnd C_bl
Rb_89_99 bit_89_99 bit_89_100 R_bl
Rbb_89_99 bitb_89_99 bitb_89_100 R_bl
Cb_89_99 bit_89_99 gnd C_bl
Cbb_89_99 bitb_89_99 gnd C_bl
Rb_90_0 bit_90_0 bit_90_1 R_bl
Rbb_90_0 bitb_90_0 bitb_90_1 R_bl
Cb_90_0 bit_90_0 gnd C_bl
Cbb_90_0 bitb_90_0 gnd C_bl
Rb_90_1 bit_90_1 bit_90_2 R_bl
Rbb_90_1 bitb_90_1 bitb_90_2 R_bl
Cb_90_1 bit_90_1 gnd C_bl
Cbb_90_1 bitb_90_1 gnd C_bl
Rb_90_2 bit_90_2 bit_90_3 R_bl
Rbb_90_2 bitb_90_2 bitb_90_3 R_bl
Cb_90_2 bit_90_2 gnd C_bl
Cbb_90_2 bitb_90_2 gnd C_bl
Rb_90_3 bit_90_3 bit_90_4 R_bl
Rbb_90_3 bitb_90_3 bitb_90_4 R_bl
Cb_90_3 bit_90_3 gnd C_bl
Cbb_90_3 bitb_90_3 gnd C_bl
Rb_90_4 bit_90_4 bit_90_5 R_bl
Rbb_90_4 bitb_90_4 bitb_90_5 R_bl
Cb_90_4 bit_90_4 gnd C_bl
Cbb_90_4 bitb_90_4 gnd C_bl
Rb_90_5 bit_90_5 bit_90_6 R_bl
Rbb_90_5 bitb_90_5 bitb_90_6 R_bl
Cb_90_5 bit_90_5 gnd C_bl
Cbb_90_5 bitb_90_5 gnd C_bl
Rb_90_6 bit_90_6 bit_90_7 R_bl
Rbb_90_6 bitb_90_6 bitb_90_7 R_bl
Cb_90_6 bit_90_6 gnd C_bl
Cbb_90_6 bitb_90_6 gnd C_bl
Rb_90_7 bit_90_7 bit_90_8 R_bl
Rbb_90_7 bitb_90_7 bitb_90_8 R_bl
Cb_90_7 bit_90_7 gnd C_bl
Cbb_90_7 bitb_90_7 gnd C_bl
Rb_90_8 bit_90_8 bit_90_9 R_bl
Rbb_90_8 bitb_90_8 bitb_90_9 R_bl
Cb_90_8 bit_90_8 gnd C_bl
Cbb_90_8 bitb_90_8 gnd C_bl
Rb_90_9 bit_90_9 bit_90_10 R_bl
Rbb_90_9 bitb_90_9 bitb_90_10 R_bl
Cb_90_9 bit_90_9 gnd C_bl
Cbb_90_9 bitb_90_9 gnd C_bl
Rb_90_10 bit_90_10 bit_90_11 R_bl
Rbb_90_10 bitb_90_10 bitb_90_11 R_bl
Cb_90_10 bit_90_10 gnd C_bl
Cbb_90_10 bitb_90_10 gnd C_bl
Rb_90_11 bit_90_11 bit_90_12 R_bl
Rbb_90_11 bitb_90_11 bitb_90_12 R_bl
Cb_90_11 bit_90_11 gnd C_bl
Cbb_90_11 bitb_90_11 gnd C_bl
Rb_90_12 bit_90_12 bit_90_13 R_bl
Rbb_90_12 bitb_90_12 bitb_90_13 R_bl
Cb_90_12 bit_90_12 gnd C_bl
Cbb_90_12 bitb_90_12 gnd C_bl
Rb_90_13 bit_90_13 bit_90_14 R_bl
Rbb_90_13 bitb_90_13 bitb_90_14 R_bl
Cb_90_13 bit_90_13 gnd C_bl
Cbb_90_13 bitb_90_13 gnd C_bl
Rb_90_14 bit_90_14 bit_90_15 R_bl
Rbb_90_14 bitb_90_14 bitb_90_15 R_bl
Cb_90_14 bit_90_14 gnd C_bl
Cbb_90_14 bitb_90_14 gnd C_bl
Rb_90_15 bit_90_15 bit_90_16 R_bl
Rbb_90_15 bitb_90_15 bitb_90_16 R_bl
Cb_90_15 bit_90_15 gnd C_bl
Cbb_90_15 bitb_90_15 gnd C_bl
Rb_90_16 bit_90_16 bit_90_17 R_bl
Rbb_90_16 bitb_90_16 bitb_90_17 R_bl
Cb_90_16 bit_90_16 gnd C_bl
Cbb_90_16 bitb_90_16 gnd C_bl
Rb_90_17 bit_90_17 bit_90_18 R_bl
Rbb_90_17 bitb_90_17 bitb_90_18 R_bl
Cb_90_17 bit_90_17 gnd C_bl
Cbb_90_17 bitb_90_17 gnd C_bl
Rb_90_18 bit_90_18 bit_90_19 R_bl
Rbb_90_18 bitb_90_18 bitb_90_19 R_bl
Cb_90_18 bit_90_18 gnd C_bl
Cbb_90_18 bitb_90_18 gnd C_bl
Rb_90_19 bit_90_19 bit_90_20 R_bl
Rbb_90_19 bitb_90_19 bitb_90_20 R_bl
Cb_90_19 bit_90_19 gnd C_bl
Cbb_90_19 bitb_90_19 gnd C_bl
Rb_90_20 bit_90_20 bit_90_21 R_bl
Rbb_90_20 bitb_90_20 bitb_90_21 R_bl
Cb_90_20 bit_90_20 gnd C_bl
Cbb_90_20 bitb_90_20 gnd C_bl
Rb_90_21 bit_90_21 bit_90_22 R_bl
Rbb_90_21 bitb_90_21 bitb_90_22 R_bl
Cb_90_21 bit_90_21 gnd C_bl
Cbb_90_21 bitb_90_21 gnd C_bl
Rb_90_22 bit_90_22 bit_90_23 R_bl
Rbb_90_22 bitb_90_22 bitb_90_23 R_bl
Cb_90_22 bit_90_22 gnd C_bl
Cbb_90_22 bitb_90_22 gnd C_bl
Rb_90_23 bit_90_23 bit_90_24 R_bl
Rbb_90_23 bitb_90_23 bitb_90_24 R_bl
Cb_90_23 bit_90_23 gnd C_bl
Cbb_90_23 bitb_90_23 gnd C_bl
Rb_90_24 bit_90_24 bit_90_25 R_bl
Rbb_90_24 bitb_90_24 bitb_90_25 R_bl
Cb_90_24 bit_90_24 gnd C_bl
Cbb_90_24 bitb_90_24 gnd C_bl
Rb_90_25 bit_90_25 bit_90_26 R_bl
Rbb_90_25 bitb_90_25 bitb_90_26 R_bl
Cb_90_25 bit_90_25 gnd C_bl
Cbb_90_25 bitb_90_25 gnd C_bl
Rb_90_26 bit_90_26 bit_90_27 R_bl
Rbb_90_26 bitb_90_26 bitb_90_27 R_bl
Cb_90_26 bit_90_26 gnd C_bl
Cbb_90_26 bitb_90_26 gnd C_bl
Rb_90_27 bit_90_27 bit_90_28 R_bl
Rbb_90_27 bitb_90_27 bitb_90_28 R_bl
Cb_90_27 bit_90_27 gnd C_bl
Cbb_90_27 bitb_90_27 gnd C_bl
Rb_90_28 bit_90_28 bit_90_29 R_bl
Rbb_90_28 bitb_90_28 bitb_90_29 R_bl
Cb_90_28 bit_90_28 gnd C_bl
Cbb_90_28 bitb_90_28 gnd C_bl
Rb_90_29 bit_90_29 bit_90_30 R_bl
Rbb_90_29 bitb_90_29 bitb_90_30 R_bl
Cb_90_29 bit_90_29 gnd C_bl
Cbb_90_29 bitb_90_29 gnd C_bl
Rb_90_30 bit_90_30 bit_90_31 R_bl
Rbb_90_30 bitb_90_30 bitb_90_31 R_bl
Cb_90_30 bit_90_30 gnd C_bl
Cbb_90_30 bitb_90_30 gnd C_bl
Rb_90_31 bit_90_31 bit_90_32 R_bl
Rbb_90_31 bitb_90_31 bitb_90_32 R_bl
Cb_90_31 bit_90_31 gnd C_bl
Cbb_90_31 bitb_90_31 gnd C_bl
Rb_90_32 bit_90_32 bit_90_33 R_bl
Rbb_90_32 bitb_90_32 bitb_90_33 R_bl
Cb_90_32 bit_90_32 gnd C_bl
Cbb_90_32 bitb_90_32 gnd C_bl
Rb_90_33 bit_90_33 bit_90_34 R_bl
Rbb_90_33 bitb_90_33 bitb_90_34 R_bl
Cb_90_33 bit_90_33 gnd C_bl
Cbb_90_33 bitb_90_33 gnd C_bl
Rb_90_34 bit_90_34 bit_90_35 R_bl
Rbb_90_34 bitb_90_34 bitb_90_35 R_bl
Cb_90_34 bit_90_34 gnd C_bl
Cbb_90_34 bitb_90_34 gnd C_bl
Rb_90_35 bit_90_35 bit_90_36 R_bl
Rbb_90_35 bitb_90_35 bitb_90_36 R_bl
Cb_90_35 bit_90_35 gnd C_bl
Cbb_90_35 bitb_90_35 gnd C_bl
Rb_90_36 bit_90_36 bit_90_37 R_bl
Rbb_90_36 bitb_90_36 bitb_90_37 R_bl
Cb_90_36 bit_90_36 gnd C_bl
Cbb_90_36 bitb_90_36 gnd C_bl
Rb_90_37 bit_90_37 bit_90_38 R_bl
Rbb_90_37 bitb_90_37 bitb_90_38 R_bl
Cb_90_37 bit_90_37 gnd C_bl
Cbb_90_37 bitb_90_37 gnd C_bl
Rb_90_38 bit_90_38 bit_90_39 R_bl
Rbb_90_38 bitb_90_38 bitb_90_39 R_bl
Cb_90_38 bit_90_38 gnd C_bl
Cbb_90_38 bitb_90_38 gnd C_bl
Rb_90_39 bit_90_39 bit_90_40 R_bl
Rbb_90_39 bitb_90_39 bitb_90_40 R_bl
Cb_90_39 bit_90_39 gnd C_bl
Cbb_90_39 bitb_90_39 gnd C_bl
Rb_90_40 bit_90_40 bit_90_41 R_bl
Rbb_90_40 bitb_90_40 bitb_90_41 R_bl
Cb_90_40 bit_90_40 gnd C_bl
Cbb_90_40 bitb_90_40 gnd C_bl
Rb_90_41 bit_90_41 bit_90_42 R_bl
Rbb_90_41 bitb_90_41 bitb_90_42 R_bl
Cb_90_41 bit_90_41 gnd C_bl
Cbb_90_41 bitb_90_41 gnd C_bl
Rb_90_42 bit_90_42 bit_90_43 R_bl
Rbb_90_42 bitb_90_42 bitb_90_43 R_bl
Cb_90_42 bit_90_42 gnd C_bl
Cbb_90_42 bitb_90_42 gnd C_bl
Rb_90_43 bit_90_43 bit_90_44 R_bl
Rbb_90_43 bitb_90_43 bitb_90_44 R_bl
Cb_90_43 bit_90_43 gnd C_bl
Cbb_90_43 bitb_90_43 gnd C_bl
Rb_90_44 bit_90_44 bit_90_45 R_bl
Rbb_90_44 bitb_90_44 bitb_90_45 R_bl
Cb_90_44 bit_90_44 gnd C_bl
Cbb_90_44 bitb_90_44 gnd C_bl
Rb_90_45 bit_90_45 bit_90_46 R_bl
Rbb_90_45 bitb_90_45 bitb_90_46 R_bl
Cb_90_45 bit_90_45 gnd C_bl
Cbb_90_45 bitb_90_45 gnd C_bl
Rb_90_46 bit_90_46 bit_90_47 R_bl
Rbb_90_46 bitb_90_46 bitb_90_47 R_bl
Cb_90_46 bit_90_46 gnd C_bl
Cbb_90_46 bitb_90_46 gnd C_bl
Rb_90_47 bit_90_47 bit_90_48 R_bl
Rbb_90_47 bitb_90_47 bitb_90_48 R_bl
Cb_90_47 bit_90_47 gnd C_bl
Cbb_90_47 bitb_90_47 gnd C_bl
Rb_90_48 bit_90_48 bit_90_49 R_bl
Rbb_90_48 bitb_90_48 bitb_90_49 R_bl
Cb_90_48 bit_90_48 gnd C_bl
Cbb_90_48 bitb_90_48 gnd C_bl
Rb_90_49 bit_90_49 bit_90_50 R_bl
Rbb_90_49 bitb_90_49 bitb_90_50 R_bl
Cb_90_49 bit_90_49 gnd C_bl
Cbb_90_49 bitb_90_49 gnd C_bl
Rb_90_50 bit_90_50 bit_90_51 R_bl
Rbb_90_50 bitb_90_50 bitb_90_51 R_bl
Cb_90_50 bit_90_50 gnd C_bl
Cbb_90_50 bitb_90_50 gnd C_bl
Rb_90_51 bit_90_51 bit_90_52 R_bl
Rbb_90_51 bitb_90_51 bitb_90_52 R_bl
Cb_90_51 bit_90_51 gnd C_bl
Cbb_90_51 bitb_90_51 gnd C_bl
Rb_90_52 bit_90_52 bit_90_53 R_bl
Rbb_90_52 bitb_90_52 bitb_90_53 R_bl
Cb_90_52 bit_90_52 gnd C_bl
Cbb_90_52 bitb_90_52 gnd C_bl
Rb_90_53 bit_90_53 bit_90_54 R_bl
Rbb_90_53 bitb_90_53 bitb_90_54 R_bl
Cb_90_53 bit_90_53 gnd C_bl
Cbb_90_53 bitb_90_53 gnd C_bl
Rb_90_54 bit_90_54 bit_90_55 R_bl
Rbb_90_54 bitb_90_54 bitb_90_55 R_bl
Cb_90_54 bit_90_54 gnd C_bl
Cbb_90_54 bitb_90_54 gnd C_bl
Rb_90_55 bit_90_55 bit_90_56 R_bl
Rbb_90_55 bitb_90_55 bitb_90_56 R_bl
Cb_90_55 bit_90_55 gnd C_bl
Cbb_90_55 bitb_90_55 gnd C_bl
Rb_90_56 bit_90_56 bit_90_57 R_bl
Rbb_90_56 bitb_90_56 bitb_90_57 R_bl
Cb_90_56 bit_90_56 gnd C_bl
Cbb_90_56 bitb_90_56 gnd C_bl
Rb_90_57 bit_90_57 bit_90_58 R_bl
Rbb_90_57 bitb_90_57 bitb_90_58 R_bl
Cb_90_57 bit_90_57 gnd C_bl
Cbb_90_57 bitb_90_57 gnd C_bl
Rb_90_58 bit_90_58 bit_90_59 R_bl
Rbb_90_58 bitb_90_58 bitb_90_59 R_bl
Cb_90_58 bit_90_58 gnd C_bl
Cbb_90_58 bitb_90_58 gnd C_bl
Rb_90_59 bit_90_59 bit_90_60 R_bl
Rbb_90_59 bitb_90_59 bitb_90_60 R_bl
Cb_90_59 bit_90_59 gnd C_bl
Cbb_90_59 bitb_90_59 gnd C_bl
Rb_90_60 bit_90_60 bit_90_61 R_bl
Rbb_90_60 bitb_90_60 bitb_90_61 R_bl
Cb_90_60 bit_90_60 gnd C_bl
Cbb_90_60 bitb_90_60 gnd C_bl
Rb_90_61 bit_90_61 bit_90_62 R_bl
Rbb_90_61 bitb_90_61 bitb_90_62 R_bl
Cb_90_61 bit_90_61 gnd C_bl
Cbb_90_61 bitb_90_61 gnd C_bl
Rb_90_62 bit_90_62 bit_90_63 R_bl
Rbb_90_62 bitb_90_62 bitb_90_63 R_bl
Cb_90_62 bit_90_62 gnd C_bl
Cbb_90_62 bitb_90_62 gnd C_bl
Rb_90_63 bit_90_63 bit_90_64 R_bl
Rbb_90_63 bitb_90_63 bitb_90_64 R_bl
Cb_90_63 bit_90_63 gnd C_bl
Cbb_90_63 bitb_90_63 gnd C_bl
Rb_90_64 bit_90_64 bit_90_65 R_bl
Rbb_90_64 bitb_90_64 bitb_90_65 R_bl
Cb_90_64 bit_90_64 gnd C_bl
Cbb_90_64 bitb_90_64 gnd C_bl
Rb_90_65 bit_90_65 bit_90_66 R_bl
Rbb_90_65 bitb_90_65 bitb_90_66 R_bl
Cb_90_65 bit_90_65 gnd C_bl
Cbb_90_65 bitb_90_65 gnd C_bl
Rb_90_66 bit_90_66 bit_90_67 R_bl
Rbb_90_66 bitb_90_66 bitb_90_67 R_bl
Cb_90_66 bit_90_66 gnd C_bl
Cbb_90_66 bitb_90_66 gnd C_bl
Rb_90_67 bit_90_67 bit_90_68 R_bl
Rbb_90_67 bitb_90_67 bitb_90_68 R_bl
Cb_90_67 bit_90_67 gnd C_bl
Cbb_90_67 bitb_90_67 gnd C_bl
Rb_90_68 bit_90_68 bit_90_69 R_bl
Rbb_90_68 bitb_90_68 bitb_90_69 R_bl
Cb_90_68 bit_90_68 gnd C_bl
Cbb_90_68 bitb_90_68 gnd C_bl
Rb_90_69 bit_90_69 bit_90_70 R_bl
Rbb_90_69 bitb_90_69 bitb_90_70 R_bl
Cb_90_69 bit_90_69 gnd C_bl
Cbb_90_69 bitb_90_69 gnd C_bl
Rb_90_70 bit_90_70 bit_90_71 R_bl
Rbb_90_70 bitb_90_70 bitb_90_71 R_bl
Cb_90_70 bit_90_70 gnd C_bl
Cbb_90_70 bitb_90_70 gnd C_bl
Rb_90_71 bit_90_71 bit_90_72 R_bl
Rbb_90_71 bitb_90_71 bitb_90_72 R_bl
Cb_90_71 bit_90_71 gnd C_bl
Cbb_90_71 bitb_90_71 gnd C_bl
Rb_90_72 bit_90_72 bit_90_73 R_bl
Rbb_90_72 bitb_90_72 bitb_90_73 R_bl
Cb_90_72 bit_90_72 gnd C_bl
Cbb_90_72 bitb_90_72 gnd C_bl
Rb_90_73 bit_90_73 bit_90_74 R_bl
Rbb_90_73 bitb_90_73 bitb_90_74 R_bl
Cb_90_73 bit_90_73 gnd C_bl
Cbb_90_73 bitb_90_73 gnd C_bl
Rb_90_74 bit_90_74 bit_90_75 R_bl
Rbb_90_74 bitb_90_74 bitb_90_75 R_bl
Cb_90_74 bit_90_74 gnd C_bl
Cbb_90_74 bitb_90_74 gnd C_bl
Rb_90_75 bit_90_75 bit_90_76 R_bl
Rbb_90_75 bitb_90_75 bitb_90_76 R_bl
Cb_90_75 bit_90_75 gnd C_bl
Cbb_90_75 bitb_90_75 gnd C_bl
Rb_90_76 bit_90_76 bit_90_77 R_bl
Rbb_90_76 bitb_90_76 bitb_90_77 R_bl
Cb_90_76 bit_90_76 gnd C_bl
Cbb_90_76 bitb_90_76 gnd C_bl
Rb_90_77 bit_90_77 bit_90_78 R_bl
Rbb_90_77 bitb_90_77 bitb_90_78 R_bl
Cb_90_77 bit_90_77 gnd C_bl
Cbb_90_77 bitb_90_77 gnd C_bl
Rb_90_78 bit_90_78 bit_90_79 R_bl
Rbb_90_78 bitb_90_78 bitb_90_79 R_bl
Cb_90_78 bit_90_78 gnd C_bl
Cbb_90_78 bitb_90_78 gnd C_bl
Rb_90_79 bit_90_79 bit_90_80 R_bl
Rbb_90_79 bitb_90_79 bitb_90_80 R_bl
Cb_90_79 bit_90_79 gnd C_bl
Cbb_90_79 bitb_90_79 gnd C_bl
Rb_90_80 bit_90_80 bit_90_81 R_bl
Rbb_90_80 bitb_90_80 bitb_90_81 R_bl
Cb_90_80 bit_90_80 gnd C_bl
Cbb_90_80 bitb_90_80 gnd C_bl
Rb_90_81 bit_90_81 bit_90_82 R_bl
Rbb_90_81 bitb_90_81 bitb_90_82 R_bl
Cb_90_81 bit_90_81 gnd C_bl
Cbb_90_81 bitb_90_81 gnd C_bl
Rb_90_82 bit_90_82 bit_90_83 R_bl
Rbb_90_82 bitb_90_82 bitb_90_83 R_bl
Cb_90_82 bit_90_82 gnd C_bl
Cbb_90_82 bitb_90_82 gnd C_bl
Rb_90_83 bit_90_83 bit_90_84 R_bl
Rbb_90_83 bitb_90_83 bitb_90_84 R_bl
Cb_90_83 bit_90_83 gnd C_bl
Cbb_90_83 bitb_90_83 gnd C_bl
Rb_90_84 bit_90_84 bit_90_85 R_bl
Rbb_90_84 bitb_90_84 bitb_90_85 R_bl
Cb_90_84 bit_90_84 gnd C_bl
Cbb_90_84 bitb_90_84 gnd C_bl
Rb_90_85 bit_90_85 bit_90_86 R_bl
Rbb_90_85 bitb_90_85 bitb_90_86 R_bl
Cb_90_85 bit_90_85 gnd C_bl
Cbb_90_85 bitb_90_85 gnd C_bl
Rb_90_86 bit_90_86 bit_90_87 R_bl
Rbb_90_86 bitb_90_86 bitb_90_87 R_bl
Cb_90_86 bit_90_86 gnd C_bl
Cbb_90_86 bitb_90_86 gnd C_bl
Rb_90_87 bit_90_87 bit_90_88 R_bl
Rbb_90_87 bitb_90_87 bitb_90_88 R_bl
Cb_90_87 bit_90_87 gnd C_bl
Cbb_90_87 bitb_90_87 gnd C_bl
Rb_90_88 bit_90_88 bit_90_89 R_bl
Rbb_90_88 bitb_90_88 bitb_90_89 R_bl
Cb_90_88 bit_90_88 gnd C_bl
Cbb_90_88 bitb_90_88 gnd C_bl
Rb_90_89 bit_90_89 bit_90_90 R_bl
Rbb_90_89 bitb_90_89 bitb_90_90 R_bl
Cb_90_89 bit_90_89 gnd C_bl
Cbb_90_89 bitb_90_89 gnd C_bl
Rb_90_90 bit_90_90 bit_90_91 R_bl
Rbb_90_90 bitb_90_90 bitb_90_91 R_bl
Cb_90_90 bit_90_90 gnd C_bl
Cbb_90_90 bitb_90_90 gnd C_bl
Rb_90_91 bit_90_91 bit_90_92 R_bl
Rbb_90_91 bitb_90_91 bitb_90_92 R_bl
Cb_90_91 bit_90_91 gnd C_bl
Cbb_90_91 bitb_90_91 gnd C_bl
Rb_90_92 bit_90_92 bit_90_93 R_bl
Rbb_90_92 bitb_90_92 bitb_90_93 R_bl
Cb_90_92 bit_90_92 gnd C_bl
Cbb_90_92 bitb_90_92 gnd C_bl
Rb_90_93 bit_90_93 bit_90_94 R_bl
Rbb_90_93 bitb_90_93 bitb_90_94 R_bl
Cb_90_93 bit_90_93 gnd C_bl
Cbb_90_93 bitb_90_93 gnd C_bl
Rb_90_94 bit_90_94 bit_90_95 R_bl
Rbb_90_94 bitb_90_94 bitb_90_95 R_bl
Cb_90_94 bit_90_94 gnd C_bl
Cbb_90_94 bitb_90_94 gnd C_bl
Rb_90_95 bit_90_95 bit_90_96 R_bl
Rbb_90_95 bitb_90_95 bitb_90_96 R_bl
Cb_90_95 bit_90_95 gnd C_bl
Cbb_90_95 bitb_90_95 gnd C_bl
Rb_90_96 bit_90_96 bit_90_97 R_bl
Rbb_90_96 bitb_90_96 bitb_90_97 R_bl
Cb_90_96 bit_90_96 gnd C_bl
Cbb_90_96 bitb_90_96 gnd C_bl
Rb_90_97 bit_90_97 bit_90_98 R_bl
Rbb_90_97 bitb_90_97 bitb_90_98 R_bl
Cb_90_97 bit_90_97 gnd C_bl
Cbb_90_97 bitb_90_97 gnd C_bl
Rb_90_98 bit_90_98 bit_90_99 R_bl
Rbb_90_98 bitb_90_98 bitb_90_99 R_bl
Cb_90_98 bit_90_98 gnd C_bl
Cbb_90_98 bitb_90_98 gnd C_bl
Rb_90_99 bit_90_99 bit_90_100 R_bl
Rbb_90_99 bitb_90_99 bitb_90_100 R_bl
Cb_90_99 bit_90_99 gnd C_bl
Cbb_90_99 bitb_90_99 gnd C_bl
Rb_91_0 bit_91_0 bit_91_1 R_bl
Rbb_91_0 bitb_91_0 bitb_91_1 R_bl
Cb_91_0 bit_91_0 gnd C_bl
Cbb_91_0 bitb_91_0 gnd C_bl
Rb_91_1 bit_91_1 bit_91_2 R_bl
Rbb_91_1 bitb_91_1 bitb_91_2 R_bl
Cb_91_1 bit_91_1 gnd C_bl
Cbb_91_1 bitb_91_1 gnd C_bl
Rb_91_2 bit_91_2 bit_91_3 R_bl
Rbb_91_2 bitb_91_2 bitb_91_3 R_bl
Cb_91_2 bit_91_2 gnd C_bl
Cbb_91_2 bitb_91_2 gnd C_bl
Rb_91_3 bit_91_3 bit_91_4 R_bl
Rbb_91_3 bitb_91_3 bitb_91_4 R_bl
Cb_91_3 bit_91_3 gnd C_bl
Cbb_91_3 bitb_91_3 gnd C_bl
Rb_91_4 bit_91_4 bit_91_5 R_bl
Rbb_91_4 bitb_91_4 bitb_91_5 R_bl
Cb_91_4 bit_91_4 gnd C_bl
Cbb_91_4 bitb_91_4 gnd C_bl
Rb_91_5 bit_91_5 bit_91_6 R_bl
Rbb_91_5 bitb_91_5 bitb_91_6 R_bl
Cb_91_5 bit_91_5 gnd C_bl
Cbb_91_5 bitb_91_5 gnd C_bl
Rb_91_6 bit_91_6 bit_91_7 R_bl
Rbb_91_6 bitb_91_6 bitb_91_7 R_bl
Cb_91_6 bit_91_6 gnd C_bl
Cbb_91_6 bitb_91_6 gnd C_bl
Rb_91_7 bit_91_7 bit_91_8 R_bl
Rbb_91_7 bitb_91_7 bitb_91_8 R_bl
Cb_91_7 bit_91_7 gnd C_bl
Cbb_91_7 bitb_91_7 gnd C_bl
Rb_91_8 bit_91_8 bit_91_9 R_bl
Rbb_91_8 bitb_91_8 bitb_91_9 R_bl
Cb_91_8 bit_91_8 gnd C_bl
Cbb_91_8 bitb_91_8 gnd C_bl
Rb_91_9 bit_91_9 bit_91_10 R_bl
Rbb_91_9 bitb_91_9 bitb_91_10 R_bl
Cb_91_9 bit_91_9 gnd C_bl
Cbb_91_9 bitb_91_9 gnd C_bl
Rb_91_10 bit_91_10 bit_91_11 R_bl
Rbb_91_10 bitb_91_10 bitb_91_11 R_bl
Cb_91_10 bit_91_10 gnd C_bl
Cbb_91_10 bitb_91_10 gnd C_bl
Rb_91_11 bit_91_11 bit_91_12 R_bl
Rbb_91_11 bitb_91_11 bitb_91_12 R_bl
Cb_91_11 bit_91_11 gnd C_bl
Cbb_91_11 bitb_91_11 gnd C_bl
Rb_91_12 bit_91_12 bit_91_13 R_bl
Rbb_91_12 bitb_91_12 bitb_91_13 R_bl
Cb_91_12 bit_91_12 gnd C_bl
Cbb_91_12 bitb_91_12 gnd C_bl
Rb_91_13 bit_91_13 bit_91_14 R_bl
Rbb_91_13 bitb_91_13 bitb_91_14 R_bl
Cb_91_13 bit_91_13 gnd C_bl
Cbb_91_13 bitb_91_13 gnd C_bl
Rb_91_14 bit_91_14 bit_91_15 R_bl
Rbb_91_14 bitb_91_14 bitb_91_15 R_bl
Cb_91_14 bit_91_14 gnd C_bl
Cbb_91_14 bitb_91_14 gnd C_bl
Rb_91_15 bit_91_15 bit_91_16 R_bl
Rbb_91_15 bitb_91_15 bitb_91_16 R_bl
Cb_91_15 bit_91_15 gnd C_bl
Cbb_91_15 bitb_91_15 gnd C_bl
Rb_91_16 bit_91_16 bit_91_17 R_bl
Rbb_91_16 bitb_91_16 bitb_91_17 R_bl
Cb_91_16 bit_91_16 gnd C_bl
Cbb_91_16 bitb_91_16 gnd C_bl
Rb_91_17 bit_91_17 bit_91_18 R_bl
Rbb_91_17 bitb_91_17 bitb_91_18 R_bl
Cb_91_17 bit_91_17 gnd C_bl
Cbb_91_17 bitb_91_17 gnd C_bl
Rb_91_18 bit_91_18 bit_91_19 R_bl
Rbb_91_18 bitb_91_18 bitb_91_19 R_bl
Cb_91_18 bit_91_18 gnd C_bl
Cbb_91_18 bitb_91_18 gnd C_bl
Rb_91_19 bit_91_19 bit_91_20 R_bl
Rbb_91_19 bitb_91_19 bitb_91_20 R_bl
Cb_91_19 bit_91_19 gnd C_bl
Cbb_91_19 bitb_91_19 gnd C_bl
Rb_91_20 bit_91_20 bit_91_21 R_bl
Rbb_91_20 bitb_91_20 bitb_91_21 R_bl
Cb_91_20 bit_91_20 gnd C_bl
Cbb_91_20 bitb_91_20 gnd C_bl
Rb_91_21 bit_91_21 bit_91_22 R_bl
Rbb_91_21 bitb_91_21 bitb_91_22 R_bl
Cb_91_21 bit_91_21 gnd C_bl
Cbb_91_21 bitb_91_21 gnd C_bl
Rb_91_22 bit_91_22 bit_91_23 R_bl
Rbb_91_22 bitb_91_22 bitb_91_23 R_bl
Cb_91_22 bit_91_22 gnd C_bl
Cbb_91_22 bitb_91_22 gnd C_bl
Rb_91_23 bit_91_23 bit_91_24 R_bl
Rbb_91_23 bitb_91_23 bitb_91_24 R_bl
Cb_91_23 bit_91_23 gnd C_bl
Cbb_91_23 bitb_91_23 gnd C_bl
Rb_91_24 bit_91_24 bit_91_25 R_bl
Rbb_91_24 bitb_91_24 bitb_91_25 R_bl
Cb_91_24 bit_91_24 gnd C_bl
Cbb_91_24 bitb_91_24 gnd C_bl
Rb_91_25 bit_91_25 bit_91_26 R_bl
Rbb_91_25 bitb_91_25 bitb_91_26 R_bl
Cb_91_25 bit_91_25 gnd C_bl
Cbb_91_25 bitb_91_25 gnd C_bl
Rb_91_26 bit_91_26 bit_91_27 R_bl
Rbb_91_26 bitb_91_26 bitb_91_27 R_bl
Cb_91_26 bit_91_26 gnd C_bl
Cbb_91_26 bitb_91_26 gnd C_bl
Rb_91_27 bit_91_27 bit_91_28 R_bl
Rbb_91_27 bitb_91_27 bitb_91_28 R_bl
Cb_91_27 bit_91_27 gnd C_bl
Cbb_91_27 bitb_91_27 gnd C_bl
Rb_91_28 bit_91_28 bit_91_29 R_bl
Rbb_91_28 bitb_91_28 bitb_91_29 R_bl
Cb_91_28 bit_91_28 gnd C_bl
Cbb_91_28 bitb_91_28 gnd C_bl
Rb_91_29 bit_91_29 bit_91_30 R_bl
Rbb_91_29 bitb_91_29 bitb_91_30 R_bl
Cb_91_29 bit_91_29 gnd C_bl
Cbb_91_29 bitb_91_29 gnd C_bl
Rb_91_30 bit_91_30 bit_91_31 R_bl
Rbb_91_30 bitb_91_30 bitb_91_31 R_bl
Cb_91_30 bit_91_30 gnd C_bl
Cbb_91_30 bitb_91_30 gnd C_bl
Rb_91_31 bit_91_31 bit_91_32 R_bl
Rbb_91_31 bitb_91_31 bitb_91_32 R_bl
Cb_91_31 bit_91_31 gnd C_bl
Cbb_91_31 bitb_91_31 gnd C_bl
Rb_91_32 bit_91_32 bit_91_33 R_bl
Rbb_91_32 bitb_91_32 bitb_91_33 R_bl
Cb_91_32 bit_91_32 gnd C_bl
Cbb_91_32 bitb_91_32 gnd C_bl
Rb_91_33 bit_91_33 bit_91_34 R_bl
Rbb_91_33 bitb_91_33 bitb_91_34 R_bl
Cb_91_33 bit_91_33 gnd C_bl
Cbb_91_33 bitb_91_33 gnd C_bl
Rb_91_34 bit_91_34 bit_91_35 R_bl
Rbb_91_34 bitb_91_34 bitb_91_35 R_bl
Cb_91_34 bit_91_34 gnd C_bl
Cbb_91_34 bitb_91_34 gnd C_bl
Rb_91_35 bit_91_35 bit_91_36 R_bl
Rbb_91_35 bitb_91_35 bitb_91_36 R_bl
Cb_91_35 bit_91_35 gnd C_bl
Cbb_91_35 bitb_91_35 gnd C_bl
Rb_91_36 bit_91_36 bit_91_37 R_bl
Rbb_91_36 bitb_91_36 bitb_91_37 R_bl
Cb_91_36 bit_91_36 gnd C_bl
Cbb_91_36 bitb_91_36 gnd C_bl
Rb_91_37 bit_91_37 bit_91_38 R_bl
Rbb_91_37 bitb_91_37 bitb_91_38 R_bl
Cb_91_37 bit_91_37 gnd C_bl
Cbb_91_37 bitb_91_37 gnd C_bl
Rb_91_38 bit_91_38 bit_91_39 R_bl
Rbb_91_38 bitb_91_38 bitb_91_39 R_bl
Cb_91_38 bit_91_38 gnd C_bl
Cbb_91_38 bitb_91_38 gnd C_bl
Rb_91_39 bit_91_39 bit_91_40 R_bl
Rbb_91_39 bitb_91_39 bitb_91_40 R_bl
Cb_91_39 bit_91_39 gnd C_bl
Cbb_91_39 bitb_91_39 gnd C_bl
Rb_91_40 bit_91_40 bit_91_41 R_bl
Rbb_91_40 bitb_91_40 bitb_91_41 R_bl
Cb_91_40 bit_91_40 gnd C_bl
Cbb_91_40 bitb_91_40 gnd C_bl
Rb_91_41 bit_91_41 bit_91_42 R_bl
Rbb_91_41 bitb_91_41 bitb_91_42 R_bl
Cb_91_41 bit_91_41 gnd C_bl
Cbb_91_41 bitb_91_41 gnd C_bl
Rb_91_42 bit_91_42 bit_91_43 R_bl
Rbb_91_42 bitb_91_42 bitb_91_43 R_bl
Cb_91_42 bit_91_42 gnd C_bl
Cbb_91_42 bitb_91_42 gnd C_bl
Rb_91_43 bit_91_43 bit_91_44 R_bl
Rbb_91_43 bitb_91_43 bitb_91_44 R_bl
Cb_91_43 bit_91_43 gnd C_bl
Cbb_91_43 bitb_91_43 gnd C_bl
Rb_91_44 bit_91_44 bit_91_45 R_bl
Rbb_91_44 bitb_91_44 bitb_91_45 R_bl
Cb_91_44 bit_91_44 gnd C_bl
Cbb_91_44 bitb_91_44 gnd C_bl
Rb_91_45 bit_91_45 bit_91_46 R_bl
Rbb_91_45 bitb_91_45 bitb_91_46 R_bl
Cb_91_45 bit_91_45 gnd C_bl
Cbb_91_45 bitb_91_45 gnd C_bl
Rb_91_46 bit_91_46 bit_91_47 R_bl
Rbb_91_46 bitb_91_46 bitb_91_47 R_bl
Cb_91_46 bit_91_46 gnd C_bl
Cbb_91_46 bitb_91_46 gnd C_bl
Rb_91_47 bit_91_47 bit_91_48 R_bl
Rbb_91_47 bitb_91_47 bitb_91_48 R_bl
Cb_91_47 bit_91_47 gnd C_bl
Cbb_91_47 bitb_91_47 gnd C_bl
Rb_91_48 bit_91_48 bit_91_49 R_bl
Rbb_91_48 bitb_91_48 bitb_91_49 R_bl
Cb_91_48 bit_91_48 gnd C_bl
Cbb_91_48 bitb_91_48 gnd C_bl
Rb_91_49 bit_91_49 bit_91_50 R_bl
Rbb_91_49 bitb_91_49 bitb_91_50 R_bl
Cb_91_49 bit_91_49 gnd C_bl
Cbb_91_49 bitb_91_49 gnd C_bl
Rb_91_50 bit_91_50 bit_91_51 R_bl
Rbb_91_50 bitb_91_50 bitb_91_51 R_bl
Cb_91_50 bit_91_50 gnd C_bl
Cbb_91_50 bitb_91_50 gnd C_bl
Rb_91_51 bit_91_51 bit_91_52 R_bl
Rbb_91_51 bitb_91_51 bitb_91_52 R_bl
Cb_91_51 bit_91_51 gnd C_bl
Cbb_91_51 bitb_91_51 gnd C_bl
Rb_91_52 bit_91_52 bit_91_53 R_bl
Rbb_91_52 bitb_91_52 bitb_91_53 R_bl
Cb_91_52 bit_91_52 gnd C_bl
Cbb_91_52 bitb_91_52 gnd C_bl
Rb_91_53 bit_91_53 bit_91_54 R_bl
Rbb_91_53 bitb_91_53 bitb_91_54 R_bl
Cb_91_53 bit_91_53 gnd C_bl
Cbb_91_53 bitb_91_53 gnd C_bl
Rb_91_54 bit_91_54 bit_91_55 R_bl
Rbb_91_54 bitb_91_54 bitb_91_55 R_bl
Cb_91_54 bit_91_54 gnd C_bl
Cbb_91_54 bitb_91_54 gnd C_bl
Rb_91_55 bit_91_55 bit_91_56 R_bl
Rbb_91_55 bitb_91_55 bitb_91_56 R_bl
Cb_91_55 bit_91_55 gnd C_bl
Cbb_91_55 bitb_91_55 gnd C_bl
Rb_91_56 bit_91_56 bit_91_57 R_bl
Rbb_91_56 bitb_91_56 bitb_91_57 R_bl
Cb_91_56 bit_91_56 gnd C_bl
Cbb_91_56 bitb_91_56 gnd C_bl
Rb_91_57 bit_91_57 bit_91_58 R_bl
Rbb_91_57 bitb_91_57 bitb_91_58 R_bl
Cb_91_57 bit_91_57 gnd C_bl
Cbb_91_57 bitb_91_57 gnd C_bl
Rb_91_58 bit_91_58 bit_91_59 R_bl
Rbb_91_58 bitb_91_58 bitb_91_59 R_bl
Cb_91_58 bit_91_58 gnd C_bl
Cbb_91_58 bitb_91_58 gnd C_bl
Rb_91_59 bit_91_59 bit_91_60 R_bl
Rbb_91_59 bitb_91_59 bitb_91_60 R_bl
Cb_91_59 bit_91_59 gnd C_bl
Cbb_91_59 bitb_91_59 gnd C_bl
Rb_91_60 bit_91_60 bit_91_61 R_bl
Rbb_91_60 bitb_91_60 bitb_91_61 R_bl
Cb_91_60 bit_91_60 gnd C_bl
Cbb_91_60 bitb_91_60 gnd C_bl
Rb_91_61 bit_91_61 bit_91_62 R_bl
Rbb_91_61 bitb_91_61 bitb_91_62 R_bl
Cb_91_61 bit_91_61 gnd C_bl
Cbb_91_61 bitb_91_61 gnd C_bl
Rb_91_62 bit_91_62 bit_91_63 R_bl
Rbb_91_62 bitb_91_62 bitb_91_63 R_bl
Cb_91_62 bit_91_62 gnd C_bl
Cbb_91_62 bitb_91_62 gnd C_bl
Rb_91_63 bit_91_63 bit_91_64 R_bl
Rbb_91_63 bitb_91_63 bitb_91_64 R_bl
Cb_91_63 bit_91_63 gnd C_bl
Cbb_91_63 bitb_91_63 gnd C_bl
Rb_91_64 bit_91_64 bit_91_65 R_bl
Rbb_91_64 bitb_91_64 bitb_91_65 R_bl
Cb_91_64 bit_91_64 gnd C_bl
Cbb_91_64 bitb_91_64 gnd C_bl
Rb_91_65 bit_91_65 bit_91_66 R_bl
Rbb_91_65 bitb_91_65 bitb_91_66 R_bl
Cb_91_65 bit_91_65 gnd C_bl
Cbb_91_65 bitb_91_65 gnd C_bl
Rb_91_66 bit_91_66 bit_91_67 R_bl
Rbb_91_66 bitb_91_66 bitb_91_67 R_bl
Cb_91_66 bit_91_66 gnd C_bl
Cbb_91_66 bitb_91_66 gnd C_bl
Rb_91_67 bit_91_67 bit_91_68 R_bl
Rbb_91_67 bitb_91_67 bitb_91_68 R_bl
Cb_91_67 bit_91_67 gnd C_bl
Cbb_91_67 bitb_91_67 gnd C_bl
Rb_91_68 bit_91_68 bit_91_69 R_bl
Rbb_91_68 bitb_91_68 bitb_91_69 R_bl
Cb_91_68 bit_91_68 gnd C_bl
Cbb_91_68 bitb_91_68 gnd C_bl
Rb_91_69 bit_91_69 bit_91_70 R_bl
Rbb_91_69 bitb_91_69 bitb_91_70 R_bl
Cb_91_69 bit_91_69 gnd C_bl
Cbb_91_69 bitb_91_69 gnd C_bl
Rb_91_70 bit_91_70 bit_91_71 R_bl
Rbb_91_70 bitb_91_70 bitb_91_71 R_bl
Cb_91_70 bit_91_70 gnd C_bl
Cbb_91_70 bitb_91_70 gnd C_bl
Rb_91_71 bit_91_71 bit_91_72 R_bl
Rbb_91_71 bitb_91_71 bitb_91_72 R_bl
Cb_91_71 bit_91_71 gnd C_bl
Cbb_91_71 bitb_91_71 gnd C_bl
Rb_91_72 bit_91_72 bit_91_73 R_bl
Rbb_91_72 bitb_91_72 bitb_91_73 R_bl
Cb_91_72 bit_91_72 gnd C_bl
Cbb_91_72 bitb_91_72 gnd C_bl
Rb_91_73 bit_91_73 bit_91_74 R_bl
Rbb_91_73 bitb_91_73 bitb_91_74 R_bl
Cb_91_73 bit_91_73 gnd C_bl
Cbb_91_73 bitb_91_73 gnd C_bl
Rb_91_74 bit_91_74 bit_91_75 R_bl
Rbb_91_74 bitb_91_74 bitb_91_75 R_bl
Cb_91_74 bit_91_74 gnd C_bl
Cbb_91_74 bitb_91_74 gnd C_bl
Rb_91_75 bit_91_75 bit_91_76 R_bl
Rbb_91_75 bitb_91_75 bitb_91_76 R_bl
Cb_91_75 bit_91_75 gnd C_bl
Cbb_91_75 bitb_91_75 gnd C_bl
Rb_91_76 bit_91_76 bit_91_77 R_bl
Rbb_91_76 bitb_91_76 bitb_91_77 R_bl
Cb_91_76 bit_91_76 gnd C_bl
Cbb_91_76 bitb_91_76 gnd C_bl
Rb_91_77 bit_91_77 bit_91_78 R_bl
Rbb_91_77 bitb_91_77 bitb_91_78 R_bl
Cb_91_77 bit_91_77 gnd C_bl
Cbb_91_77 bitb_91_77 gnd C_bl
Rb_91_78 bit_91_78 bit_91_79 R_bl
Rbb_91_78 bitb_91_78 bitb_91_79 R_bl
Cb_91_78 bit_91_78 gnd C_bl
Cbb_91_78 bitb_91_78 gnd C_bl
Rb_91_79 bit_91_79 bit_91_80 R_bl
Rbb_91_79 bitb_91_79 bitb_91_80 R_bl
Cb_91_79 bit_91_79 gnd C_bl
Cbb_91_79 bitb_91_79 gnd C_bl
Rb_91_80 bit_91_80 bit_91_81 R_bl
Rbb_91_80 bitb_91_80 bitb_91_81 R_bl
Cb_91_80 bit_91_80 gnd C_bl
Cbb_91_80 bitb_91_80 gnd C_bl
Rb_91_81 bit_91_81 bit_91_82 R_bl
Rbb_91_81 bitb_91_81 bitb_91_82 R_bl
Cb_91_81 bit_91_81 gnd C_bl
Cbb_91_81 bitb_91_81 gnd C_bl
Rb_91_82 bit_91_82 bit_91_83 R_bl
Rbb_91_82 bitb_91_82 bitb_91_83 R_bl
Cb_91_82 bit_91_82 gnd C_bl
Cbb_91_82 bitb_91_82 gnd C_bl
Rb_91_83 bit_91_83 bit_91_84 R_bl
Rbb_91_83 bitb_91_83 bitb_91_84 R_bl
Cb_91_83 bit_91_83 gnd C_bl
Cbb_91_83 bitb_91_83 gnd C_bl
Rb_91_84 bit_91_84 bit_91_85 R_bl
Rbb_91_84 bitb_91_84 bitb_91_85 R_bl
Cb_91_84 bit_91_84 gnd C_bl
Cbb_91_84 bitb_91_84 gnd C_bl
Rb_91_85 bit_91_85 bit_91_86 R_bl
Rbb_91_85 bitb_91_85 bitb_91_86 R_bl
Cb_91_85 bit_91_85 gnd C_bl
Cbb_91_85 bitb_91_85 gnd C_bl
Rb_91_86 bit_91_86 bit_91_87 R_bl
Rbb_91_86 bitb_91_86 bitb_91_87 R_bl
Cb_91_86 bit_91_86 gnd C_bl
Cbb_91_86 bitb_91_86 gnd C_bl
Rb_91_87 bit_91_87 bit_91_88 R_bl
Rbb_91_87 bitb_91_87 bitb_91_88 R_bl
Cb_91_87 bit_91_87 gnd C_bl
Cbb_91_87 bitb_91_87 gnd C_bl
Rb_91_88 bit_91_88 bit_91_89 R_bl
Rbb_91_88 bitb_91_88 bitb_91_89 R_bl
Cb_91_88 bit_91_88 gnd C_bl
Cbb_91_88 bitb_91_88 gnd C_bl
Rb_91_89 bit_91_89 bit_91_90 R_bl
Rbb_91_89 bitb_91_89 bitb_91_90 R_bl
Cb_91_89 bit_91_89 gnd C_bl
Cbb_91_89 bitb_91_89 gnd C_bl
Rb_91_90 bit_91_90 bit_91_91 R_bl
Rbb_91_90 bitb_91_90 bitb_91_91 R_bl
Cb_91_90 bit_91_90 gnd C_bl
Cbb_91_90 bitb_91_90 gnd C_bl
Rb_91_91 bit_91_91 bit_91_92 R_bl
Rbb_91_91 bitb_91_91 bitb_91_92 R_bl
Cb_91_91 bit_91_91 gnd C_bl
Cbb_91_91 bitb_91_91 gnd C_bl
Rb_91_92 bit_91_92 bit_91_93 R_bl
Rbb_91_92 bitb_91_92 bitb_91_93 R_bl
Cb_91_92 bit_91_92 gnd C_bl
Cbb_91_92 bitb_91_92 gnd C_bl
Rb_91_93 bit_91_93 bit_91_94 R_bl
Rbb_91_93 bitb_91_93 bitb_91_94 R_bl
Cb_91_93 bit_91_93 gnd C_bl
Cbb_91_93 bitb_91_93 gnd C_bl
Rb_91_94 bit_91_94 bit_91_95 R_bl
Rbb_91_94 bitb_91_94 bitb_91_95 R_bl
Cb_91_94 bit_91_94 gnd C_bl
Cbb_91_94 bitb_91_94 gnd C_bl
Rb_91_95 bit_91_95 bit_91_96 R_bl
Rbb_91_95 bitb_91_95 bitb_91_96 R_bl
Cb_91_95 bit_91_95 gnd C_bl
Cbb_91_95 bitb_91_95 gnd C_bl
Rb_91_96 bit_91_96 bit_91_97 R_bl
Rbb_91_96 bitb_91_96 bitb_91_97 R_bl
Cb_91_96 bit_91_96 gnd C_bl
Cbb_91_96 bitb_91_96 gnd C_bl
Rb_91_97 bit_91_97 bit_91_98 R_bl
Rbb_91_97 bitb_91_97 bitb_91_98 R_bl
Cb_91_97 bit_91_97 gnd C_bl
Cbb_91_97 bitb_91_97 gnd C_bl
Rb_91_98 bit_91_98 bit_91_99 R_bl
Rbb_91_98 bitb_91_98 bitb_91_99 R_bl
Cb_91_98 bit_91_98 gnd C_bl
Cbb_91_98 bitb_91_98 gnd C_bl
Rb_91_99 bit_91_99 bit_91_100 R_bl
Rbb_91_99 bitb_91_99 bitb_91_100 R_bl
Cb_91_99 bit_91_99 gnd C_bl
Cbb_91_99 bitb_91_99 gnd C_bl
Rb_92_0 bit_92_0 bit_92_1 R_bl
Rbb_92_0 bitb_92_0 bitb_92_1 R_bl
Cb_92_0 bit_92_0 gnd C_bl
Cbb_92_0 bitb_92_0 gnd C_bl
Rb_92_1 bit_92_1 bit_92_2 R_bl
Rbb_92_1 bitb_92_1 bitb_92_2 R_bl
Cb_92_1 bit_92_1 gnd C_bl
Cbb_92_1 bitb_92_1 gnd C_bl
Rb_92_2 bit_92_2 bit_92_3 R_bl
Rbb_92_2 bitb_92_2 bitb_92_3 R_bl
Cb_92_2 bit_92_2 gnd C_bl
Cbb_92_2 bitb_92_2 gnd C_bl
Rb_92_3 bit_92_3 bit_92_4 R_bl
Rbb_92_3 bitb_92_3 bitb_92_4 R_bl
Cb_92_3 bit_92_3 gnd C_bl
Cbb_92_3 bitb_92_3 gnd C_bl
Rb_92_4 bit_92_4 bit_92_5 R_bl
Rbb_92_4 bitb_92_4 bitb_92_5 R_bl
Cb_92_4 bit_92_4 gnd C_bl
Cbb_92_4 bitb_92_4 gnd C_bl
Rb_92_5 bit_92_5 bit_92_6 R_bl
Rbb_92_5 bitb_92_5 bitb_92_6 R_bl
Cb_92_5 bit_92_5 gnd C_bl
Cbb_92_5 bitb_92_5 gnd C_bl
Rb_92_6 bit_92_6 bit_92_7 R_bl
Rbb_92_6 bitb_92_6 bitb_92_7 R_bl
Cb_92_6 bit_92_6 gnd C_bl
Cbb_92_6 bitb_92_6 gnd C_bl
Rb_92_7 bit_92_7 bit_92_8 R_bl
Rbb_92_7 bitb_92_7 bitb_92_8 R_bl
Cb_92_7 bit_92_7 gnd C_bl
Cbb_92_7 bitb_92_7 gnd C_bl
Rb_92_8 bit_92_8 bit_92_9 R_bl
Rbb_92_8 bitb_92_8 bitb_92_9 R_bl
Cb_92_8 bit_92_8 gnd C_bl
Cbb_92_8 bitb_92_8 gnd C_bl
Rb_92_9 bit_92_9 bit_92_10 R_bl
Rbb_92_9 bitb_92_9 bitb_92_10 R_bl
Cb_92_9 bit_92_9 gnd C_bl
Cbb_92_9 bitb_92_9 gnd C_bl
Rb_92_10 bit_92_10 bit_92_11 R_bl
Rbb_92_10 bitb_92_10 bitb_92_11 R_bl
Cb_92_10 bit_92_10 gnd C_bl
Cbb_92_10 bitb_92_10 gnd C_bl
Rb_92_11 bit_92_11 bit_92_12 R_bl
Rbb_92_11 bitb_92_11 bitb_92_12 R_bl
Cb_92_11 bit_92_11 gnd C_bl
Cbb_92_11 bitb_92_11 gnd C_bl
Rb_92_12 bit_92_12 bit_92_13 R_bl
Rbb_92_12 bitb_92_12 bitb_92_13 R_bl
Cb_92_12 bit_92_12 gnd C_bl
Cbb_92_12 bitb_92_12 gnd C_bl
Rb_92_13 bit_92_13 bit_92_14 R_bl
Rbb_92_13 bitb_92_13 bitb_92_14 R_bl
Cb_92_13 bit_92_13 gnd C_bl
Cbb_92_13 bitb_92_13 gnd C_bl
Rb_92_14 bit_92_14 bit_92_15 R_bl
Rbb_92_14 bitb_92_14 bitb_92_15 R_bl
Cb_92_14 bit_92_14 gnd C_bl
Cbb_92_14 bitb_92_14 gnd C_bl
Rb_92_15 bit_92_15 bit_92_16 R_bl
Rbb_92_15 bitb_92_15 bitb_92_16 R_bl
Cb_92_15 bit_92_15 gnd C_bl
Cbb_92_15 bitb_92_15 gnd C_bl
Rb_92_16 bit_92_16 bit_92_17 R_bl
Rbb_92_16 bitb_92_16 bitb_92_17 R_bl
Cb_92_16 bit_92_16 gnd C_bl
Cbb_92_16 bitb_92_16 gnd C_bl
Rb_92_17 bit_92_17 bit_92_18 R_bl
Rbb_92_17 bitb_92_17 bitb_92_18 R_bl
Cb_92_17 bit_92_17 gnd C_bl
Cbb_92_17 bitb_92_17 gnd C_bl
Rb_92_18 bit_92_18 bit_92_19 R_bl
Rbb_92_18 bitb_92_18 bitb_92_19 R_bl
Cb_92_18 bit_92_18 gnd C_bl
Cbb_92_18 bitb_92_18 gnd C_bl
Rb_92_19 bit_92_19 bit_92_20 R_bl
Rbb_92_19 bitb_92_19 bitb_92_20 R_bl
Cb_92_19 bit_92_19 gnd C_bl
Cbb_92_19 bitb_92_19 gnd C_bl
Rb_92_20 bit_92_20 bit_92_21 R_bl
Rbb_92_20 bitb_92_20 bitb_92_21 R_bl
Cb_92_20 bit_92_20 gnd C_bl
Cbb_92_20 bitb_92_20 gnd C_bl
Rb_92_21 bit_92_21 bit_92_22 R_bl
Rbb_92_21 bitb_92_21 bitb_92_22 R_bl
Cb_92_21 bit_92_21 gnd C_bl
Cbb_92_21 bitb_92_21 gnd C_bl
Rb_92_22 bit_92_22 bit_92_23 R_bl
Rbb_92_22 bitb_92_22 bitb_92_23 R_bl
Cb_92_22 bit_92_22 gnd C_bl
Cbb_92_22 bitb_92_22 gnd C_bl
Rb_92_23 bit_92_23 bit_92_24 R_bl
Rbb_92_23 bitb_92_23 bitb_92_24 R_bl
Cb_92_23 bit_92_23 gnd C_bl
Cbb_92_23 bitb_92_23 gnd C_bl
Rb_92_24 bit_92_24 bit_92_25 R_bl
Rbb_92_24 bitb_92_24 bitb_92_25 R_bl
Cb_92_24 bit_92_24 gnd C_bl
Cbb_92_24 bitb_92_24 gnd C_bl
Rb_92_25 bit_92_25 bit_92_26 R_bl
Rbb_92_25 bitb_92_25 bitb_92_26 R_bl
Cb_92_25 bit_92_25 gnd C_bl
Cbb_92_25 bitb_92_25 gnd C_bl
Rb_92_26 bit_92_26 bit_92_27 R_bl
Rbb_92_26 bitb_92_26 bitb_92_27 R_bl
Cb_92_26 bit_92_26 gnd C_bl
Cbb_92_26 bitb_92_26 gnd C_bl
Rb_92_27 bit_92_27 bit_92_28 R_bl
Rbb_92_27 bitb_92_27 bitb_92_28 R_bl
Cb_92_27 bit_92_27 gnd C_bl
Cbb_92_27 bitb_92_27 gnd C_bl
Rb_92_28 bit_92_28 bit_92_29 R_bl
Rbb_92_28 bitb_92_28 bitb_92_29 R_bl
Cb_92_28 bit_92_28 gnd C_bl
Cbb_92_28 bitb_92_28 gnd C_bl
Rb_92_29 bit_92_29 bit_92_30 R_bl
Rbb_92_29 bitb_92_29 bitb_92_30 R_bl
Cb_92_29 bit_92_29 gnd C_bl
Cbb_92_29 bitb_92_29 gnd C_bl
Rb_92_30 bit_92_30 bit_92_31 R_bl
Rbb_92_30 bitb_92_30 bitb_92_31 R_bl
Cb_92_30 bit_92_30 gnd C_bl
Cbb_92_30 bitb_92_30 gnd C_bl
Rb_92_31 bit_92_31 bit_92_32 R_bl
Rbb_92_31 bitb_92_31 bitb_92_32 R_bl
Cb_92_31 bit_92_31 gnd C_bl
Cbb_92_31 bitb_92_31 gnd C_bl
Rb_92_32 bit_92_32 bit_92_33 R_bl
Rbb_92_32 bitb_92_32 bitb_92_33 R_bl
Cb_92_32 bit_92_32 gnd C_bl
Cbb_92_32 bitb_92_32 gnd C_bl
Rb_92_33 bit_92_33 bit_92_34 R_bl
Rbb_92_33 bitb_92_33 bitb_92_34 R_bl
Cb_92_33 bit_92_33 gnd C_bl
Cbb_92_33 bitb_92_33 gnd C_bl
Rb_92_34 bit_92_34 bit_92_35 R_bl
Rbb_92_34 bitb_92_34 bitb_92_35 R_bl
Cb_92_34 bit_92_34 gnd C_bl
Cbb_92_34 bitb_92_34 gnd C_bl
Rb_92_35 bit_92_35 bit_92_36 R_bl
Rbb_92_35 bitb_92_35 bitb_92_36 R_bl
Cb_92_35 bit_92_35 gnd C_bl
Cbb_92_35 bitb_92_35 gnd C_bl
Rb_92_36 bit_92_36 bit_92_37 R_bl
Rbb_92_36 bitb_92_36 bitb_92_37 R_bl
Cb_92_36 bit_92_36 gnd C_bl
Cbb_92_36 bitb_92_36 gnd C_bl
Rb_92_37 bit_92_37 bit_92_38 R_bl
Rbb_92_37 bitb_92_37 bitb_92_38 R_bl
Cb_92_37 bit_92_37 gnd C_bl
Cbb_92_37 bitb_92_37 gnd C_bl
Rb_92_38 bit_92_38 bit_92_39 R_bl
Rbb_92_38 bitb_92_38 bitb_92_39 R_bl
Cb_92_38 bit_92_38 gnd C_bl
Cbb_92_38 bitb_92_38 gnd C_bl
Rb_92_39 bit_92_39 bit_92_40 R_bl
Rbb_92_39 bitb_92_39 bitb_92_40 R_bl
Cb_92_39 bit_92_39 gnd C_bl
Cbb_92_39 bitb_92_39 gnd C_bl
Rb_92_40 bit_92_40 bit_92_41 R_bl
Rbb_92_40 bitb_92_40 bitb_92_41 R_bl
Cb_92_40 bit_92_40 gnd C_bl
Cbb_92_40 bitb_92_40 gnd C_bl
Rb_92_41 bit_92_41 bit_92_42 R_bl
Rbb_92_41 bitb_92_41 bitb_92_42 R_bl
Cb_92_41 bit_92_41 gnd C_bl
Cbb_92_41 bitb_92_41 gnd C_bl
Rb_92_42 bit_92_42 bit_92_43 R_bl
Rbb_92_42 bitb_92_42 bitb_92_43 R_bl
Cb_92_42 bit_92_42 gnd C_bl
Cbb_92_42 bitb_92_42 gnd C_bl
Rb_92_43 bit_92_43 bit_92_44 R_bl
Rbb_92_43 bitb_92_43 bitb_92_44 R_bl
Cb_92_43 bit_92_43 gnd C_bl
Cbb_92_43 bitb_92_43 gnd C_bl
Rb_92_44 bit_92_44 bit_92_45 R_bl
Rbb_92_44 bitb_92_44 bitb_92_45 R_bl
Cb_92_44 bit_92_44 gnd C_bl
Cbb_92_44 bitb_92_44 gnd C_bl
Rb_92_45 bit_92_45 bit_92_46 R_bl
Rbb_92_45 bitb_92_45 bitb_92_46 R_bl
Cb_92_45 bit_92_45 gnd C_bl
Cbb_92_45 bitb_92_45 gnd C_bl
Rb_92_46 bit_92_46 bit_92_47 R_bl
Rbb_92_46 bitb_92_46 bitb_92_47 R_bl
Cb_92_46 bit_92_46 gnd C_bl
Cbb_92_46 bitb_92_46 gnd C_bl
Rb_92_47 bit_92_47 bit_92_48 R_bl
Rbb_92_47 bitb_92_47 bitb_92_48 R_bl
Cb_92_47 bit_92_47 gnd C_bl
Cbb_92_47 bitb_92_47 gnd C_bl
Rb_92_48 bit_92_48 bit_92_49 R_bl
Rbb_92_48 bitb_92_48 bitb_92_49 R_bl
Cb_92_48 bit_92_48 gnd C_bl
Cbb_92_48 bitb_92_48 gnd C_bl
Rb_92_49 bit_92_49 bit_92_50 R_bl
Rbb_92_49 bitb_92_49 bitb_92_50 R_bl
Cb_92_49 bit_92_49 gnd C_bl
Cbb_92_49 bitb_92_49 gnd C_bl
Rb_92_50 bit_92_50 bit_92_51 R_bl
Rbb_92_50 bitb_92_50 bitb_92_51 R_bl
Cb_92_50 bit_92_50 gnd C_bl
Cbb_92_50 bitb_92_50 gnd C_bl
Rb_92_51 bit_92_51 bit_92_52 R_bl
Rbb_92_51 bitb_92_51 bitb_92_52 R_bl
Cb_92_51 bit_92_51 gnd C_bl
Cbb_92_51 bitb_92_51 gnd C_bl
Rb_92_52 bit_92_52 bit_92_53 R_bl
Rbb_92_52 bitb_92_52 bitb_92_53 R_bl
Cb_92_52 bit_92_52 gnd C_bl
Cbb_92_52 bitb_92_52 gnd C_bl
Rb_92_53 bit_92_53 bit_92_54 R_bl
Rbb_92_53 bitb_92_53 bitb_92_54 R_bl
Cb_92_53 bit_92_53 gnd C_bl
Cbb_92_53 bitb_92_53 gnd C_bl
Rb_92_54 bit_92_54 bit_92_55 R_bl
Rbb_92_54 bitb_92_54 bitb_92_55 R_bl
Cb_92_54 bit_92_54 gnd C_bl
Cbb_92_54 bitb_92_54 gnd C_bl
Rb_92_55 bit_92_55 bit_92_56 R_bl
Rbb_92_55 bitb_92_55 bitb_92_56 R_bl
Cb_92_55 bit_92_55 gnd C_bl
Cbb_92_55 bitb_92_55 gnd C_bl
Rb_92_56 bit_92_56 bit_92_57 R_bl
Rbb_92_56 bitb_92_56 bitb_92_57 R_bl
Cb_92_56 bit_92_56 gnd C_bl
Cbb_92_56 bitb_92_56 gnd C_bl
Rb_92_57 bit_92_57 bit_92_58 R_bl
Rbb_92_57 bitb_92_57 bitb_92_58 R_bl
Cb_92_57 bit_92_57 gnd C_bl
Cbb_92_57 bitb_92_57 gnd C_bl
Rb_92_58 bit_92_58 bit_92_59 R_bl
Rbb_92_58 bitb_92_58 bitb_92_59 R_bl
Cb_92_58 bit_92_58 gnd C_bl
Cbb_92_58 bitb_92_58 gnd C_bl
Rb_92_59 bit_92_59 bit_92_60 R_bl
Rbb_92_59 bitb_92_59 bitb_92_60 R_bl
Cb_92_59 bit_92_59 gnd C_bl
Cbb_92_59 bitb_92_59 gnd C_bl
Rb_92_60 bit_92_60 bit_92_61 R_bl
Rbb_92_60 bitb_92_60 bitb_92_61 R_bl
Cb_92_60 bit_92_60 gnd C_bl
Cbb_92_60 bitb_92_60 gnd C_bl
Rb_92_61 bit_92_61 bit_92_62 R_bl
Rbb_92_61 bitb_92_61 bitb_92_62 R_bl
Cb_92_61 bit_92_61 gnd C_bl
Cbb_92_61 bitb_92_61 gnd C_bl
Rb_92_62 bit_92_62 bit_92_63 R_bl
Rbb_92_62 bitb_92_62 bitb_92_63 R_bl
Cb_92_62 bit_92_62 gnd C_bl
Cbb_92_62 bitb_92_62 gnd C_bl
Rb_92_63 bit_92_63 bit_92_64 R_bl
Rbb_92_63 bitb_92_63 bitb_92_64 R_bl
Cb_92_63 bit_92_63 gnd C_bl
Cbb_92_63 bitb_92_63 gnd C_bl
Rb_92_64 bit_92_64 bit_92_65 R_bl
Rbb_92_64 bitb_92_64 bitb_92_65 R_bl
Cb_92_64 bit_92_64 gnd C_bl
Cbb_92_64 bitb_92_64 gnd C_bl
Rb_92_65 bit_92_65 bit_92_66 R_bl
Rbb_92_65 bitb_92_65 bitb_92_66 R_bl
Cb_92_65 bit_92_65 gnd C_bl
Cbb_92_65 bitb_92_65 gnd C_bl
Rb_92_66 bit_92_66 bit_92_67 R_bl
Rbb_92_66 bitb_92_66 bitb_92_67 R_bl
Cb_92_66 bit_92_66 gnd C_bl
Cbb_92_66 bitb_92_66 gnd C_bl
Rb_92_67 bit_92_67 bit_92_68 R_bl
Rbb_92_67 bitb_92_67 bitb_92_68 R_bl
Cb_92_67 bit_92_67 gnd C_bl
Cbb_92_67 bitb_92_67 gnd C_bl
Rb_92_68 bit_92_68 bit_92_69 R_bl
Rbb_92_68 bitb_92_68 bitb_92_69 R_bl
Cb_92_68 bit_92_68 gnd C_bl
Cbb_92_68 bitb_92_68 gnd C_bl
Rb_92_69 bit_92_69 bit_92_70 R_bl
Rbb_92_69 bitb_92_69 bitb_92_70 R_bl
Cb_92_69 bit_92_69 gnd C_bl
Cbb_92_69 bitb_92_69 gnd C_bl
Rb_92_70 bit_92_70 bit_92_71 R_bl
Rbb_92_70 bitb_92_70 bitb_92_71 R_bl
Cb_92_70 bit_92_70 gnd C_bl
Cbb_92_70 bitb_92_70 gnd C_bl
Rb_92_71 bit_92_71 bit_92_72 R_bl
Rbb_92_71 bitb_92_71 bitb_92_72 R_bl
Cb_92_71 bit_92_71 gnd C_bl
Cbb_92_71 bitb_92_71 gnd C_bl
Rb_92_72 bit_92_72 bit_92_73 R_bl
Rbb_92_72 bitb_92_72 bitb_92_73 R_bl
Cb_92_72 bit_92_72 gnd C_bl
Cbb_92_72 bitb_92_72 gnd C_bl
Rb_92_73 bit_92_73 bit_92_74 R_bl
Rbb_92_73 bitb_92_73 bitb_92_74 R_bl
Cb_92_73 bit_92_73 gnd C_bl
Cbb_92_73 bitb_92_73 gnd C_bl
Rb_92_74 bit_92_74 bit_92_75 R_bl
Rbb_92_74 bitb_92_74 bitb_92_75 R_bl
Cb_92_74 bit_92_74 gnd C_bl
Cbb_92_74 bitb_92_74 gnd C_bl
Rb_92_75 bit_92_75 bit_92_76 R_bl
Rbb_92_75 bitb_92_75 bitb_92_76 R_bl
Cb_92_75 bit_92_75 gnd C_bl
Cbb_92_75 bitb_92_75 gnd C_bl
Rb_92_76 bit_92_76 bit_92_77 R_bl
Rbb_92_76 bitb_92_76 bitb_92_77 R_bl
Cb_92_76 bit_92_76 gnd C_bl
Cbb_92_76 bitb_92_76 gnd C_bl
Rb_92_77 bit_92_77 bit_92_78 R_bl
Rbb_92_77 bitb_92_77 bitb_92_78 R_bl
Cb_92_77 bit_92_77 gnd C_bl
Cbb_92_77 bitb_92_77 gnd C_bl
Rb_92_78 bit_92_78 bit_92_79 R_bl
Rbb_92_78 bitb_92_78 bitb_92_79 R_bl
Cb_92_78 bit_92_78 gnd C_bl
Cbb_92_78 bitb_92_78 gnd C_bl
Rb_92_79 bit_92_79 bit_92_80 R_bl
Rbb_92_79 bitb_92_79 bitb_92_80 R_bl
Cb_92_79 bit_92_79 gnd C_bl
Cbb_92_79 bitb_92_79 gnd C_bl
Rb_92_80 bit_92_80 bit_92_81 R_bl
Rbb_92_80 bitb_92_80 bitb_92_81 R_bl
Cb_92_80 bit_92_80 gnd C_bl
Cbb_92_80 bitb_92_80 gnd C_bl
Rb_92_81 bit_92_81 bit_92_82 R_bl
Rbb_92_81 bitb_92_81 bitb_92_82 R_bl
Cb_92_81 bit_92_81 gnd C_bl
Cbb_92_81 bitb_92_81 gnd C_bl
Rb_92_82 bit_92_82 bit_92_83 R_bl
Rbb_92_82 bitb_92_82 bitb_92_83 R_bl
Cb_92_82 bit_92_82 gnd C_bl
Cbb_92_82 bitb_92_82 gnd C_bl
Rb_92_83 bit_92_83 bit_92_84 R_bl
Rbb_92_83 bitb_92_83 bitb_92_84 R_bl
Cb_92_83 bit_92_83 gnd C_bl
Cbb_92_83 bitb_92_83 gnd C_bl
Rb_92_84 bit_92_84 bit_92_85 R_bl
Rbb_92_84 bitb_92_84 bitb_92_85 R_bl
Cb_92_84 bit_92_84 gnd C_bl
Cbb_92_84 bitb_92_84 gnd C_bl
Rb_92_85 bit_92_85 bit_92_86 R_bl
Rbb_92_85 bitb_92_85 bitb_92_86 R_bl
Cb_92_85 bit_92_85 gnd C_bl
Cbb_92_85 bitb_92_85 gnd C_bl
Rb_92_86 bit_92_86 bit_92_87 R_bl
Rbb_92_86 bitb_92_86 bitb_92_87 R_bl
Cb_92_86 bit_92_86 gnd C_bl
Cbb_92_86 bitb_92_86 gnd C_bl
Rb_92_87 bit_92_87 bit_92_88 R_bl
Rbb_92_87 bitb_92_87 bitb_92_88 R_bl
Cb_92_87 bit_92_87 gnd C_bl
Cbb_92_87 bitb_92_87 gnd C_bl
Rb_92_88 bit_92_88 bit_92_89 R_bl
Rbb_92_88 bitb_92_88 bitb_92_89 R_bl
Cb_92_88 bit_92_88 gnd C_bl
Cbb_92_88 bitb_92_88 gnd C_bl
Rb_92_89 bit_92_89 bit_92_90 R_bl
Rbb_92_89 bitb_92_89 bitb_92_90 R_bl
Cb_92_89 bit_92_89 gnd C_bl
Cbb_92_89 bitb_92_89 gnd C_bl
Rb_92_90 bit_92_90 bit_92_91 R_bl
Rbb_92_90 bitb_92_90 bitb_92_91 R_bl
Cb_92_90 bit_92_90 gnd C_bl
Cbb_92_90 bitb_92_90 gnd C_bl
Rb_92_91 bit_92_91 bit_92_92 R_bl
Rbb_92_91 bitb_92_91 bitb_92_92 R_bl
Cb_92_91 bit_92_91 gnd C_bl
Cbb_92_91 bitb_92_91 gnd C_bl
Rb_92_92 bit_92_92 bit_92_93 R_bl
Rbb_92_92 bitb_92_92 bitb_92_93 R_bl
Cb_92_92 bit_92_92 gnd C_bl
Cbb_92_92 bitb_92_92 gnd C_bl
Rb_92_93 bit_92_93 bit_92_94 R_bl
Rbb_92_93 bitb_92_93 bitb_92_94 R_bl
Cb_92_93 bit_92_93 gnd C_bl
Cbb_92_93 bitb_92_93 gnd C_bl
Rb_92_94 bit_92_94 bit_92_95 R_bl
Rbb_92_94 bitb_92_94 bitb_92_95 R_bl
Cb_92_94 bit_92_94 gnd C_bl
Cbb_92_94 bitb_92_94 gnd C_bl
Rb_92_95 bit_92_95 bit_92_96 R_bl
Rbb_92_95 bitb_92_95 bitb_92_96 R_bl
Cb_92_95 bit_92_95 gnd C_bl
Cbb_92_95 bitb_92_95 gnd C_bl
Rb_92_96 bit_92_96 bit_92_97 R_bl
Rbb_92_96 bitb_92_96 bitb_92_97 R_bl
Cb_92_96 bit_92_96 gnd C_bl
Cbb_92_96 bitb_92_96 gnd C_bl
Rb_92_97 bit_92_97 bit_92_98 R_bl
Rbb_92_97 bitb_92_97 bitb_92_98 R_bl
Cb_92_97 bit_92_97 gnd C_bl
Cbb_92_97 bitb_92_97 gnd C_bl
Rb_92_98 bit_92_98 bit_92_99 R_bl
Rbb_92_98 bitb_92_98 bitb_92_99 R_bl
Cb_92_98 bit_92_98 gnd C_bl
Cbb_92_98 bitb_92_98 gnd C_bl
Rb_92_99 bit_92_99 bit_92_100 R_bl
Rbb_92_99 bitb_92_99 bitb_92_100 R_bl
Cb_92_99 bit_92_99 gnd C_bl
Cbb_92_99 bitb_92_99 gnd C_bl
Rb_93_0 bit_93_0 bit_93_1 R_bl
Rbb_93_0 bitb_93_0 bitb_93_1 R_bl
Cb_93_0 bit_93_0 gnd C_bl
Cbb_93_0 bitb_93_0 gnd C_bl
Rb_93_1 bit_93_1 bit_93_2 R_bl
Rbb_93_1 bitb_93_1 bitb_93_2 R_bl
Cb_93_1 bit_93_1 gnd C_bl
Cbb_93_1 bitb_93_1 gnd C_bl
Rb_93_2 bit_93_2 bit_93_3 R_bl
Rbb_93_2 bitb_93_2 bitb_93_3 R_bl
Cb_93_2 bit_93_2 gnd C_bl
Cbb_93_2 bitb_93_2 gnd C_bl
Rb_93_3 bit_93_3 bit_93_4 R_bl
Rbb_93_3 bitb_93_3 bitb_93_4 R_bl
Cb_93_3 bit_93_3 gnd C_bl
Cbb_93_3 bitb_93_3 gnd C_bl
Rb_93_4 bit_93_4 bit_93_5 R_bl
Rbb_93_4 bitb_93_4 bitb_93_5 R_bl
Cb_93_4 bit_93_4 gnd C_bl
Cbb_93_4 bitb_93_4 gnd C_bl
Rb_93_5 bit_93_5 bit_93_6 R_bl
Rbb_93_5 bitb_93_5 bitb_93_6 R_bl
Cb_93_5 bit_93_5 gnd C_bl
Cbb_93_5 bitb_93_5 gnd C_bl
Rb_93_6 bit_93_6 bit_93_7 R_bl
Rbb_93_6 bitb_93_6 bitb_93_7 R_bl
Cb_93_6 bit_93_6 gnd C_bl
Cbb_93_6 bitb_93_6 gnd C_bl
Rb_93_7 bit_93_7 bit_93_8 R_bl
Rbb_93_7 bitb_93_7 bitb_93_8 R_bl
Cb_93_7 bit_93_7 gnd C_bl
Cbb_93_7 bitb_93_7 gnd C_bl
Rb_93_8 bit_93_8 bit_93_9 R_bl
Rbb_93_8 bitb_93_8 bitb_93_9 R_bl
Cb_93_8 bit_93_8 gnd C_bl
Cbb_93_8 bitb_93_8 gnd C_bl
Rb_93_9 bit_93_9 bit_93_10 R_bl
Rbb_93_9 bitb_93_9 bitb_93_10 R_bl
Cb_93_9 bit_93_9 gnd C_bl
Cbb_93_9 bitb_93_9 gnd C_bl
Rb_93_10 bit_93_10 bit_93_11 R_bl
Rbb_93_10 bitb_93_10 bitb_93_11 R_bl
Cb_93_10 bit_93_10 gnd C_bl
Cbb_93_10 bitb_93_10 gnd C_bl
Rb_93_11 bit_93_11 bit_93_12 R_bl
Rbb_93_11 bitb_93_11 bitb_93_12 R_bl
Cb_93_11 bit_93_11 gnd C_bl
Cbb_93_11 bitb_93_11 gnd C_bl
Rb_93_12 bit_93_12 bit_93_13 R_bl
Rbb_93_12 bitb_93_12 bitb_93_13 R_bl
Cb_93_12 bit_93_12 gnd C_bl
Cbb_93_12 bitb_93_12 gnd C_bl
Rb_93_13 bit_93_13 bit_93_14 R_bl
Rbb_93_13 bitb_93_13 bitb_93_14 R_bl
Cb_93_13 bit_93_13 gnd C_bl
Cbb_93_13 bitb_93_13 gnd C_bl
Rb_93_14 bit_93_14 bit_93_15 R_bl
Rbb_93_14 bitb_93_14 bitb_93_15 R_bl
Cb_93_14 bit_93_14 gnd C_bl
Cbb_93_14 bitb_93_14 gnd C_bl
Rb_93_15 bit_93_15 bit_93_16 R_bl
Rbb_93_15 bitb_93_15 bitb_93_16 R_bl
Cb_93_15 bit_93_15 gnd C_bl
Cbb_93_15 bitb_93_15 gnd C_bl
Rb_93_16 bit_93_16 bit_93_17 R_bl
Rbb_93_16 bitb_93_16 bitb_93_17 R_bl
Cb_93_16 bit_93_16 gnd C_bl
Cbb_93_16 bitb_93_16 gnd C_bl
Rb_93_17 bit_93_17 bit_93_18 R_bl
Rbb_93_17 bitb_93_17 bitb_93_18 R_bl
Cb_93_17 bit_93_17 gnd C_bl
Cbb_93_17 bitb_93_17 gnd C_bl
Rb_93_18 bit_93_18 bit_93_19 R_bl
Rbb_93_18 bitb_93_18 bitb_93_19 R_bl
Cb_93_18 bit_93_18 gnd C_bl
Cbb_93_18 bitb_93_18 gnd C_bl
Rb_93_19 bit_93_19 bit_93_20 R_bl
Rbb_93_19 bitb_93_19 bitb_93_20 R_bl
Cb_93_19 bit_93_19 gnd C_bl
Cbb_93_19 bitb_93_19 gnd C_bl
Rb_93_20 bit_93_20 bit_93_21 R_bl
Rbb_93_20 bitb_93_20 bitb_93_21 R_bl
Cb_93_20 bit_93_20 gnd C_bl
Cbb_93_20 bitb_93_20 gnd C_bl
Rb_93_21 bit_93_21 bit_93_22 R_bl
Rbb_93_21 bitb_93_21 bitb_93_22 R_bl
Cb_93_21 bit_93_21 gnd C_bl
Cbb_93_21 bitb_93_21 gnd C_bl
Rb_93_22 bit_93_22 bit_93_23 R_bl
Rbb_93_22 bitb_93_22 bitb_93_23 R_bl
Cb_93_22 bit_93_22 gnd C_bl
Cbb_93_22 bitb_93_22 gnd C_bl
Rb_93_23 bit_93_23 bit_93_24 R_bl
Rbb_93_23 bitb_93_23 bitb_93_24 R_bl
Cb_93_23 bit_93_23 gnd C_bl
Cbb_93_23 bitb_93_23 gnd C_bl
Rb_93_24 bit_93_24 bit_93_25 R_bl
Rbb_93_24 bitb_93_24 bitb_93_25 R_bl
Cb_93_24 bit_93_24 gnd C_bl
Cbb_93_24 bitb_93_24 gnd C_bl
Rb_93_25 bit_93_25 bit_93_26 R_bl
Rbb_93_25 bitb_93_25 bitb_93_26 R_bl
Cb_93_25 bit_93_25 gnd C_bl
Cbb_93_25 bitb_93_25 gnd C_bl
Rb_93_26 bit_93_26 bit_93_27 R_bl
Rbb_93_26 bitb_93_26 bitb_93_27 R_bl
Cb_93_26 bit_93_26 gnd C_bl
Cbb_93_26 bitb_93_26 gnd C_bl
Rb_93_27 bit_93_27 bit_93_28 R_bl
Rbb_93_27 bitb_93_27 bitb_93_28 R_bl
Cb_93_27 bit_93_27 gnd C_bl
Cbb_93_27 bitb_93_27 gnd C_bl
Rb_93_28 bit_93_28 bit_93_29 R_bl
Rbb_93_28 bitb_93_28 bitb_93_29 R_bl
Cb_93_28 bit_93_28 gnd C_bl
Cbb_93_28 bitb_93_28 gnd C_bl
Rb_93_29 bit_93_29 bit_93_30 R_bl
Rbb_93_29 bitb_93_29 bitb_93_30 R_bl
Cb_93_29 bit_93_29 gnd C_bl
Cbb_93_29 bitb_93_29 gnd C_bl
Rb_93_30 bit_93_30 bit_93_31 R_bl
Rbb_93_30 bitb_93_30 bitb_93_31 R_bl
Cb_93_30 bit_93_30 gnd C_bl
Cbb_93_30 bitb_93_30 gnd C_bl
Rb_93_31 bit_93_31 bit_93_32 R_bl
Rbb_93_31 bitb_93_31 bitb_93_32 R_bl
Cb_93_31 bit_93_31 gnd C_bl
Cbb_93_31 bitb_93_31 gnd C_bl
Rb_93_32 bit_93_32 bit_93_33 R_bl
Rbb_93_32 bitb_93_32 bitb_93_33 R_bl
Cb_93_32 bit_93_32 gnd C_bl
Cbb_93_32 bitb_93_32 gnd C_bl
Rb_93_33 bit_93_33 bit_93_34 R_bl
Rbb_93_33 bitb_93_33 bitb_93_34 R_bl
Cb_93_33 bit_93_33 gnd C_bl
Cbb_93_33 bitb_93_33 gnd C_bl
Rb_93_34 bit_93_34 bit_93_35 R_bl
Rbb_93_34 bitb_93_34 bitb_93_35 R_bl
Cb_93_34 bit_93_34 gnd C_bl
Cbb_93_34 bitb_93_34 gnd C_bl
Rb_93_35 bit_93_35 bit_93_36 R_bl
Rbb_93_35 bitb_93_35 bitb_93_36 R_bl
Cb_93_35 bit_93_35 gnd C_bl
Cbb_93_35 bitb_93_35 gnd C_bl
Rb_93_36 bit_93_36 bit_93_37 R_bl
Rbb_93_36 bitb_93_36 bitb_93_37 R_bl
Cb_93_36 bit_93_36 gnd C_bl
Cbb_93_36 bitb_93_36 gnd C_bl
Rb_93_37 bit_93_37 bit_93_38 R_bl
Rbb_93_37 bitb_93_37 bitb_93_38 R_bl
Cb_93_37 bit_93_37 gnd C_bl
Cbb_93_37 bitb_93_37 gnd C_bl
Rb_93_38 bit_93_38 bit_93_39 R_bl
Rbb_93_38 bitb_93_38 bitb_93_39 R_bl
Cb_93_38 bit_93_38 gnd C_bl
Cbb_93_38 bitb_93_38 gnd C_bl
Rb_93_39 bit_93_39 bit_93_40 R_bl
Rbb_93_39 bitb_93_39 bitb_93_40 R_bl
Cb_93_39 bit_93_39 gnd C_bl
Cbb_93_39 bitb_93_39 gnd C_bl
Rb_93_40 bit_93_40 bit_93_41 R_bl
Rbb_93_40 bitb_93_40 bitb_93_41 R_bl
Cb_93_40 bit_93_40 gnd C_bl
Cbb_93_40 bitb_93_40 gnd C_bl
Rb_93_41 bit_93_41 bit_93_42 R_bl
Rbb_93_41 bitb_93_41 bitb_93_42 R_bl
Cb_93_41 bit_93_41 gnd C_bl
Cbb_93_41 bitb_93_41 gnd C_bl
Rb_93_42 bit_93_42 bit_93_43 R_bl
Rbb_93_42 bitb_93_42 bitb_93_43 R_bl
Cb_93_42 bit_93_42 gnd C_bl
Cbb_93_42 bitb_93_42 gnd C_bl
Rb_93_43 bit_93_43 bit_93_44 R_bl
Rbb_93_43 bitb_93_43 bitb_93_44 R_bl
Cb_93_43 bit_93_43 gnd C_bl
Cbb_93_43 bitb_93_43 gnd C_bl
Rb_93_44 bit_93_44 bit_93_45 R_bl
Rbb_93_44 bitb_93_44 bitb_93_45 R_bl
Cb_93_44 bit_93_44 gnd C_bl
Cbb_93_44 bitb_93_44 gnd C_bl
Rb_93_45 bit_93_45 bit_93_46 R_bl
Rbb_93_45 bitb_93_45 bitb_93_46 R_bl
Cb_93_45 bit_93_45 gnd C_bl
Cbb_93_45 bitb_93_45 gnd C_bl
Rb_93_46 bit_93_46 bit_93_47 R_bl
Rbb_93_46 bitb_93_46 bitb_93_47 R_bl
Cb_93_46 bit_93_46 gnd C_bl
Cbb_93_46 bitb_93_46 gnd C_bl
Rb_93_47 bit_93_47 bit_93_48 R_bl
Rbb_93_47 bitb_93_47 bitb_93_48 R_bl
Cb_93_47 bit_93_47 gnd C_bl
Cbb_93_47 bitb_93_47 gnd C_bl
Rb_93_48 bit_93_48 bit_93_49 R_bl
Rbb_93_48 bitb_93_48 bitb_93_49 R_bl
Cb_93_48 bit_93_48 gnd C_bl
Cbb_93_48 bitb_93_48 gnd C_bl
Rb_93_49 bit_93_49 bit_93_50 R_bl
Rbb_93_49 bitb_93_49 bitb_93_50 R_bl
Cb_93_49 bit_93_49 gnd C_bl
Cbb_93_49 bitb_93_49 gnd C_bl
Rb_93_50 bit_93_50 bit_93_51 R_bl
Rbb_93_50 bitb_93_50 bitb_93_51 R_bl
Cb_93_50 bit_93_50 gnd C_bl
Cbb_93_50 bitb_93_50 gnd C_bl
Rb_93_51 bit_93_51 bit_93_52 R_bl
Rbb_93_51 bitb_93_51 bitb_93_52 R_bl
Cb_93_51 bit_93_51 gnd C_bl
Cbb_93_51 bitb_93_51 gnd C_bl
Rb_93_52 bit_93_52 bit_93_53 R_bl
Rbb_93_52 bitb_93_52 bitb_93_53 R_bl
Cb_93_52 bit_93_52 gnd C_bl
Cbb_93_52 bitb_93_52 gnd C_bl
Rb_93_53 bit_93_53 bit_93_54 R_bl
Rbb_93_53 bitb_93_53 bitb_93_54 R_bl
Cb_93_53 bit_93_53 gnd C_bl
Cbb_93_53 bitb_93_53 gnd C_bl
Rb_93_54 bit_93_54 bit_93_55 R_bl
Rbb_93_54 bitb_93_54 bitb_93_55 R_bl
Cb_93_54 bit_93_54 gnd C_bl
Cbb_93_54 bitb_93_54 gnd C_bl
Rb_93_55 bit_93_55 bit_93_56 R_bl
Rbb_93_55 bitb_93_55 bitb_93_56 R_bl
Cb_93_55 bit_93_55 gnd C_bl
Cbb_93_55 bitb_93_55 gnd C_bl
Rb_93_56 bit_93_56 bit_93_57 R_bl
Rbb_93_56 bitb_93_56 bitb_93_57 R_bl
Cb_93_56 bit_93_56 gnd C_bl
Cbb_93_56 bitb_93_56 gnd C_bl
Rb_93_57 bit_93_57 bit_93_58 R_bl
Rbb_93_57 bitb_93_57 bitb_93_58 R_bl
Cb_93_57 bit_93_57 gnd C_bl
Cbb_93_57 bitb_93_57 gnd C_bl
Rb_93_58 bit_93_58 bit_93_59 R_bl
Rbb_93_58 bitb_93_58 bitb_93_59 R_bl
Cb_93_58 bit_93_58 gnd C_bl
Cbb_93_58 bitb_93_58 gnd C_bl
Rb_93_59 bit_93_59 bit_93_60 R_bl
Rbb_93_59 bitb_93_59 bitb_93_60 R_bl
Cb_93_59 bit_93_59 gnd C_bl
Cbb_93_59 bitb_93_59 gnd C_bl
Rb_93_60 bit_93_60 bit_93_61 R_bl
Rbb_93_60 bitb_93_60 bitb_93_61 R_bl
Cb_93_60 bit_93_60 gnd C_bl
Cbb_93_60 bitb_93_60 gnd C_bl
Rb_93_61 bit_93_61 bit_93_62 R_bl
Rbb_93_61 bitb_93_61 bitb_93_62 R_bl
Cb_93_61 bit_93_61 gnd C_bl
Cbb_93_61 bitb_93_61 gnd C_bl
Rb_93_62 bit_93_62 bit_93_63 R_bl
Rbb_93_62 bitb_93_62 bitb_93_63 R_bl
Cb_93_62 bit_93_62 gnd C_bl
Cbb_93_62 bitb_93_62 gnd C_bl
Rb_93_63 bit_93_63 bit_93_64 R_bl
Rbb_93_63 bitb_93_63 bitb_93_64 R_bl
Cb_93_63 bit_93_63 gnd C_bl
Cbb_93_63 bitb_93_63 gnd C_bl
Rb_93_64 bit_93_64 bit_93_65 R_bl
Rbb_93_64 bitb_93_64 bitb_93_65 R_bl
Cb_93_64 bit_93_64 gnd C_bl
Cbb_93_64 bitb_93_64 gnd C_bl
Rb_93_65 bit_93_65 bit_93_66 R_bl
Rbb_93_65 bitb_93_65 bitb_93_66 R_bl
Cb_93_65 bit_93_65 gnd C_bl
Cbb_93_65 bitb_93_65 gnd C_bl
Rb_93_66 bit_93_66 bit_93_67 R_bl
Rbb_93_66 bitb_93_66 bitb_93_67 R_bl
Cb_93_66 bit_93_66 gnd C_bl
Cbb_93_66 bitb_93_66 gnd C_bl
Rb_93_67 bit_93_67 bit_93_68 R_bl
Rbb_93_67 bitb_93_67 bitb_93_68 R_bl
Cb_93_67 bit_93_67 gnd C_bl
Cbb_93_67 bitb_93_67 gnd C_bl
Rb_93_68 bit_93_68 bit_93_69 R_bl
Rbb_93_68 bitb_93_68 bitb_93_69 R_bl
Cb_93_68 bit_93_68 gnd C_bl
Cbb_93_68 bitb_93_68 gnd C_bl
Rb_93_69 bit_93_69 bit_93_70 R_bl
Rbb_93_69 bitb_93_69 bitb_93_70 R_bl
Cb_93_69 bit_93_69 gnd C_bl
Cbb_93_69 bitb_93_69 gnd C_bl
Rb_93_70 bit_93_70 bit_93_71 R_bl
Rbb_93_70 bitb_93_70 bitb_93_71 R_bl
Cb_93_70 bit_93_70 gnd C_bl
Cbb_93_70 bitb_93_70 gnd C_bl
Rb_93_71 bit_93_71 bit_93_72 R_bl
Rbb_93_71 bitb_93_71 bitb_93_72 R_bl
Cb_93_71 bit_93_71 gnd C_bl
Cbb_93_71 bitb_93_71 gnd C_bl
Rb_93_72 bit_93_72 bit_93_73 R_bl
Rbb_93_72 bitb_93_72 bitb_93_73 R_bl
Cb_93_72 bit_93_72 gnd C_bl
Cbb_93_72 bitb_93_72 gnd C_bl
Rb_93_73 bit_93_73 bit_93_74 R_bl
Rbb_93_73 bitb_93_73 bitb_93_74 R_bl
Cb_93_73 bit_93_73 gnd C_bl
Cbb_93_73 bitb_93_73 gnd C_bl
Rb_93_74 bit_93_74 bit_93_75 R_bl
Rbb_93_74 bitb_93_74 bitb_93_75 R_bl
Cb_93_74 bit_93_74 gnd C_bl
Cbb_93_74 bitb_93_74 gnd C_bl
Rb_93_75 bit_93_75 bit_93_76 R_bl
Rbb_93_75 bitb_93_75 bitb_93_76 R_bl
Cb_93_75 bit_93_75 gnd C_bl
Cbb_93_75 bitb_93_75 gnd C_bl
Rb_93_76 bit_93_76 bit_93_77 R_bl
Rbb_93_76 bitb_93_76 bitb_93_77 R_bl
Cb_93_76 bit_93_76 gnd C_bl
Cbb_93_76 bitb_93_76 gnd C_bl
Rb_93_77 bit_93_77 bit_93_78 R_bl
Rbb_93_77 bitb_93_77 bitb_93_78 R_bl
Cb_93_77 bit_93_77 gnd C_bl
Cbb_93_77 bitb_93_77 gnd C_bl
Rb_93_78 bit_93_78 bit_93_79 R_bl
Rbb_93_78 bitb_93_78 bitb_93_79 R_bl
Cb_93_78 bit_93_78 gnd C_bl
Cbb_93_78 bitb_93_78 gnd C_bl
Rb_93_79 bit_93_79 bit_93_80 R_bl
Rbb_93_79 bitb_93_79 bitb_93_80 R_bl
Cb_93_79 bit_93_79 gnd C_bl
Cbb_93_79 bitb_93_79 gnd C_bl
Rb_93_80 bit_93_80 bit_93_81 R_bl
Rbb_93_80 bitb_93_80 bitb_93_81 R_bl
Cb_93_80 bit_93_80 gnd C_bl
Cbb_93_80 bitb_93_80 gnd C_bl
Rb_93_81 bit_93_81 bit_93_82 R_bl
Rbb_93_81 bitb_93_81 bitb_93_82 R_bl
Cb_93_81 bit_93_81 gnd C_bl
Cbb_93_81 bitb_93_81 gnd C_bl
Rb_93_82 bit_93_82 bit_93_83 R_bl
Rbb_93_82 bitb_93_82 bitb_93_83 R_bl
Cb_93_82 bit_93_82 gnd C_bl
Cbb_93_82 bitb_93_82 gnd C_bl
Rb_93_83 bit_93_83 bit_93_84 R_bl
Rbb_93_83 bitb_93_83 bitb_93_84 R_bl
Cb_93_83 bit_93_83 gnd C_bl
Cbb_93_83 bitb_93_83 gnd C_bl
Rb_93_84 bit_93_84 bit_93_85 R_bl
Rbb_93_84 bitb_93_84 bitb_93_85 R_bl
Cb_93_84 bit_93_84 gnd C_bl
Cbb_93_84 bitb_93_84 gnd C_bl
Rb_93_85 bit_93_85 bit_93_86 R_bl
Rbb_93_85 bitb_93_85 bitb_93_86 R_bl
Cb_93_85 bit_93_85 gnd C_bl
Cbb_93_85 bitb_93_85 gnd C_bl
Rb_93_86 bit_93_86 bit_93_87 R_bl
Rbb_93_86 bitb_93_86 bitb_93_87 R_bl
Cb_93_86 bit_93_86 gnd C_bl
Cbb_93_86 bitb_93_86 gnd C_bl
Rb_93_87 bit_93_87 bit_93_88 R_bl
Rbb_93_87 bitb_93_87 bitb_93_88 R_bl
Cb_93_87 bit_93_87 gnd C_bl
Cbb_93_87 bitb_93_87 gnd C_bl
Rb_93_88 bit_93_88 bit_93_89 R_bl
Rbb_93_88 bitb_93_88 bitb_93_89 R_bl
Cb_93_88 bit_93_88 gnd C_bl
Cbb_93_88 bitb_93_88 gnd C_bl
Rb_93_89 bit_93_89 bit_93_90 R_bl
Rbb_93_89 bitb_93_89 bitb_93_90 R_bl
Cb_93_89 bit_93_89 gnd C_bl
Cbb_93_89 bitb_93_89 gnd C_bl
Rb_93_90 bit_93_90 bit_93_91 R_bl
Rbb_93_90 bitb_93_90 bitb_93_91 R_bl
Cb_93_90 bit_93_90 gnd C_bl
Cbb_93_90 bitb_93_90 gnd C_bl
Rb_93_91 bit_93_91 bit_93_92 R_bl
Rbb_93_91 bitb_93_91 bitb_93_92 R_bl
Cb_93_91 bit_93_91 gnd C_bl
Cbb_93_91 bitb_93_91 gnd C_bl
Rb_93_92 bit_93_92 bit_93_93 R_bl
Rbb_93_92 bitb_93_92 bitb_93_93 R_bl
Cb_93_92 bit_93_92 gnd C_bl
Cbb_93_92 bitb_93_92 gnd C_bl
Rb_93_93 bit_93_93 bit_93_94 R_bl
Rbb_93_93 bitb_93_93 bitb_93_94 R_bl
Cb_93_93 bit_93_93 gnd C_bl
Cbb_93_93 bitb_93_93 gnd C_bl
Rb_93_94 bit_93_94 bit_93_95 R_bl
Rbb_93_94 bitb_93_94 bitb_93_95 R_bl
Cb_93_94 bit_93_94 gnd C_bl
Cbb_93_94 bitb_93_94 gnd C_bl
Rb_93_95 bit_93_95 bit_93_96 R_bl
Rbb_93_95 bitb_93_95 bitb_93_96 R_bl
Cb_93_95 bit_93_95 gnd C_bl
Cbb_93_95 bitb_93_95 gnd C_bl
Rb_93_96 bit_93_96 bit_93_97 R_bl
Rbb_93_96 bitb_93_96 bitb_93_97 R_bl
Cb_93_96 bit_93_96 gnd C_bl
Cbb_93_96 bitb_93_96 gnd C_bl
Rb_93_97 bit_93_97 bit_93_98 R_bl
Rbb_93_97 bitb_93_97 bitb_93_98 R_bl
Cb_93_97 bit_93_97 gnd C_bl
Cbb_93_97 bitb_93_97 gnd C_bl
Rb_93_98 bit_93_98 bit_93_99 R_bl
Rbb_93_98 bitb_93_98 bitb_93_99 R_bl
Cb_93_98 bit_93_98 gnd C_bl
Cbb_93_98 bitb_93_98 gnd C_bl
Rb_93_99 bit_93_99 bit_93_100 R_bl
Rbb_93_99 bitb_93_99 bitb_93_100 R_bl
Cb_93_99 bit_93_99 gnd C_bl
Cbb_93_99 bitb_93_99 gnd C_bl
Rb_94_0 bit_94_0 bit_94_1 R_bl
Rbb_94_0 bitb_94_0 bitb_94_1 R_bl
Cb_94_0 bit_94_0 gnd C_bl
Cbb_94_0 bitb_94_0 gnd C_bl
Rb_94_1 bit_94_1 bit_94_2 R_bl
Rbb_94_1 bitb_94_1 bitb_94_2 R_bl
Cb_94_1 bit_94_1 gnd C_bl
Cbb_94_1 bitb_94_1 gnd C_bl
Rb_94_2 bit_94_2 bit_94_3 R_bl
Rbb_94_2 bitb_94_2 bitb_94_3 R_bl
Cb_94_2 bit_94_2 gnd C_bl
Cbb_94_2 bitb_94_2 gnd C_bl
Rb_94_3 bit_94_3 bit_94_4 R_bl
Rbb_94_3 bitb_94_3 bitb_94_4 R_bl
Cb_94_3 bit_94_3 gnd C_bl
Cbb_94_3 bitb_94_3 gnd C_bl
Rb_94_4 bit_94_4 bit_94_5 R_bl
Rbb_94_4 bitb_94_4 bitb_94_5 R_bl
Cb_94_4 bit_94_4 gnd C_bl
Cbb_94_4 bitb_94_4 gnd C_bl
Rb_94_5 bit_94_5 bit_94_6 R_bl
Rbb_94_5 bitb_94_5 bitb_94_6 R_bl
Cb_94_5 bit_94_5 gnd C_bl
Cbb_94_5 bitb_94_5 gnd C_bl
Rb_94_6 bit_94_6 bit_94_7 R_bl
Rbb_94_6 bitb_94_6 bitb_94_7 R_bl
Cb_94_6 bit_94_6 gnd C_bl
Cbb_94_6 bitb_94_6 gnd C_bl
Rb_94_7 bit_94_7 bit_94_8 R_bl
Rbb_94_7 bitb_94_7 bitb_94_8 R_bl
Cb_94_7 bit_94_7 gnd C_bl
Cbb_94_7 bitb_94_7 gnd C_bl
Rb_94_8 bit_94_8 bit_94_9 R_bl
Rbb_94_8 bitb_94_8 bitb_94_9 R_bl
Cb_94_8 bit_94_8 gnd C_bl
Cbb_94_8 bitb_94_8 gnd C_bl
Rb_94_9 bit_94_9 bit_94_10 R_bl
Rbb_94_9 bitb_94_9 bitb_94_10 R_bl
Cb_94_9 bit_94_9 gnd C_bl
Cbb_94_9 bitb_94_9 gnd C_bl
Rb_94_10 bit_94_10 bit_94_11 R_bl
Rbb_94_10 bitb_94_10 bitb_94_11 R_bl
Cb_94_10 bit_94_10 gnd C_bl
Cbb_94_10 bitb_94_10 gnd C_bl
Rb_94_11 bit_94_11 bit_94_12 R_bl
Rbb_94_11 bitb_94_11 bitb_94_12 R_bl
Cb_94_11 bit_94_11 gnd C_bl
Cbb_94_11 bitb_94_11 gnd C_bl
Rb_94_12 bit_94_12 bit_94_13 R_bl
Rbb_94_12 bitb_94_12 bitb_94_13 R_bl
Cb_94_12 bit_94_12 gnd C_bl
Cbb_94_12 bitb_94_12 gnd C_bl
Rb_94_13 bit_94_13 bit_94_14 R_bl
Rbb_94_13 bitb_94_13 bitb_94_14 R_bl
Cb_94_13 bit_94_13 gnd C_bl
Cbb_94_13 bitb_94_13 gnd C_bl
Rb_94_14 bit_94_14 bit_94_15 R_bl
Rbb_94_14 bitb_94_14 bitb_94_15 R_bl
Cb_94_14 bit_94_14 gnd C_bl
Cbb_94_14 bitb_94_14 gnd C_bl
Rb_94_15 bit_94_15 bit_94_16 R_bl
Rbb_94_15 bitb_94_15 bitb_94_16 R_bl
Cb_94_15 bit_94_15 gnd C_bl
Cbb_94_15 bitb_94_15 gnd C_bl
Rb_94_16 bit_94_16 bit_94_17 R_bl
Rbb_94_16 bitb_94_16 bitb_94_17 R_bl
Cb_94_16 bit_94_16 gnd C_bl
Cbb_94_16 bitb_94_16 gnd C_bl
Rb_94_17 bit_94_17 bit_94_18 R_bl
Rbb_94_17 bitb_94_17 bitb_94_18 R_bl
Cb_94_17 bit_94_17 gnd C_bl
Cbb_94_17 bitb_94_17 gnd C_bl
Rb_94_18 bit_94_18 bit_94_19 R_bl
Rbb_94_18 bitb_94_18 bitb_94_19 R_bl
Cb_94_18 bit_94_18 gnd C_bl
Cbb_94_18 bitb_94_18 gnd C_bl
Rb_94_19 bit_94_19 bit_94_20 R_bl
Rbb_94_19 bitb_94_19 bitb_94_20 R_bl
Cb_94_19 bit_94_19 gnd C_bl
Cbb_94_19 bitb_94_19 gnd C_bl
Rb_94_20 bit_94_20 bit_94_21 R_bl
Rbb_94_20 bitb_94_20 bitb_94_21 R_bl
Cb_94_20 bit_94_20 gnd C_bl
Cbb_94_20 bitb_94_20 gnd C_bl
Rb_94_21 bit_94_21 bit_94_22 R_bl
Rbb_94_21 bitb_94_21 bitb_94_22 R_bl
Cb_94_21 bit_94_21 gnd C_bl
Cbb_94_21 bitb_94_21 gnd C_bl
Rb_94_22 bit_94_22 bit_94_23 R_bl
Rbb_94_22 bitb_94_22 bitb_94_23 R_bl
Cb_94_22 bit_94_22 gnd C_bl
Cbb_94_22 bitb_94_22 gnd C_bl
Rb_94_23 bit_94_23 bit_94_24 R_bl
Rbb_94_23 bitb_94_23 bitb_94_24 R_bl
Cb_94_23 bit_94_23 gnd C_bl
Cbb_94_23 bitb_94_23 gnd C_bl
Rb_94_24 bit_94_24 bit_94_25 R_bl
Rbb_94_24 bitb_94_24 bitb_94_25 R_bl
Cb_94_24 bit_94_24 gnd C_bl
Cbb_94_24 bitb_94_24 gnd C_bl
Rb_94_25 bit_94_25 bit_94_26 R_bl
Rbb_94_25 bitb_94_25 bitb_94_26 R_bl
Cb_94_25 bit_94_25 gnd C_bl
Cbb_94_25 bitb_94_25 gnd C_bl
Rb_94_26 bit_94_26 bit_94_27 R_bl
Rbb_94_26 bitb_94_26 bitb_94_27 R_bl
Cb_94_26 bit_94_26 gnd C_bl
Cbb_94_26 bitb_94_26 gnd C_bl
Rb_94_27 bit_94_27 bit_94_28 R_bl
Rbb_94_27 bitb_94_27 bitb_94_28 R_bl
Cb_94_27 bit_94_27 gnd C_bl
Cbb_94_27 bitb_94_27 gnd C_bl
Rb_94_28 bit_94_28 bit_94_29 R_bl
Rbb_94_28 bitb_94_28 bitb_94_29 R_bl
Cb_94_28 bit_94_28 gnd C_bl
Cbb_94_28 bitb_94_28 gnd C_bl
Rb_94_29 bit_94_29 bit_94_30 R_bl
Rbb_94_29 bitb_94_29 bitb_94_30 R_bl
Cb_94_29 bit_94_29 gnd C_bl
Cbb_94_29 bitb_94_29 gnd C_bl
Rb_94_30 bit_94_30 bit_94_31 R_bl
Rbb_94_30 bitb_94_30 bitb_94_31 R_bl
Cb_94_30 bit_94_30 gnd C_bl
Cbb_94_30 bitb_94_30 gnd C_bl
Rb_94_31 bit_94_31 bit_94_32 R_bl
Rbb_94_31 bitb_94_31 bitb_94_32 R_bl
Cb_94_31 bit_94_31 gnd C_bl
Cbb_94_31 bitb_94_31 gnd C_bl
Rb_94_32 bit_94_32 bit_94_33 R_bl
Rbb_94_32 bitb_94_32 bitb_94_33 R_bl
Cb_94_32 bit_94_32 gnd C_bl
Cbb_94_32 bitb_94_32 gnd C_bl
Rb_94_33 bit_94_33 bit_94_34 R_bl
Rbb_94_33 bitb_94_33 bitb_94_34 R_bl
Cb_94_33 bit_94_33 gnd C_bl
Cbb_94_33 bitb_94_33 gnd C_bl
Rb_94_34 bit_94_34 bit_94_35 R_bl
Rbb_94_34 bitb_94_34 bitb_94_35 R_bl
Cb_94_34 bit_94_34 gnd C_bl
Cbb_94_34 bitb_94_34 gnd C_bl
Rb_94_35 bit_94_35 bit_94_36 R_bl
Rbb_94_35 bitb_94_35 bitb_94_36 R_bl
Cb_94_35 bit_94_35 gnd C_bl
Cbb_94_35 bitb_94_35 gnd C_bl
Rb_94_36 bit_94_36 bit_94_37 R_bl
Rbb_94_36 bitb_94_36 bitb_94_37 R_bl
Cb_94_36 bit_94_36 gnd C_bl
Cbb_94_36 bitb_94_36 gnd C_bl
Rb_94_37 bit_94_37 bit_94_38 R_bl
Rbb_94_37 bitb_94_37 bitb_94_38 R_bl
Cb_94_37 bit_94_37 gnd C_bl
Cbb_94_37 bitb_94_37 gnd C_bl
Rb_94_38 bit_94_38 bit_94_39 R_bl
Rbb_94_38 bitb_94_38 bitb_94_39 R_bl
Cb_94_38 bit_94_38 gnd C_bl
Cbb_94_38 bitb_94_38 gnd C_bl
Rb_94_39 bit_94_39 bit_94_40 R_bl
Rbb_94_39 bitb_94_39 bitb_94_40 R_bl
Cb_94_39 bit_94_39 gnd C_bl
Cbb_94_39 bitb_94_39 gnd C_bl
Rb_94_40 bit_94_40 bit_94_41 R_bl
Rbb_94_40 bitb_94_40 bitb_94_41 R_bl
Cb_94_40 bit_94_40 gnd C_bl
Cbb_94_40 bitb_94_40 gnd C_bl
Rb_94_41 bit_94_41 bit_94_42 R_bl
Rbb_94_41 bitb_94_41 bitb_94_42 R_bl
Cb_94_41 bit_94_41 gnd C_bl
Cbb_94_41 bitb_94_41 gnd C_bl
Rb_94_42 bit_94_42 bit_94_43 R_bl
Rbb_94_42 bitb_94_42 bitb_94_43 R_bl
Cb_94_42 bit_94_42 gnd C_bl
Cbb_94_42 bitb_94_42 gnd C_bl
Rb_94_43 bit_94_43 bit_94_44 R_bl
Rbb_94_43 bitb_94_43 bitb_94_44 R_bl
Cb_94_43 bit_94_43 gnd C_bl
Cbb_94_43 bitb_94_43 gnd C_bl
Rb_94_44 bit_94_44 bit_94_45 R_bl
Rbb_94_44 bitb_94_44 bitb_94_45 R_bl
Cb_94_44 bit_94_44 gnd C_bl
Cbb_94_44 bitb_94_44 gnd C_bl
Rb_94_45 bit_94_45 bit_94_46 R_bl
Rbb_94_45 bitb_94_45 bitb_94_46 R_bl
Cb_94_45 bit_94_45 gnd C_bl
Cbb_94_45 bitb_94_45 gnd C_bl
Rb_94_46 bit_94_46 bit_94_47 R_bl
Rbb_94_46 bitb_94_46 bitb_94_47 R_bl
Cb_94_46 bit_94_46 gnd C_bl
Cbb_94_46 bitb_94_46 gnd C_bl
Rb_94_47 bit_94_47 bit_94_48 R_bl
Rbb_94_47 bitb_94_47 bitb_94_48 R_bl
Cb_94_47 bit_94_47 gnd C_bl
Cbb_94_47 bitb_94_47 gnd C_bl
Rb_94_48 bit_94_48 bit_94_49 R_bl
Rbb_94_48 bitb_94_48 bitb_94_49 R_bl
Cb_94_48 bit_94_48 gnd C_bl
Cbb_94_48 bitb_94_48 gnd C_bl
Rb_94_49 bit_94_49 bit_94_50 R_bl
Rbb_94_49 bitb_94_49 bitb_94_50 R_bl
Cb_94_49 bit_94_49 gnd C_bl
Cbb_94_49 bitb_94_49 gnd C_bl
Rb_94_50 bit_94_50 bit_94_51 R_bl
Rbb_94_50 bitb_94_50 bitb_94_51 R_bl
Cb_94_50 bit_94_50 gnd C_bl
Cbb_94_50 bitb_94_50 gnd C_bl
Rb_94_51 bit_94_51 bit_94_52 R_bl
Rbb_94_51 bitb_94_51 bitb_94_52 R_bl
Cb_94_51 bit_94_51 gnd C_bl
Cbb_94_51 bitb_94_51 gnd C_bl
Rb_94_52 bit_94_52 bit_94_53 R_bl
Rbb_94_52 bitb_94_52 bitb_94_53 R_bl
Cb_94_52 bit_94_52 gnd C_bl
Cbb_94_52 bitb_94_52 gnd C_bl
Rb_94_53 bit_94_53 bit_94_54 R_bl
Rbb_94_53 bitb_94_53 bitb_94_54 R_bl
Cb_94_53 bit_94_53 gnd C_bl
Cbb_94_53 bitb_94_53 gnd C_bl
Rb_94_54 bit_94_54 bit_94_55 R_bl
Rbb_94_54 bitb_94_54 bitb_94_55 R_bl
Cb_94_54 bit_94_54 gnd C_bl
Cbb_94_54 bitb_94_54 gnd C_bl
Rb_94_55 bit_94_55 bit_94_56 R_bl
Rbb_94_55 bitb_94_55 bitb_94_56 R_bl
Cb_94_55 bit_94_55 gnd C_bl
Cbb_94_55 bitb_94_55 gnd C_bl
Rb_94_56 bit_94_56 bit_94_57 R_bl
Rbb_94_56 bitb_94_56 bitb_94_57 R_bl
Cb_94_56 bit_94_56 gnd C_bl
Cbb_94_56 bitb_94_56 gnd C_bl
Rb_94_57 bit_94_57 bit_94_58 R_bl
Rbb_94_57 bitb_94_57 bitb_94_58 R_bl
Cb_94_57 bit_94_57 gnd C_bl
Cbb_94_57 bitb_94_57 gnd C_bl
Rb_94_58 bit_94_58 bit_94_59 R_bl
Rbb_94_58 bitb_94_58 bitb_94_59 R_bl
Cb_94_58 bit_94_58 gnd C_bl
Cbb_94_58 bitb_94_58 gnd C_bl
Rb_94_59 bit_94_59 bit_94_60 R_bl
Rbb_94_59 bitb_94_59 bitb_94_60 R_bl
Cb_94_59 bit_94_59 gnd C_bl
Cbb_94_59 bitb_94_59 gnd C_bl
Rb_94_60 bit_94_60 bit_94_61 R_bl
Rbb_94_60 bitb_94_60 bitb_94_61 R_bl
Cb_94_60 bit_94_60 gnd C_bl
Cbb_94_60 bitb_94_60 gnd C_bl
Rb_94_61 bit_94_61 bit_94_62 R_bl
Rbb_94_61 bitb_94_61 bitb_94_62 R_bl
Cb_94_61 bit_94_61 gnd C_bl
Cbb_94_61 bitb_94_61 gnd C_bl
Rb_94_62 bit_94_62 bit_94_63 R_bl
Rbb_94_62 bitb_94_62 bitb_94_63 R_bl
Cb_94_62 bit_94_62 gnd C_bl
Cbb_94_62 bitb_94_62 gnd C_bl
Rb_94_63 bit_94_63 bit_94_64 R_bl
Rbb_94_63 bitb_94_63 bitb_94_64 R_bl
Cb_94_63 bit_94_63 gnd C_bl
Cbb_94_63 bitb_94_63 gnd C_bl
Rb_94_64 bit_94_64 bit_94_65 R_bl
Rbb_94_64 bitb_94_64 bitb_94_65 R_bl
Cb_94_64 bit_94_64 gnd C_bl
Cbb_94_64 bitb_94_64 gnd C_bl
Rb_94_65 bit_94_65 bit_94_66 R_bl
Rbb_94_65 bitb_94_65 bitb_94_66 R_bl
Cb_94_65 bit_94_65 gnd C_bl
Cbb_94_65 bitb_94_65 gnd C_bl
Rb_94_66 bit_94_66 bit_94_67 R_bl
Rbb_94_66 bitb_94_66 bitb_94_67 R_bl
Cb_94_66 bit_94_66 gnd C_bl
Cbb_94_66 bitb_94_66 gnd C_bl
Rb_94_67 bit_94_67 bit_94_68 R_bl
Rbb_94_67 bitb_94_67 bitb_94_68 R_bl
Cb_94_67 bit_94_67 gnd C_bl
Cbb_94_67 bitb_94_67 gnd C_bl
Rb_94_68 bit_94_68 bit_94_69 R_bl
Rbb_94_68 bitb_94_68 bitb_94_69 R_bl
Cb_94_68 bit_94_68 gnd C_bl
Cbb_94_68 bitb_94_68 gnd C_bl
Rb_94_69 bit_94_69 bit_94_70 R_bl
Rbb_94_69 bitb_94_69 bitb_94_70 R_bl
Cb_94_69 bit_94_69 gnd C_bl
Cbb_94_69 bitb_94_69 gnd C_bl
Rb_94_70 bit_94_70 bit_94_71 R_bl
Rbb_94_70 bitb_94_70 bitb_94_71 R_bl
Cb_94_70 bit_94_70 gnd C_bl
Cbb_94_70 bitb_94_70 gnd C_bl
Rb_94_71 bit_94_71 bit_94_72 R_bl
Rbb_94_71 bitb_94_71 bitb_94_72 R_bl
Cb_94_71 bit_94_71 gnd C_bl
Cbb_94_71 bitb_94_71 gnd C_bl
Rb_94_72 bit_94_72 bit_94_73 R_bl
Rbb_94_72 bitb_94_72 bitb_94_73 R_bl
Cb_94_72 bit_94_72 gnd C_bl
Cbb_94_72 bitb_94_72 gnd C_bl
Rb_94_73 bit_94_73 bit_94_74 R_bl
Rbb_94_73 bitb_94_73 bitb_94_74 R_bl
Cb_94_73 bit_94_73 gnd C_bl
Cbb_94_73 bitb_94_73 gnd C_bl
Rb_94_74 bit_94_74 bit_94_75 R_bl
Rbb_94_74 bitb_94_74 bitb_94_75 R_bl
Cb_94_74 bit_94_74 gnd C_bl
Cbb_94_74 bitb_94_74 gnd C_bl
Rb_94_75 bit_94_75 bit_94_76 R_bl
Rbb_94_75 bitb_94_75 bitb_94_76 R_bl
Cb_94_75 bit_94_75 gnd C_bl
Cbb_94_75 bitb_94_75 gnd C_bl
Rb_94_76 bit_94_76 bit_94_77 R_bl
Rbb_94_76 bitb_94_76 bitb_94_77 R_bl
Cb_94_76 bit_94_76 gnd C_bl
Cbb_94_76 bitb_94_76 gnd C_bl
Rb_94_77 bit_94_77 bit_94_78 R_bl
Rbb_94_77 bitb_94_77 bitb_94_78 R_bl
Cb_94_77 bit_94_77 gnd C_bl
Cbb_94_77 bitb_94_77 gnd C_bl
Rb_94_78 bit_94_78 bit_94_79 R_bl
Rbb_94_78 bitb_94_78 bitb_94_79 R_bl
Cb_94_78 bit_94_78 gnd C_bl
Cbb_94_78 bitb_94_78 gnd C_bl
Rb_94_79 bit_94_79 bit_94_80 R_bl
Rbb_94_79 bitb_94_79 bitb_94_80 R_bl
Cb_94_79 bit_94_79 gnd C_bl
Cbb_94_79 bitb_94_79 gnd C_bl
Rb_94_80 bit_94_80 bit_94_81 R_bl
Rbb_94_80 bitb_94_80 bitb_94_81 R_bl
Cb_94_80 bit_94_80 gnd C_bl
Cbb_94_80 bitb_94_80 gnd C_bl
Rb_94_81 bit_94_81 bit_94_82 R_bl
Rbb_94_81 bitb_94_81 bitb_94_82 R_bl
Cb_94_81 bit_94_81 gnd C_bl
Cbb_94_81 bitb_94_81 gnd C_bl
Rb_94_82 bit_94_82 bit_94_83 R_bl
Rbb_94_82 bitb_94_82 bitb_94_83 R_bl
Cb_94_82 bit_94_82 gnd C_bl
Cbb_94_82 bitb_94_82 gnd C_bl
Rb_94_83 bit_94_83 bit_94_84 R_bl
Rbb_94_83 bitb_94_83 bitb_94_84 R_bl
Cb_94_83 bit_94_83 gnd C_bl
Cbb_94_83 bitb_94_83 gnd C_bl
Rb_94_84 bit_94_84 bit_94_85 R_bl
Rbb_94_84 bitb_94_84 bitb_94_85 R_bl
Cb_94_84 bit_94_84 gnd C_bl
Cbb_94_84 bitb_94_84 gnd C_bl
Rb_94_85 bit_94_85 bit_94_86 R_bl
Rbb_94_85 bitb_94_85 bitb_94_86 R_bl
Cb_94_85 bit_94_85 gnd C_bl
Cbb_94_85 bitb_94_85 gnd C_bl
Rb_94_86 bit_94_86 bit_94_87 R_bl
Rbb_94_86 bitb_94_86 bitb_94_87 R_bl
Cb_94_86 bit_94_86 gnd C_bl
Cbb_94_86 bitb_94_86 gnd C_bl
Rb_94_87 bit_94_87 bit_94_88 R_bl
Rbb_94_87 bitb_94_87 bitb_94_88 R_bl
Cb_94_87 bit_94_87 gnd C_bl
Cbb_94_87 bitb_94_87 gnd C_bl
Rb_94_88 bit_94_88 bit_94_89 R_bl
Rbb_94_88 bitb_94_88 bitb_94_89 R_bl
Cb_94_88 bit_94_88 gnd C_bl
Cbb_94_88 bitb_94_88 gnd C_bl
Rb_94_89 bit_94_89 bit_94_90 R_bl
Rbb_94_89 bitb_94_89 bitb_94_90 R_bl
Cb_94_89 bit_94_89 gnd C_bl
Cbb_94_89 bitb_94_89 gnd C_bl
Rb_94_90 bit_94_90 bit_94_91 R_bl
Rbb_94_90 bitb_94_90 bitb_94_91 R_bl
Cb_94_90 bit_94_90 gnd C_bl
Cbb_94_90 bitb_94_90 gnd C_bl
Rb_94_91 bit_94_91 bit_94_92 R_bl
Rbb_94_91 bitb_94_91 bitb_94_92 R_bl
Cb_94_91 bit_94_91 gnd C_bl
Cbb_94_91 bitb_94_91 gnd C_bl
Rb_94_92 bit_94_92 bit_94_93 R_bl
Rbb_94_92 bitb_94_92 bitb_94_93 R_bl
Cb_94_92 bit_94_92 gnd C_bl
Cbb_94_92 bitb_94_92 gnd C_bl
Rb_94_93 bit_94_93 bit_94_94 R_bl
Rbb_94_93 bitb_94_93 bitb_94_94 R_bl
Cb_94_93 bit_94_93 gnd C_bl
Cbb_94_93 bitb_94_93 gnd C_bl
Rb_94_94 bit_94_94 bit_94_95 R_bl
Rbb_94_94 bitb_94_94 bitb_94_95 R_bl
Cb_94_94 bit_94_94 gnd C_bl
Cbb_94_94 bitb_94_94 gnd C_bl
Rb_94_95 bit_94_95 bit_94_96 R_bl
Rbb_94_95 bitb_94_95 bitb_94_96 R_bl
Cb_94_95 bit_94_95 gnd C_bl
Cbb_94_95 bitb_94_95 gnd C_bl
Rb_94_96 bit_94_96 bit_94_97 R_bl
Rbb_94_96 bitb_94_96 bitb_94_97 R_bl
Cb_94_96 bit_94_96 gnd C_bl
Cbb_94_96 bitb_94_96 gnd C_bl
Rb_94_97 bit_94_97 bit_94_98 R_bl
Rbb_94_97 bitb_94_97 bitb_94_98 R_bl
Cb_94_97 bit_94_97 gnd C_bl
Cbb_94_97 bitb_94_97 gnd C_bl
Rb_94_98 bit_94_98 bit_94_99 R_bl
Rbb_94_98 bitb_94_98 bitb_94_99 R_bl
Cb_94_98 bit_94_98 gnd C_bl
Cbb_94_98 bitb_94_98 gnd C_bl
Rb_94_99 bit_94_99 bit_94_100 R_bl
Rbb_94_99 bitb_94_99 bitb_94_100 R_bl
Cb_94_99 bit_94_99 gnd C_bl
Cbb_94_99 bitb_94_99 gnd C_bl
Rb_95_0 bit_95_0 bit_95_1 R_bl
Rbb_95_0 bitb_95_0 bitb_95_1 R_bl
Cb_95_0 bit_95_0 gnd C_bl
Cbb_95_0 bitb_95_0 gnd C_bl
Rb_95_1 bit_95_1 bit_95_2 R_bl
Rbb_95_1 bitb_95_1 bitb_95_2 R_bl
Cb_95_1 bit_95_1 gnd C_bl
Cbb_95_1 bitb_95_1 gnd C_bl
Rb_95_2 bit_95_2 bit_95_3 R_bl
Rbb_95_2 bitb_95_2 bitb_95_3 R_bl
Cb_95_2 bit_95_2 gnd C_bl
Cbb_95_2 bitb_95_2 gnd C_bl
Rb_95_3 bit_95_3 bit_95_4 R_bl
Rbb_95_3 bitb_95_3 bitb_95_4 R_bl
Cb_95_3 bit_95_3 gnd C_bl
Cbb_95_3 bitb_95_3 gnd C_bl
Rb_95_4 bit_95_4 bit_95_5 R_bl
Rbb_95_4 bitb_95_4 bitb_95_5 R_bl
Cb_95_4 bit_95_4 gnd C_bl
Cbb_95_4 bitb_95_4 gnd C_bl
Rb_95_5 bit_95_5 bit_95_6 R_bl
Rbb_95_5 bitb_95_5 bitb_95_6 R_bl
Cb_95_5 bit_95_5 gnd C_bl
Cbb_95_5 bitb_95_5 gnd C_bl
Rb_95_6 bit_95_6 bit_95_7 R_bl
Rbb_95_6 bitb_95_6 bitb_95_7 R_bl
Cb_95_6 bit_95_6 gnd C_bl
Cbb_95_6 bitb_95_6 gnd C_bl
Rb_95_7 bit_95_7 bit_95_8 R_bl
Rbb_95_7 bitb_95_7 bitb_95_8 R_bl
Cb_95_7 bit_95_7 gnd C_bl
Cbb_95_7 bitb_95_7 gnd C_bl
Rb_95_8 bit_95_8 bit_95_9 R_bl
Rbb_95_8 bitb_95_8 bitb_95_9 R_bl
Cb_95_8 bit_95_8 gnd C_bl
Cbb_95_8 bitb_95_8 gnd C_bl
Rb_95_9 bit_95_9 bit_95_10 R_bl
Rbb_95_9 bitb_95_9 bitb_95_10 R_bl
Cb_95_9 bit_95_9 gnd C_bl
Cbb_95_9 bitb_95_9 gnd C_bl
Rb_95_10 bit_95_10 bit_95_11 R_bl
Rbb_95_10 bitb_95_10 bitb_95_11 R_bl
Cb_95_10 bit_95_10 gnd C_bl
Cbb_95_10 bitb_95_10 gnd C_bl
Rb_95_11 bit_95_11 bit_95_12 R_bl
Rbb_95_11 bitb_95_11 bitb_95_12 R_bl
Cb_95_11 bit_95_11 gnd C_bl
Cbb_95_11 bitb_95_11 gnd C_bl
Rb_95_12 bit_95_12 bit_95_13 R_bl
Rbb_95_12 bitb_95_12 bitb_95_13 R_bl
Cb_95_12 bit_95_12 gnd C_bl
Cbb_95_12 bitb_95_12 gnd C_bl
Rb_95_13 bit_95_13 bit_95_14 R_bl
Rbb_95_13 bitb_95_13 bitb_95_14 R_bl
Cb_95_13 bit_95_13 gnd C_bl
Cbb_95_13 bitb_95_13 gnd C_bl
Rb_95_14 bit_95_14 bit_95_15 R_bl
Rbb_95_14 bitb_95_14 bitb_95_15 R_bl
Cb_95_14 bit_95_14 gnd C_bl
Cbb_95_14 bitb_95_14 gnd C_bl
Rb_95_15 bit_95_15 bit_95_16 R_bl
Rbb_95_15 bitb_95_15 bitb_95_16 R_bl
Cb_95_15 bit_95_15 gnd C_bl
Cbb_95_15 bitb_95_15 gnd C_bl
Rb_95_16 bit_95_16 bit_95_17 R_bl
Rbb_95_16 bitb_95_16 bitb_95_17 R_bl
Cb_95_16 bit_95_16 gnd C_bl
Cbb_95_16 bitb_95_16 gnd C_bl
Rb_95_17 bit_95_17 bit_95_18 R_bl
Rbb_95_17 bitb_95_17 bitb_95_18 R_bl
Cb_95_17 bit_95_17 gnd C_bl
Cbb_95_17 bitb_95_17 gnd C_bl
Rb_95_18 bit_95_18 bit_95_19 R_bl
Rbb_95_18 bitb_95_18 bitb_95_19 R_bl
Cb_95_18 bit_95_18 gnd C_bl
Cbb_95_18 bitb_95_18 gnd C_bl
Rb_95_19 bit_95_19 bit_95_20 R_bl
Rbb_95_19 bitb_95_19 bitb_95_20 R_bl
Cb_95_19 bit_95_19 gnd C_bl
Cbb_95_19 bitb_95_19 gnd C_bl
Rb_95_20 bit_95_20 bit_95_21 R_bl
Rbb_95_20 bitb_95_20 bitb_95_21 R_bl
Cb_95_20 bit_95_20 gnd C_bl
Cbb_95_20 bitb_95_20 gnd C_bl
Rb_95_21 bit_95_21 bit_95_22 R_bl
Rbb_95_21 bitb_95_21 bitb_95_22 R_bl
Cb_95_21 bit_95_21 gnd C_bl
Cbb_95_21 bitb_95_21 gnd C_bl
Rb_95_22 bit_95_22 bit_95_23 R_bl
Rbb_95_22 bitb_95_22 bitb_95_23 R_bl
Cb_95_22 bit_95_22 gnd C_bl
Cbb_95_22 bitb_95_22 gnd C_bl
Rb_95_23 bit_95_23 bit_95_24 R_bl
Rbb_95_23 bitb_95_23 bitb_95_24 R_bl
Cb_95_23 bit_95_23 gnd C_bl
Cbb_95_23 bitb_95_23 gnd C_bl
Rb_95_24 bit_95_24 bit_95_25 R_bl
Rbb_95_24 bitb_95_24 bitb_95_25 R_bl
Cb_95_24 bit_95_24 gnd C_bl
Cbb_95_24 bitb_95_24 gnd C_bl
Rb_95_25 bit_95_25 bit_95_26 R_bl
Rbb_95_25 bitb_95_25 bitb_95_26 R_bl
Cb_95_25 bit_95_25 gnd C_bl
Cbb_95_25 bitb_95_25 gnd C_bl
Rb_95_26 bit_95_26 bit_95_27 R_bl
Rbb_95_26 bitb_95_26 bitb_95_27 R_bl
Cb_95_26 bit_95_26 gnd C_bl
Cbb_95_26 bitb_95_26 gnd C_bl
Rb_95_27 bit_95_27 bit_95_28 R_bl
Rbb_95_27 bitb_95_27 bitb_95_28 R_bl
Cb_95_27 bit_95_27 gnd C_bl
Cbb_95_27 bitb_95_27 gnd C_bl
Rb_95_28 bit_95_28 bit_95_29 R_bl
Rbb_95_28 bitb_95_28 bitb_95_29 R_bl
Cb_95_28 bit_95_28 gnd C_bl
Cbb_95_28 bitb_95_28 gnd C_bl
Rb_95_29 bit_95_29 bit_95_30 R_bl
Rbb_95_29 bitb_95_29 bitb_95_30 R_bl
Cb_95_29 bit_95_29 gnd C_bl
Cbb_95_29 bitb_95_29 gnd C_bl
Rb_95_30 bit_95_30 bit_95_31 R_bl
Rbb_95_30 bitb_95_30 bitb_95_31 R_bl
Cb_95_30 bit_95_30 gnd C_bl
Cbb_95_30 bitb_95_30 gnd C_bl
Rb_95_31 bit_95_31 bit_95_32 R_bl
Rbb_95_31 bitb_95_31 bitb_95_32 R_bl
Cb_95_31 bit_95_31 gnd C_bl
Cbb_95_31 bitb_95_31 gnd C_bl
Rb_95_32 bit_95_32 bit_95_33 R_bl
Rbb_95_32 bitb_95_32 bitb_95_33 R_bl
Cb_95_32 bit_95_32 gnd C_bl
Cbb_95_32 bitb_95_32 gnd C_bl
Rb_95_33 bit_95_33 bit_95_34 R_bl
Rbb_95_33 bitb_95_33 bitb_95_34 R_bl
Cb_95_33 bit_95_33 gnd C_bl
Cbb_95_33 bitb_95_33 gnd C_bl
Rb_95_34 bit_95_34 bit_95_35 R_bl
Rbb_95_34 bitb_95_34 bitb_95_35 R_bl
Cb_95_34 bit_95_34 gnd C_bl
Cbb_95_34 bitb_95_34 gnd C_bl
Rb_95_35 bit_95_35 bit_95_36 R_bl
Rbb_95_35 bitb_95_35 bitb_95_36 R_bl
Cb_95_35 bit_95_35 gnd C_bl
Cbb_95_35 bitb_95_35 gnd C_bl
Rb_95_36 bit_95_36 bit_95_37 R_bl
Rbb_95_36 bitb_95_36 bitb_95_37 R_bl
Cb_95_36 bit_95_36 gnd C_bl
Cbb_95_36 bitb_95_36 gnd C_bl
Rb_95_37 bit_95_37 bit_95_38 R_bl
Rbb_95_37 bitb_95_37 bitb_95_38 R_bl
Cb_95_37 bit_95_37 gnd C_bl
Cbb_95_37 bitb_95_37 gnd C_bl
Rb_95_38 bit_95_38 bit_95_39 R_bl
Rbb_95_38 bitb_95_38 bitb_95_39 R_bl
Cb_95_38 bit_95_38 gnd C_bl
Cbb_95_38 bitb_95_38 gnd C_bl
Rb_95_39 bit_95_39 bit_95_40 R_bl
Rbb_95_39 bitb_95_39 bitb_95_40 R_bl
Cb_95_39 bit_95_39 gnd C_bl
Cbb_95_39 bitb_95_39 gnd C_bl
Rb_95_40 bit_95_40 bit_95_41 R_bl
Rbb_95_40 bitb_95_40 bitb_95_41 R_bl
Cb_95_40 bit_95_40 gnd C_bl
Cbb_95_40 bitb_95_40 gnd C_bl
Rb_95_41 bit_95_41 bit_95_42 R_bl
Rbb_95_41 bitb_95_41 bitb_95_42 R_bl
Cb_95_41 bit_95_41 gnd C_bl
Cbb_95_41 bitb_95_41 gnd C_bl
Rb_95_42 bit_95_42 bit_95_43 R_bl
Rbb_95_42 bitb_95_42 bitb_95_43 R_bl
Cb_95_42 bit_95_42 gnd C_bl
Cbb_95_42 bitb_95_42 gnd C_bl
Rb_95_43 bit_95_43 bit_95_44 R_bl
Rbb_95_43 bitb_95_43 bitb_95_44 R_bl
Cb_95_43 bit_95_43 gnd C_bl
Cbb_95_43 bitb_95_43 gnd C_bl
Rb_95_44 bit_95_44 bit_95_45 R_bl
Rbb_95_44 bitb_95_44 bitb_95_45 R_bl
Cb_95_44 bit_95_44 gnd C_bl
Cbb_95_44 bitb_95_44 gnd C_bl
Rb_95_45 bit_95_45 bit_95_46 R_bl
Rbb_95_45 bitb_95_45 bitb_95_46 R_bl
Cb_95_45 bit_95_45 gnd C_bl
Cbb_95_45 bitb_95_45 gnd C_bl
Rb_95_46 bit_95_46 bit_95_47 R_bl
Rbb_95_46 bitb_95_46 bitb_95_47 R_bl
Cb_95_46 bit_95_46 gnd C_bl
Cbb_95_46 bitb_95_46 gnd C_bl
Rb_95_47 bit_95_47 bit_95_48 R_bl
Rbb_95_47 bitb_95_47 bitb_95_48 R_bl
Cb_95_47 bit_95_47 gnd C_bl
Cbb_95_47 bitb_95_47 gnd C_bl
Rb_95_48 bit_95_48 bit_95_49 R_bl
Rbb_95_48 bitb_95_48 bitb_95_49 R_bl
Cb_95_48 bit_95_48 gnd C_bl
Cbb_95_48 bitb_95_48 gnd C_bl
Rb_95_49 bit_95_49 bit_95_50 R_bl
Rbb_95_49 bitb_95_49 bitb_95_50 R_bl
Cb_95_49 bit_95_49 gnd C_bl
Cbb_95_49 bitb_95_49 gnd C_bl
Rb_95_50 bit_95_50 bit_95_51 R_bl
Rbb_95_50 bitb_95_50 bitb_95_51 R_bl
Cb_95_50 bit_95_50 gnd C_bl
Cbb_95_50 bitb_95_50 gnd C_bl
Rb_95_51 bit_95_51 bit_95_52 R_bl
Rbb_95_51 bitb_95_51 bitb_95_52 R_bl
Cb_95_51 bit_95_51 gnd C_bl
Cbb_95_51 bitb_95_51 gnd C_bl
Rb_95_52 bit_95_52 bit_95_53 R_bl
Rbb_95_52 bitb_95_52 bitb_95_53 R_bl
Cb_95_52 bit_95_52 gnd C_bl
Cbb_95_52 bitb_95_52 gnd C_bl
Rb_95_53 bit_95_53 bit_95_54 R_bl
Rbb_95_53 bitb_95_53 bitb_95_54 R_bl
Cb_95_53 bit_95_53 gnd C_bl
Cbb_95_53 bitb_95_53 gnd C_bl
Rb_95_54 bit_95_54 bit_95_55 R_bl
Rbb_95_54 bitb_95_54 bitb_95_55 R_bl
Cb_95_54 bit_95_54 gnd C_bl
Cbb_95_54 bitb_95_54 gnd C_bl
Rb_95_55 bit_95_55 bit_95_56 R_bl
Rbb_95_55 bitb_95_55 bitb_95_56 R_bl
Cb_95_55 bit_95_55 gnd C_bl
Cbb_95_55 bitb_95_55 gnd C_bl
Rb_95_56 bit_95_56 bit_95_57 R_bl
Rbb_95_56 bitb_95_56 bitb_95_57 R_bl
Cb_95_56 bit_95_56 gnd C_bl
Cbb_95_56 bitb_95_56 gnd C_bl
Rb_95_57 bit_95_57 bit_95_58 R_bl
Rbb_95_57 bitb_95_57 bitb_95_58 R_bl
Cb_95_57 bit_95_57 gnd C_bl
Cbb_95_57 bitb_95_57 gnd C_bl
Rb_95_58 bit_95_58 bit_95_59 R_bl
Rbb_95_58 bitb_95_58 bitb_95_59 R_bl
Cb_95_58 bit_95_58 gnd C_bl
Cbb_95_58 bitb_95_58 gnd C_bl
Rb_95_59 bit_95_59 bit_95_60 R_bl
Rbb_95_59 bitb_95_59 bitb_95_60 R_bl
Cb_95_59 bit_95_59 gnd C_bl
Cbb_95_59 bitb_95_59 gnd C_bl
Rb_95_60 bit_95_60 bit_95_61 R_bl
Rbb_95_60 bitb_95_60 bitb_95_61 R_bl
Cb_95_60 bit_95_60 gnd C_bl
Cbb_95_60 bitb_95_60 gnd C_bl
Rb_95_61 bit_95_61 bit_95_62 R_bl
Rbb_95_61 bitb_95_61 bitb_95_62 R_bl
Cb_95_61 bit_95_61 gnd C_bl
Cbb_95_61 bitb_95_61 gnd C_bl
Rb_95_62 bit_95_62 bit_95_63 R_bl
Rbb_95_62 bitb_95_62 bitb_95_63 R_bl
Cb_95_62 bit_95_62 gnd C_bl
Cbb_95_62 bitb_95_62 gnd C_bl
Rb_95_63 bit_95_63 bit_95_64 R_bl
Rbb_95_63 bitb_95_63 bitb_95_64 R_bl
Cb_95_63 bit_95_63 gnd C_bl
Cbb_95_63 bitb_95_63 gnd C_bl
Rb_95_64 bit_95_64 bit_95_65 R_bl
Rbb_95_64 bitb_95_64 bitb_95_65 R_bl
Cb_95_64 bit_95_64 gnd C_bl
Cbb_95_64 bitb_95_64 gnd C_bl
Rb_95_65 bit_95_65 bit_95_66 R_bl
Rbb_95_65 bitb_95_65 bitb_95_66 R_bl
Cb_95_65 bit_95_65 gnd C_bl
Cbb_95_65 bitb_95_65 gnd C_bl
Rb_95_66 bit_95_66 bit_95_67 R_bl
Rbb_95_66 bitb_95_66 bitb_95_67 R_bl
Cb_95_66 bit_95_66 gnd C_bl
Cbb_95_66 bitb_95_66 gnd C_bl
Rb_95_67 bit_95_67 bit_95_68 R_bl
Rbb_95_67 bitb_95_67 bitb_95_68 R_bl
Cb_95_67 bit_95_67 gnd C_bl
Cbb_95_67 bitb_95_67 gnd C_bl
Rb_95_68 bit_95_68 bit_95_69 R_bl
Rbb_95_68 bitb_95_68 bitb_95_69 R_bl
Cb_95_68 bit_95_68 gnd C_bl
Cbb_95_68 bitb_95_68 gnd C_bl
Rb_95_69 bit_95_69 bit_95_70 R_bl
Rbb_95_69 bitb_95_69 bitb_95_70 R_bl
Cb_95_69 bit_95_69 gnd C_bl
Cbb_95_69 bitb_95_69 gnd C_bl
Rb_95_70 bit_95_70 bit_95_71 R_bl
Rbb_95_70 bitb_95_70 bitb_95_71 R_bl
Cb_95_70 bit_95_70 gnd C_bl
Cbb_95_70 bitb_95_70 gnd C_bl
Rb_95_71 bit_95_71 bit_95_72 R_bl
Rbb_95_71 bitb_95_71 bitb_95_72 R_bl
Cb_95_71 bit_95_71 gnd C_bl
Cbb_95_71 bitb_95_71 gnd C_bl
Rb_95_72 bit_95_72 bit_95_73 R_bl
Rbb_95_72 bitb_95_72 bitb_95_73 R_bl
Cb_95_72 bit_95_72 gnd C_bl
Cbb_95_72 bitb_95_72 gnd C_bl
Rb_95_73 bit_95_73 bit_95_74 R_bl
Rbb_95_73 bitb_95_73 bitb_95_74 R_bl
Cb_95_73 bit_95_73 gnd C_bl
Cbb_95_73 bitb_95_73 gnd C_bl
Rb_95_74 bit_95_74 bit_95_75 R_bl
Rbb_95_74 bitb_95_74 bitb_95_75 R_bl
Cb_95_74 bit_95_74 gnd C_bl
Cbb_95_74 bitb_95_74 gnd C_bl
Rb_95_75 bit_95_75 bit_95_76 R_bl
Rbb_95_75 bitb_95_75 bitb_95_76 R_bl
Cb_95_75 bit_95_75 gnd C_bl
Cbb_95_75 bitb_95_75 gnd C_bl
Rb_95_76 bit_95_76 bit_95_77 R_bl
Rbb_95_76 bitb_95_76 bitb_95_77 R_bl
Cb_95_76 bit_95_76 gnd C_bl
Cbb_95_76 bitb_95_76 gnd C_bl
Rb_95_77 bit_95_77 bit_95_78 R_bl
Rbb_95_77 bitb_95_77 bitb_95_78 R_bl
Cb_95_77 bit_95_77 gnd C_bl
Cbb_95_77 bitb_95_77 gnd C_bl
Rb_95_78 bit_95_78 bit_95_79 R_bl
Rbb_95_78 bitb_95_78 bitb_95_79 R_bl
Cb_95_78 bit_95_78 gnd C_bl
Cbb_95_78 bitb_95_78 gnd C_bl
Rb_95_79 bit_95_79 bit_95_80 R_bl
Rbb_95_79 bitb_95_79 bitb_95_80 R_bl
Cb_95_79 bit_95_79 gnd C_bl
Cbb_95_79 bitb_95_79 gnd C_bl
Rb_95_80 bit_95_80 bit_95_81 R_bl
Rbb_95_80 bitb_95_80 bitb_95_81 R_bl
Cb_95_80 bit_95_80 gnd C_bl
Cbb_95_80 bitb_95_80 gnd C_bl
Rb_95_81 bit_95_81 bit_95_82 R_bl
Rbb_95_81 bitb_95_81 bitb_95_82 R_bl
Cb_95_81 bit_95_81 gnd C_bl
Cbb_95_81 bitb_95_81 gnd C_bl
Rb_95_82 bit_95_82 bit_95_83 R_bl
Rbb_95_82 bitb_95_82 bitb_95_83 R_bl
Cb_95_82 bit_95_82 gnd C_bl
Cbb_95_82 bitb_95_82 gnd C_bl
Rb_95_83 bit_95_83 bit_95_84 R_bl
Rbb_95_83 bitb_95_83 bitb_95_84 R_bl
Cb_95_83 bit_95_83 gnd C_bl
Cbb_95_83 bitb_95_83 gnd C_bl
Rb_95_84 bit_95_84 bit_95_85 R_bl
Rbb_95_84 bitb_95_84 bitb_95_85 R_bl
Cb_95_84 bit_95_84 gnd C_bl
Cbb_95_84 bitb_95_84 gnd C_bl
Rb_95_85 bit_95_85 bit_95_86 R_bl
Rbb_95_85 bitb_95_85 bitb_95_86 R_bl
Cb_95_85 bit_95_85 gnd C_bl
Cbb_95_85 bitb_95_85 gnd C_bl
Rb_95_86 bit_95_86 bit_95_87 R_bl
Rbb_95_86 bitb_95_86 bitb_95_87 R_bl
Cb_95_86 bit_95_86 gnd C_bl
Cbb_95_86 bitb_95_86 gnd C_bl
Rb_95_87 bit_95_87 bit_95_88 R_bl
Rbb_95_87 bitb_95_87 bitb_95_88 R_bl
Cb_95_87 bit_95_87 gnd C_bl
Cbb_95_87 bitb_95_87 gnd C_bl
Rb_95_88 bit_95_88 bit_95_89 R_bl
Rbb_95_88 bitb_95_88 bitb_95_89 R_bl
Cb_95_88 bit_95_88 gnd C_bl
Cbb_95_88 bitb_95_88 gnd C_bl
Rb_95_89 bit_95_89 bit_95_90 R_bl
Rbb_95_89 bitb_95_89 bitb_95_90 R_bl
Cb_95_89 bit_95_89 gnd C_bl
Cbb_95_89 bitb_95_89 gnd C_bl
Rb_95_90 bit_95_90 bit_95_91 R_bl
Rbb_95_90 bitb_95_90 bitb_95_91 R_bl
Cb_95_90 bit_95_90 gnd C_bl
Cbb_95_90 bitb_95_90 gnd C_bl
Rb_95_91 bit_95_91 bit_95_92 R_bl
Rbb_95_91 bitb_95_91 bitb_95_92 R_bl
Cb_95_91 bit_95_91 gnd C_bl
Cbb_95_91 bitb_95_91 gnd C_bl
Rb_95_92 bit_95_92 bit_95_93 R_bl
Rbb_95_92 bitb_95_92 bitb_95_93 R_bl
Cb_95_92 bit_95_92 gnd C_bl
Cbb_95_92 bitb_95_92 gnd C_bl
Rb_95_93 bit_95_93 bit_95_94 R_bl
Rbb_95_93 bitb_95_93 bitb_95_94 R_bl
Cb_95_93 bit_95_93 gnd C_bl
Cbb_95_93 bitb_95_93 gnd C_bl
Rb_95_94 bit_95_94 bit_95_95 R_bl
Rbb_95_94 bitb_95_94 bitb_95_95 R_bl
Cb_95_94 bit_95_94 gnd C_bl
Cbb_95_94 bitb_95_94 gnd C_bl
Rb_95_95 bit_95_95 bit_95_96 R_bl
Rbb_95_95 bitb_95_95 bitb_95_96 R_bl
Cb_95_95 bit_95_95 gnd C_bl
Cbb_95_95 bitb_95_95 gnd C_bl
Rb_95_96 bit_95_96 bit_95_97 R_bl
Rbb_95_96 bitb_95_96 bitb_95_97 R_bl
Cb_95_96 bit_95_96 gnd C_bl
Cbb_95_96 bitb_95_96 gnd C_bl
Rb_95_97 bit_95_97 bit_95_98 R_bl
Rbb_95_97 bitb_95_97 bitb_95_98 R_bl
Cb_95_97 bit_95_97 gnd C_bl
Cbb_95_97 bitb_95_97 gnd C_bl
Rb_95_98 bit_95_98 bit_95_99 R_bl
Rbb_95_98 bitb_95_98 bitb_95_99 R_bl
Cb_95_98 bit_95_98 gnd C_bl
Cbb_95_98 bitb_95_98 gnd C_bl
Rb_95_99 bit_95_99 bit_95_100 R_bl
Rbb_95_99 bitb_95_99 bitb_95_100 R_bl
Cb_95_99 bit_95_99 gnd C_bl
Cbb_95_99 bitb_95_99 gnd C_bl
Rb_96_0 bit_96_0 bit_96_1 R_bl
Rbb_96_0 bitb_96_0 bitb_96_1 R_bl
Cb_96_0 bit_96_0 gnd C_bl
Cbb_96_0 bitb_96_0 gnd C_bl
Rb_96_1 bit_96_1 bit_96_2 R_bl
Rbb_96_1 bitb_96_1 bitb_96_2 R_bl
Cb_96_1 bit_96_1 gnd C_bl
Cbb_96_1 bitb_96_1 gnd C_bl
Rb_96_2 bit_96_2 bit_96_3 R_bl
Rbb_96_2 bitb_96_2 bitb_96_3 R_bl
Cb_96_2 bit_96_2 gnd C_bl
Cbb_96_2 bitb_96_2 gnd C_bl
Rb_96_3 bit_96_3 bit_96_4 R_bl
Rbb_96_3 bitb_96_3 bitb_96_4 R_bl
Cb_96_3 bit_96_3 gnd C_bl
Cbb_96_3 bitb_96_3 gnd C_bl
Rb_96_4 bit_96_4 bit_96_5 R_bl
Rbb_96_4 bitb_96_4 bitb_96_5 R_bl
Cb_96_4 bit_96_4 gnd C_bl
Cbb_96_4 bitb_96_4 gnd C_bl
Rb_96_5 bit_96_5 bit_96_6 R_bl
Rbb_96_5 bitb_96_5 bitb_96_6 R_bl
Cb_96_5 bit_96_5 gnd C_bl
Cbb_96_5 bitb_96_5 gnd C_bl
Rb_96_6 bit_96_6 bit_96_7 R_bl
Rbb_96_6 bitb_96_6 bitb_96_7 R_bl
Cb_96_6 bit_96_6 gnd C_bl
Cbb_96_6 bitb_96_6 gnd C_bl
Rb_96_7 bit_96_7 bit_96_8 R_bl
Rbb_96_7 bitb_96_7 bitb_96_8 R_bl
Cb_96_7 bit_96_7 gnd C_bl
Cbb_96_7 bitb_96_7 gnd C_bl
Rb_96_8 bit_96_8 bit_96_9 R_bl
Rbb_96_8 bitb_96_8 bitb_96_9 R_bl
Cb_96_8 bit_96_8 gnd C_bl
Cbb_96_8 bitb_96_8 gnd C_bl
Rb_96_9 bit_96_9 bit_96_10 R_bl
Rbb_96_9 bitb_96_9 bitb_96_10 R_bl
Cb_96_9 bit_96_9 gnd C_bl
Cbb_96_9 bitb_96_9 gnd C_bl
Rb_96_10 bit_96_10 bit_96_11 R_bl
Rbb_96_10 bitb_96_10 bitb_96_11 R_bl
Cb_96_10 bit_96_10 gnd C_bl
Cbb_96_10 bitb_96_10 gnd C_bl
Rb_96_11 bit_96_11 bit_96_12 R_bl
Rbb_96_11 bitb_96_11 bitb_96_12 R_bl
Cb_96_11 bit_96_11 gnd C_bl
Cbb_96_11 bitb_96_11 gnd C_bl
Rb_96_12 bit_96_12 bit_96_13 R_bl
Rbb_96_12 bitb_96_12 bitb_96_13 R_bl
Cb_96_12 bit_96_12 gnd C_bl
Cbb_96_12 bitb_96_12 gnd C_bl
Rb_96_13 bit_96_13 bit_96_14 R_bl
Rbb_96_13 bitb_96_13 bitb_96_14 R_bl
Cb_96_13 bit_96_13 gnd C_bl
Cbb_96_13 bitb_96_13 gnd C_bl
Rb_96_14 bit_96_14 bit_96_15 R_bl
Rbb_96_14 bitb_96_14 bitb_96_15 R_bl
Cb_96_14 bit_96_14 gnd C_bl
Cbb_96_14 bitb_96_14 gnd C_bl
Rb_96_15 bit_96_15 bit_96_16 R_bl
Rbb_96_15 bitb_96_15 bitb_96_16 R_bl
Cb_96_15 bit_96_15 gnd C_bl
Cbb_96_15 bitb_96_15 gnd C_bl
Rb_96_16 bit_96_16 bit_96_17 R_bl
Rbb_96_16 bitb_96_16 bitb_96_17 R_bl
Cb_96_16 bit_96_16 gnd C_bl
Cbb_96_16 bitb_96_16 gnd C_bl
Rb_96_17 bit_96_17 bit_96_18 R_bl
Rbb_96_17 bitb_96_17 bitb_96_18 R_bl
Cb_96_17 bit_96_17 gnd C_bl
Cbb_96_17 bitb_96_17 gnd C_bl
Rb_96_18 bit_96_18 bit_96_19 R_bl
Rbb_96_18 bitb_96_18 bitb_96_19 R_bl
Cb_96_18 bit_96_18 gnd C_bl
Cbb_96_18 bitb_96_18 gnd C_bl
Rb_96_19 bit_96_19 bit_96_20 R_bl
Rbb_96_19 bitb_96_19 bitb_96_20 R_bl
Cb_96_19 bit_96_19 gnd C_bl
Cbb_96_19 bitb_96_19 gnd C_bl
Rb_96_20 bit_96_20 bit_96_21 R_bl
Rbb_96_20 bitb_96_20 bitb_96_21 R_bl
Cb_96_20 bit_96_20 gnd C_bl
Cbb_96_20 bitb_96_20 gnd C_bl
Rb_96_21 bit_96_21 bit_96_22 R_bl
Rbb_96_21 bitb_96_21 bitb_96_22 R_bl
Cb_96_21 bit_96_21 gnd C_bl
Cbb_96_21 bitb_96_21 gnd C_bl
Rb_96_22 bit_96_22 bit_96_23 R_bl
Rbb_96_22 bitb_96_22 bitb_96_23 R_bl
Cb_96_22 bit_96_22 gnd C_bl
Cbb_96_22 bitb_96_22 gnd C_bl
Rb_96_23 bit_96_23 bit_96_24 R_bl
Rbb_96_23 bitb_96_23 bitb_96_24 R_bl
Cb_96_23 bit_96_23 gnd C_bl
Cbb_96_23 bitb_96_23 gnd C_bl
Rb_96_24 bit_96_24 bit_96_25 R_bl
Rbb_96_24 bitb_96_24 bitb_96_25 R_bl
Cb_96_24 bit_96_24 gnd C_bl
Cbb_96_24 bitb_96_24 gnd C_bl
Rb_96_25 bit_96_25 bit_96_26 R_bl
Rbb_96_25 bitb_96_25 bitb_96_26 R_bl
Cb_96_25 bit_96_25 gnd C_bl
Cbb_96_25 bitb_96_25 gnd C_bl
Rb_96_26 bit_96_26 bit_96_27 R_bl
Rbb_96_26 bitb_96_26 bitb_96_27 R_bl
Cb_96_26 bit_96_26 gnd C_bl
Cbb_96_26 bitb_96_26 gnd C_bl
Rb_96_27 bit_96_27 bit_96_28 R_bl
Rbb_96_27 bitb_96_27 bitb_96_28 R_bl
Cb_96_27 bit_96_27 gnd C_bl
Cbb_96_27 bitb_96_27 gnd C_bl
Rb_96_28 bit_96_28 bit_96_29 R_bl
Rbb_96_28 bitb_96_28 bitb_96_29 R_bl
Cb_96_28 bit_96_28 gnd C_bl
Cbb_96_28 bitb_96_28 gnd C_bl
Rb_96_29 bit_96_29 bit_96_30 R_bl
Rbb_96_29 bitb_96_29 bitb_96_30 R_bl
Cb_96_29 bit_96_29 gnd C_bl
Cbb_96_29 bitb_96_29 gnd C_bl
Rb_96_30 bit_96_30 bit_96_31 R_bl
Rbb_96_30 bitb_96_30 bitb_96_31 R_bl
Cb_96_30 bit_96_30 gnd C_bl
Cbb_96_30 bitb_96_30 gnd C_bl
Rb_96_31 bit_96_31 bit_96_32 R_bl
Rbb_96_31 bitb_96_31 bitb_96_32 R_bl
Cb_96_31 bit_96_31 gnd C_bl
Cbb_96_31 bitb_96_31 gnd C_bl
Rb_96_32 bit_96_32 bit_96_33 R_bl
Rbb_96_32 bitb_96_32 bitb_96_33 R_bl
Cb_96_32 bit_96_32 gnd C_bl
Cbb_96_32 bitb_96_32 gnd C_bl
Rb_96_33 bit_96_33 bit_96_34 R_bl
Rbb_96_33 bitb_96_33 bitb_96_34 R_bl
Cb_96_33 bit_96_33 gnd C_bl
Cbb_96_33 bitb_96_33 gnd C_bl
Rb_96_34 bit_96_34 bit_96_35 R_bl
Rbb_96_34 bitb_96_34 bitb_96_35 R_bl
Cb_96_34 bit_96_34 gnd C_bl
Cbb_96_34 bitb_96_34 gnd C_bl
Rb_96_35 bit_96_35 bit_96_36 R_bl
Rbb_96_35 bitb_96_35 bitb_96_36 R_bl
Cb_96_35 bit_96_35 gnd C_bl
Cbb_96_35 bitb_96_35 gnd C_bl
Rb_96_36 bit_96_36 bit_96_37 R_bl
Rbb_96_36 bitb_96_36 bitb_96_37 R_bl
Cb_96_36 bit_96_36 gnd C_bl
Cbb_96_36 bitb_96_36 gnd C_bl
Rb_96_37 bit_96_37 bit_96_38 R_bl
Rbb_96_37 bitb_96_37 bitb_96_38 R_bl
Cb_96_37 bit_96_37 gnd C_bl
Cbb_96_37 bitb_96_37 gnd C_bl
Rb_96_38 bit_96_38 bit_96_39 R_bl
Rbb_96_38 bitb_96_38 bitb_96_39 R_bl
Cb_96_38 bit_96_38 gnd C_bl
Cbb_96_38 bitb_96_38 gnd C_bl
Rb_96_39 bit_96_39 bit_96_40 R_bl
Rbb_96_39 bitb_96_39 bitb_96_40 R_bl
Cb_96_39 bit_96_39 gnd C_bl
Cbb_96_39 bitb_96_39 gnd C_bl
Rb_96_40 bit_96_40 bit_96_41 R_bl
Rbb_96_40 bitb_96_40 bitb_96_41 R_bl
Cb_96_40 bit_96_40 gnd C_bl
Cbb_96_40 bitb_96_40 gnd C_bl
Rb_96_41 bit_96_41 bit_96_42 R_bl
Rbb_96_41 bitb_96_41 bitb_96_42 R_bl
Cb_96_41 bit_96_41 gnd C_bl
Cbb_96_41 bitb_96_41 gnd C_bl
Rb_96_42 bit_96_42 bit_96_43 R_bl
Rbb_96_42 bitb_96_42 bitb_96_43 R_bl
Cb_96_42 bit_96_42 gnd C_bl
Cbb_96_42 bitb_96_42 gnd C_bl
Rb_96_43 bit_96_43 bit_96_44 R_bl
Rbb_96_43 bitb_96_43 bitb_96_44 R_bl
Cb_96_43 bit_96_43 gnd C_bl
Cbb_96_43 bitb_96_43 gnd C_bl
Rb_96_44 bit_96_44 bit_96_45 R_bl
Rbb_96_44 bitb_96_44 bitb_96_45 R_bl
Cb_96_44 bit_96_44 gnd C_bl
Cbb_96_44 bitb_96_44 gnd C_bl
Rb_96_45 bit_96_45 bit_96_46 R_bl
Rbb_96_45 bitb_96_45 bitb_96_46 R_bl
Cb_96_45 bit_96_45 gnd C_bl
Cbb_96_45 bitb_96_45 gnd C_bl
Rb_96_46 bit_96_46 bit_96_47 R_bl
Rbb_96_46 bitb_96_46 bitb_96_47 R_bl
Cb_96_46 bit_96_46 gnd C_bl
Cbb_96_46 bitb_96_46 gnd C_bl
Rb_96_47 bit_96_47 bit_96_48 R_bl
Rbb_96_47 bitb_96_47 bitb_96_48 R_bl
Cb_96_47 bit_96_47 gnd C_bl
Cbb_96_47 bitb_96_47 gnd C_bl
Rb_96_48 bit_96_48 bit_96_49 R_bl
Rbb_96_48 bitb_96_48 bitb_96_49 R_bl
Cb_96_48 bit_96_48 gnd C_bl
Cbb_96_48 bitb_96_48 gnd C_bl
Rb_96_49 bit_96_49 bit_96_50 R_bl
Rbb_96_49 bitb_96_49 bitb_96_50 R_bl
Cb_96_49 bit_96_49 gnd C_bl
Cbb_96_49 bitb_96_49 gnd C_bl
Rb_96_50 bit_96_50 bit_96_51 R_bl
Rbb_96_50 bitb_96_50 bitb_96_51 R_bl
Cb_96_50 bit_96_50 gnd C_bl
Cbb_96_50 bitb_96_50 gnd C_bl
Rb_96_51 bit_96_51 bit_96_52 R_bl
Rbb_96_51 bitb_96_51 bitb_96_52 R_bl
Cb_96_51 bit_96_51 gnd C_bl
Cbb_96_51 bitb_96_51 gnd C_bl
Rb_96_52 bit_96_52 bit_96_53 R_bl
Rbb_96_52 bitb_96_52 bitb_96_53 R_bl
Cb_96_52 bit_96_52 gnd C_bl
Cbb_96_52 bitb_96_52 gnd C_bl
Rb_96_53 bit_96_53 bit_96_54 R_bl
Rbb_96_53 bitb_96_53 bitb_96_54 R_bl
Cb_96_53 bit_96_53 gnd C_bl
Cbb_96_53 bitb_96_53 gnd C_bl
Rb_96_54 bit_96_54 bit_96_55 R_bl
Rbb_96_54 bitb_96_54 bitb_96_55 R_bl
Cb_96_54 bit_96_54 gnd C_bl
Cbb_96_54 bitb_96_54 gnd C_bl
Rb_96_55 bit_96_55 bit_96_56 R_bl
Rbb_96_55 bitb_96_55 bitb_96_56 R_bl
Cb_96_55 bit_96_55 gnd C_bl
Cbb_96_55 bitb_96_55 gnd C_bl
Rb_96_56 bit_96_56 bit_96_57 R_bl
Rbb_96_56 bitb_96_56 bitb_96_57 R_bl
Cb_96_56 bit_96_56 gnd C_bl
Cbb_96_56 bitb_96_56 gnd C_bl
Rb_96_57 bit_96_57 bit_96_58 R_bl
Rbb_96_57 bitb_96_57 bitb_96_58 R_bl
Cb_96_57 bit_96_57 gnd C_bl
Cbb_96_57 bitb_96_57 gnd C_bl
Rb_96_58 bit_96_58 bit_96_59 R_bl
Rbb_96_58 bitb_96_58 bitb_96_59 R_bl
Cb_96_58 bit_96_58 gnd C_bl
Cbb_96_58 bitb_96_58 gnd C_bl
Rb_96_59 bit_96_59 bit_96_60 R_bl
Rbb_96_59 bitb_96_59 bitb_96_60 R_bl
Cb_96_59 bit_96_59 gnd C_bl
Cbb_96_59 bitb_96_59 gnd C_bl
Rb_96_60 bit_96_60 bit_96_61 R_bl
Rbb_96_60 bitb_96_60 bitb_96_61 R_bl
Cb_96_60 bit_96_60 gnd C_bl
Cbb_96_60 bitb_96_60 gnd C_bl
Rb_96_61 bit_96_61 bit_96_62 R_bl
Rbb_96_61 bitb_96_61 bitb_96_62 R_bl
Cb_96_61 bit_96_61 gnd C_bl
Cbb_96_61 bitb_96_61 gnd C_bl
Rb_96_62 bit_96_62 bit_96_63 R_bl
Rbb_96_62 bitb_96_62 bitb_96_63 R_bl
Cb_96_62 bit_96_62 gnd C_bl
Cbb_96_62 bitb_96_62 gnd C_bl
Rb_96_63 bit_96_63 bit_96_64 R_bl
Rbb_96_63 bitb_96_63 bitb_96_64 R_bl
Cb_96_63 bit_96_63 gnd C_bl
Cbb_96_63 bitb_96_63 gnd C_bl
Rb_96_64 bit_96_64 bit_96_65 R_bl
Rbb_96_64 bitb_96_64 bitb_96_65 R_bl
Cb_96_64 bit_96_64 gnd C_bl
Cbb_96_64 bitb_96_64 gnd C_bl
Rb_96_65 bit_96_65 bit_96_66 R_bl
Rbb_96_65 bitb_96_65 bitb_96_66 R_bl
Cb_96_65 bit_96_65 gnd C_bl
Cbb_96_65 bitb_96_65 gnd C_bl
Rb_96_66 bit_96_66 bit_96_67 R_bl
Rbb_96_66 bitb_96_66 bitb_96_67 R_bl
Cb_96_66 bit_96_66 gnd C_bl
Cbb_96_66 bitb_96_66 gnd C_bl
Rb_96_67 bit_96_67 bit_96_68 R_bl
Rbb_96_67 bitb_96_67 bitb_96_68 R_bl
Cb_96_67 bit_96_67 gnd C_bl
Cbb_96_67 bitb_96_67 gnd C_bl
Rb_96_68 bit_96_68 bit_96_69 R_bl
Rbb_96_68 bitb_96_68 bitb_96_69 R_bl
Cb_96_68 bit_96_68 gnd C_bl
Cbb_96_68 bitb_96_68 gnd C_bl
Rb_96_69 bit_96_69 bit_96_70 R_bl
Rbb_96_69 bitb_96_69 bitb_96_70 R_bl
Cb_96_69 bit_96_69 gnd C_bl
Cbb_96_69 bitb_96_69 gnd C_bl
Rb_96_70 bit_96_70 bit_96_71 R_bl
Rbb_96_70 bitb_96_70 bitb_96_71 R_bl
Cb_96_70 bit_96_70 gnd C_bl
Cbb_96_70 bitb_96_70 gnd C_bl
Rb_96_71 bit_96_71 bit_96_72 R_bl
Rbb_96_71 bitb_96_71 bitb_96_72 R_bl
Cb_96_71 bit_96_71 gnd C_bl
Cbb_96_71 bitb_96_71 gnd C_bl
Rb_96_72 bit_96_72 bit_96_73 R_bl
Rbb_96_72 bitb_96_72 bitb_96_73 R_bl
Cb_96_72 bit_96_72 gnd C_bl
Cbb_96_72 bitb_96_72 gnd C_bl
Rb_96_73 bit_96_73 bit_96_74 R_bl
Rbb_96_73 bitb_96_73 bitb_96_74 R_bl
Cb_96_73 bit_96_73 gnd C_bl
Cbb_96_73 bitb_96_73 gnd C_bl
Rb_96_74 bit_96_74 bit_96_75 R_bl
Rbb_96_74 bitb_96_74 bitb_96_75 R_bl
Cb_96_74 bit_96_74 gnd C_bl
Cbb_96_74 bitb_96_74 gnd C_bl
Rb_96_75 bit_96_75 bit_96_76 R_bl
Rbb_96_75 bitb_96_75 bitb_96_76 R_bl
Cb_96_75 bit_96_75 gnd C_bl
Cbb_96_75 bitb_96_75 gnd C_bl
Rb_96_76 bit_96_76 bit_96_77 R_bl
Rbb_96_76 bitb_96_76 bitb_96_77 R_bl
Cb_96_76 bit_96_76 gnd C_bl
Cbb_96_76 bitb_96_76 gnd C_bl
Rb_96_77 bit_96_77 bit_96_78 R_bl
Rbb_96_77 bitb_96_77 bitb_96_78 R_bl
Cb_96_77 bit_96_77 gnd C_bl
Cbb_96_77 bitb_96_77 gnd C_bl
Rb_96_78 bit_96_78 bit_96_79 R_bl
Rbb_96_78 bitb_96_78 bitb_96_79 R_bl
Cb_96_78 bit_96_78 gnd C_bl
Cbb_96_78 bitb_96_78 gnd C_bl
Rb_96_79 bit_96_79 bit_96_80 R_bl
Rbb_96_79 bitb_96_79 bitb_96_80 R_bl
Cb_96_79 bit_96_79 gnd C_bl
Cbb_96_79 bitb_96_79 gnd C_bl
Rb_96_80 bit_96_80 bit_96_81 R_bl
Rbb_96_80 bitb_96_80 bitb_96_81 R_bl
Cb_96_80 bit_96_80 gnd C_bl
Cbb_96_80 bitb_96_80 gnd C_bl
Rb_96_81 bit_96_81 bit_96_82 R_bl
Rbb_96_81 bitb_96_81 bitb_96_82 R_bl
Cb_96_81 bit_96_81 gnd C_bl
Cbb_96_81 bitb_96_81 gnd C_bl
Rb_96_82 bit_96_82 bit_96_83 R_bl
Rbb_96_82 bitb_96_82 bitb_96_83 R_bl
Cb_96_82 bit_96_82 gnd C_bl
Cbb_96_82 bitb_96_82 gnd C_bl
Rb_96_83 bit_96_83 bit_96_84 R_bl
Rbb_96_83 bitb_96_83 bitb_96_84 R_bl
Cb_96_83 bit_96_83 gnd C_bl
Cbb_96_83 bitb_96_83 gnd C_bl
Rb_96_84 bit_96_84 bit_96_85 R_bl
Rbb_96_84 bitb_96_84 bitb_96_85 R_bl
Cb_96_84 bit_96_84 gnd C_bl
Cbb_96_84 bitb_96_84 gnd C_bl
Rb_96_85 bit_96_85 bit_96_86 R_bl
Rbb_96_85 bitb_96_85 bitb_96_86 R_bl
Cb_96_85 bit_96_85 gnd C_bl
Cbb_96_85 bitb_96_85 gnd C_bl
Rb_96_86 bit_96_86 bit_96_87 R_bl
Rbb_96_86 bitb_96_86 bitb_96_87 R_bl
Cb_96_86 bit_96_86 gnd C_bl
Cbb_96_86 bitb_96_86 gnd C_bl
Rb_96_87 bit_96_87 bit_96_88 R_bl
Rbb_96_87 bitb_96_87 bitb_96_88 R_bl
Cb_96_87 bit_96_87 gnd C_bl
Cbb_96_87 bitb_96_87 gnd C_bl
Rb_96_88 bit_96_88 bit_96_89 R_bl
Rbb_96_88 bitb_96_88 bitb_96_89 R_bl
Cb_96_88 bit_96_88 gnd C_bl
Cbb_96_88 bitb_96_88 gnd C_bl
Rb_96_89 bit_96_89 bit_96_90 R_bl
Rbb_96_89 bitb_96_89 bitb_96_90 R_bl
Cb_96_89 bit_96_89 gnd C_bl
Cbb_96_89 bitb_96_89 gnd C_bl
Rb_96_90 bit_96_90 bit_96_91 R_bl
Rbb_96_90 bitb_96_90 bitb_96_91 R_bl
Cb_96_90 bit_96_90 gnd C_bl
Cbb_96_90 bitb_96_90 gnd C_bl
Rb_96_91 bit_96_91 bit_96_92 R_bl
Rbb_96_91 bitb_96_91 bitb_96_92 R_bl
Cb_96_91 bit_96_91 gnd C_bl
Cbb_96_91 bitb_96_91 gnd C_bl
Rb_96_92 bit_96_92 bit_96_93 R_bl
Rbb_96_92 bitb_96_92 bitb_96_93 R_bl
Cb_96_92 bit_96_92 gnd C_bl
Cbb_96_92 bitb_96_92 gnd C_bl
Rb_96_93 bit_96_93 bit_96_94 R_bl
Rbb_96_93 bitb_96_93 bitb_96_94 R_bl
Cb_96_93 bit_96_93 gnd C_bl
Cbb_96_93 bitb_96_93 gnd C_bl
Rb_96_94 bit_96_94 bit_96_95 R_bl
Rbb_96_94 bitb_96_94 bitb_96_95 R_bl
Cb_96_94 bit_96_94 gnd C_bl
Cbb_96_94 bitb_96_94 gnd C_bl
Rb_96_95 bit_96_95 bit_96_96 R_bl
Rbb_96_95 bitb_96_95 bitb_96_96 R_bl
Cb_96_95 bit_96_95 gnd C_bl
Cbb_96_95 bitb_96_95 gnd C_bl
Rb_96_96 bit_96_96 bit_96_97 R_bl
Rbb_96_96 bitb_96_96 bitb_96_97 R_bl
Cb_96_96 bit_96_96 gnd C_bl
Cbb_96_96 bitb_96_96 gnd C_bl
Rb_96_97 bit_96_97 bit_96_98 R_bl
Rbb_96_97 bitb_96_97 bitb_96_98 R_bl
Cb_96_97 bit_96_97 gnd C_bl
Cbb_96_97 bitb_96_97 gnd C_bl
Rb_96_98 bit_96_98 bit_96_99 R_bl
Rbb_96_98 bitb_96_98 bitb_96_99 R_bl
Cb_96_98 bit_96_98 gnd C_bl
Cbb_96_98 bitb_96_98 gnd C_bl
Rb_96_99 bit_96_99 bit_96_100 R_bl
Rbb_96_99 bitb_96_99 bitb_96_100 R_bl
Cb_96_99 bit_96_99 gnd C_bl
Cbb_96_99 bitb_96_99 gnd C_bl
Rb_97_0 bit_97_0 bit_97_1 R_bl
Rbb_97_0 bitb_97_0 bitb_97_1 R_bl
Cb_97_0 bit_97_0 gnd C_bl
Cbb_97_0 bitb_97_0 gnd C_bl
Rb_97_1 bit_97_1 bit_97_2 R_bl
Rbb_97_1 bitb_97_1 bitb_97_2 R_bl
Cb_97_1 bit_97_1 gnd C_bl
Cbb_97_1 bitb_97_1 gnd C_bl
Rb_97_2 bit_97_2 bit_97_3 R_bl
Rbb_97_2 bitb_97_2 bitb_97_3 R_bl
Cb_97_2 bit_97_2 gnd C_bl
Cbb_97_2 bitb_97_2 gnd C_bl
Rb_97_3 bit_97_3 bit_97_4 R_bl
Rbb_97_3 bitb_97_3 bitb_97_4 R_bl
Cb_97_3 bit_97_3 gnd C_bl
Cbb_97_3 bitb_97_3 gnd C_bl
Rb_97_4 bit_97_4 bit_97_5 R_bl
Rbb_97_4 bitb_97_4 bitb_97_5 R_bl
Cb_97_4 bit_97_4 gnd C_bl
Cbb_97_4 bitb_97_4 gnd C_bl
Rb_97_5 bit_97_5 bit_97_6 R_bl
Rbb_97_5 bitb_97_5 bitb_97_6 R_bl
Cb_97_5 bit_97_5 gnd C_bl
Cbb_97_5 bitb_97_5 gnd C_bl
Rb_97_6 bit_97_6 bit_97_7 R_bl
Rbb_97_6 bitb_97_6 bitb_97_7 R_bl
Cb_97_6 bit_97_6 gnd C_bl
Cbb_97_6 bitb_97_6 gnd C_bl
Rb_97_7 bit_97_7 bit_97_8 R_bl
Rbb_97_7 bitb_97_7 bitb_97_8 R_bl
Cb_97_7 bit_97_7 gnd C_bl
Cbb_97_7 bitb_97_7 gnd C_bl
Rb_97_8 bit_97_8 bit_97_9 R_bl
Rbb_97_8 bitb_97_8 bitb_97_9 R_bl
Cb_97_8 bit_97_8 gnd C_bl
Cbb_97_8 bitb_97_8 gnd C_bl
Rb_97_9 bit_97_9 bit_97_10 R_bl
Rbb_97_9 bitb_97_9 bitb_97_10 R_bl
Cb_97_9 bit_97_9 gnd C_bl
Cbb_97_9 bitb_97_9 gnd C_bl
Rb_97_10 bit_97_10 bit_97_11 R_bl
Rbb_97_10 bitb_97_10 bitb_97_11 R_bl
Cb_97_10 bit_97_10 gnd C_bl
Cbb_97_10 bitb_97_10 gnd C_bl
Rb_97_11 bit_97_11 bit_97_12 R_bl
Rbb_97_11 bitb_97_11 bitb_97_12 R_bl
Cb_97_11 bit_97_11 gnd C_bl
Cbb_97_11 bitb_97_11 gnd C_bl
Rb_97_12 bit_97_12 bit_97_13 R_bl
Rbb_97_12 bitb_97_12 bitb_97_13 R_bl
Cb_97_12 bit_97_12 gnd C_bl
Cbb_97_12 bitb_97_12 gnd C_bl
Rb_97_13 bit_97_13 bit_97_14 R_bl
Rbb_97_13 bitb_97_13 bitb_97_14 R_bl
Cb_97_13 bit_97_13 gnd C_bl
Cbb_97_13 bitb_97_13 gnd C_bl
Rb_97_14 bit_97_14 bit_97_15 R_bl
Rbb_97_14 bitb_97_14 bitb_97_15 R_bl
Cb_97_14 bit_97_14 gnd C_bl
Cbb_97_14 bitb_97_14 gnd C_bl
Rb_97_15 bit_97_15 bit_97_16 R_bl
Rbb_97_15 bitb_97_15 bitb_97_16 R_bl
Cb_97_15 bit_97_15 gnd C_bl
Cbb_97_15 bitb_97_15 gnd C_bl
Rb_97_16 bit_97_16 bit_97_17 R_bl
Rbb_97_16 bitb_97_16 bitb_97_17 R_bl
Cb_97_16 bit_97_16 gnd C_bl
Cbb_97_16 bitb_97_16 gnd C_bl
Rb_97_17 bit_97_17 bit_97_18 R_bl
Rbb_97_17 bitb_97_17 bitb_97_18 R_bl
Cb_97_17 bit_97_17 gnd C_bl
Cbb_97_17 bitb_97_17 gnd C_bl
Rb_97_18 bit_97_18 bit_97_19 R_bl
Rbb_97_18 bitb_97_18 bitb_97_19 R_bl
Cb_97_18 bit_97_18 gnd C_bl
Cbb_97_18 bitb_97_18 gnd C_bl
Rb_97_19 bit_97_19 bit_97_20 R_bl
Rbb_97_19 bitb_97_19 bitb_97_20 R_bl
Cb_97_19 bit_97_19 gnd C_bl
Cbb_97_19 bitb_97_19 gnd C_bl
Rb_97_20 bit_97_20 bit_97_21 R_bl
Rbb_97_20 bitb_97_20 bitb_97_21 R_bl
Cb_97_20 bit_97_20 gnd C_bl
Cbb_97_20 bitb_97_20 gnd C_bl
Rb_97_21 bit_97_21 bit_97_22 R_bl
Rbb_97_21 bitb_97_21 bitb_97_22 R_bl
Cb_97_21 bit_97_21 gnd C_bl
Cbb_97_21 bitb_97_21 gnd C_bl
Rb_97_22 bit_97_22 bit_97_23 R_bl
Rbb_97_22 bitb_97_22 bitb_97_23 R_bl
Cb_97_22 bit_97_22 gnd C_bl
Cbb_97_22 bitb_97_22 gnd C_bl
Rb_97_23 bit_97_23 bit_97_24 R_bl
Rbb_97_23 bitb_97_23 bitb_97_24 R_bl
Cb_97_23 bit_97_23 gnd C_bl
Cbb_97_23 bitb_97_23 gnd C_bl
Rb_97_24 bit_97_24 bit_97_25 R_bl
Rbb_97_24 bitb_97_24 bitb_97_25 R_bl
Cb_97_24 bit_97_24 gnd C_bl
Cbb_97_24 bitb_97_24 gnd C_bl
Rb_97_25 bit_97_25 bit_97_26 R_bl
Rbb_97_25 bitb_97_25 bitb_97_26 R_bl
Cb_97_25 bit_97_25 gnd C_bl
Cbb_97_25 bitb_97_25 gnd C_bl
Rb_97_26 bit_97_26 bit_97_27 R_bl
Rbb_97_26 bitb_97_26 bitb_97_27 R_bl
Cb_97_26 bit_97_26 gnd C_bl
Cbb_97_26 bitb_97_26 gnd C_bl
Rb_97_27 bit_97_27 bit_97_28 R_bl
Rbb_97_27 bitb_97_27 bitb_97_28 R_bl
Cb_97_27 bit_97_27 gnd C_bl
Cbb_97_27 bitb_97_27 gnd C_bl
Rb_97_28 bit_97_28 bit_97_29 R_bl
Rbb_97_28 bitb_97_28 bitb_97_29 R_bl
Cb_97_28 bit_97_28 gnd C_bl
Cbb_97_28 bitb_97_28 gnd C_bl
Rb_97_29 bit_97_29 bit_97_30 R_bl
Rbb_97_29 bitb_97_29 bitb_97_30 R_bl
Cb_97_29 bit_97_29 gnd C_bl
Cbb_97_29 bitb_97_29 gnd C_bl
Rb_97_30 bit_97_30 bit_97_31 R_bl
Rbb_97_30 bitb_97_30 bitb_97_31 R_bl
Cb_97_30 bit_97_30 gnd C_bl
Cbb_97_30 bitb_97_30 gnd C_bl
Rb_97_31 bit_97_31 bit_97_32 R_bl
Rbb_97_31 bitb_97_31 bitb_97_32 R_bl
Cb_97_31 bit_97_31 gnd C_bl
Cbb_97_31 bitb_97_31 gnd C_bl
Rb_97_32 bit_97_32 bit_97_33 R_bl
Rbb_97_32 bitb_97_32 bitb_97_33 R_bl
Cb_97_32 bit_97_32 gnd C_bl
Cbb_97_32 bitb_97_32 gnd C_bl
Rb_97_33 bit_97_33 bit_97_34 R_bl
Rbb_97_33 bitb_97_33 bitb_97_34 R_bl
Cb_97_33 bit_97_33 gnd C_bl
Cbb_97_33 bitb_97_33 gnd C_bl
Rb_97_34 bit_97_34 bit_97_35 R_bl
Rbb_97_34 bitb_97_34 bitb_97_35 R_bl
Cb_97_34 bit_97_34 gnd C_bl
Cbb_97_34 bitb_97_34 gnd C_bl
Rb_97_35 bit_97_35 bit_97_36 R_bl
Rbb_97_35 bitb_97_35 bitb_97_36 R_bl
Cb_97_35 bit_97_35 gnd C_bl
Cbb_97_35 bitb_97_35 gnd C_bl
Rb_97_36 bit_97_36 bit_97_37 R_bl
Rbb_97_36 bitb_97_36 bitb_97_37 R_bl
Cb_97_36 bit_97_36 gnd C_bl
Cbb_97_36 bitb_97_36 gnd C_bl
Rb_97_37 bit_97_37 bit_97_38 R_bl
Rbb_97_37 bitb_97_37 bitb_97_38 R_bl
Cb_97_37 bit_97_37 gnd C_bl
Cbb_97_37 bitb_97_37 gnd C_bl
Rb_97_38 bit_97_38 bit_97_39 R_bl
Rbb_97_38 bitb_97_38 bitb_97_39 R_bl
Cb_97_38 bit_97_38 gnd C_bl
Cbb_97_38 bitb_97_38 gnd C_bl
Rb_97_39 bit_97_39 bit_97_40 R_bl
Rbb_97_39 bitb_97_39 bitb_97_40 R_bl
Cb_97_39 bit_97_39 gnd C_bl
Cbb_97_39 bitb_97_39 gnd C_bl
Rb_97_40 bit_97_40 bit_97_41 R_bl
Rbb_97_40 bitb_97_40 bitb_97_41 R_bl
Cb_97_40 bit_97_40 gnd C_bl
Cbb_97_40 bitb_97_40 gnd C_bl
Rb_97_41 bit_97_41 bit_97_42 R_bl
Rbb_97_41 bitb_97_41 bitb_97_42 R_bl
Cb_97_41 bit_97_41 gnd C_bl
Cbb_97_41 bitb_97_41 gnd C_bl
Rb_97_42 bit_97_42 bit_97_43 R_bl
Rbb_97_42 bitb_97_42 bitb_97_43 R_bl
Cb_97_42 bit_97_42 gnd C_bl
Cbb_97_42 bitb_97_42 gnd C_bl
Rb_97_43 bit_97_43 bit_97_44 R_bl
Rbb_97_43 bitb_97_43 bitb_97_44 R_bl
Cb_97_43 bit_97_43 gnd C_bl
Cbb_97_43 bitb_97_43 gnd C_bl
Rb_97_44 bit_97_44 bit_97_45 R_bl
Rbb_97_44 bitb_97_44 bitb_97_45 R_bl
Cb_97_44 bit_97_44 gnd C_bl
Cbb_97_44 bitb_97_44 gnd C_bl
Rb_97_45 bit_97_45 bit_97_46 R_bl
Rbb_97_45 bitb_97_45 bitb_97_46 R_bl
Cb_97_45 bit_97_45 gnd C_bl
Cbb_97_45 bitb_97_45 gnd C_bl
Rb_97_46 bit_97_46 bit_97_47 R_bl
Rbb_97_46 bitb_97_46 bitb_97_47 R_bl
Cb_97_46 bit_97_46 gnd C_bl
Cbb_97_46 bitb_97_46 gnd C_bl
Rb_97_47 bit_97_47 bit_97_48 R_bl
Rbb_97_47 bitb_97_47 bitb_97_48 R_bl
Cb_97_47 bit_97_47 gnd C_bl
Cbb_97_47 bitb_97_47 gnd C_bl
Rb_97_48 bit_97_48 bit_97_49 R_bl
Rbb_97_48 bitb_97_48 bitb_97_49 R_bl
Cb_97_48 bit_97_48 gnd C_bl
Cbb_97_48 bitb_97_48 gnd C_bl
Rb_97_49 bit_97_49 bit_97_50 R_bl
Rbb_97_49 bitb_97_49 bitb_97_50 R_bl
Cb_97_49 bit_97_49 gnd C_bl
Cbb_97_49 bitb_97_49 gnd C_bl
Rb_97_50 bit_97_50 bit_97_51 R_bl
Rbb_97_50 bitb_97_50 bitb_97_51 R_bl
Cb_97_50 bit_97_50 gnd C_bl
Cbb_97_50 bitb_97_50 gnd C_bl
Rb_97_51 bit_97_51 bit_97_52 R_bl
Rbb_97_51 bitb_97_51 bitb_97_52 R_bl
Cb_97_51 bit_97_51 gnd C_bl
Cbb_97_51 bitb_97_51 gnd C_bl
Rb_97_52 bit_97_52 bit_97_53 R_bl
Rbb_97_52 bitb_97_52 bitb_97_53 R_bl
Cb_97_52 bit_97_52 gnd C_bl
Cbb_97_52 bitb_97_52 gnd C_bl
Rb_97_53 bit_97_53 bit_97_54 R_bl
Rbb_97_53 bitb_97_53 bitb_97_54 R_bl
Cb_97_53 bit_97_53 gnd C_bl
Cbb_97_53 bitb_97_53 gnd C_bl
Rb_97_54 bit_97_54 bit_97_55 R_bl
Rbb_97_54 bitb_97_54 bitb_97_55 R_bl
Cb_97_54 bit_97_54 gnd C_bl
Cbb_97_54 bitb_97_54 gnd C_bl
Rb_97_55 bit_97_55 bit_97_56 R_bl
Rbb_97_55 bitb_97_55 bitb_97_56 R_bl
Cb_97_55 bit_97_55 gnd C_bl
Cbb_97_55 bitb_97_55 gnd C_bl
Rb_97_56 bit_97_56 bit_97_57 R_bl
Rbb_97_56 bitb_97_56 bitb_97_57 R_bl
Cb_97_56 bit_97_56 gnd C_bl
Cbb_97_56 bitb_97_56 gnd C_bl
Rb_97_57 bit_97_57 bit_97_58 R_bl
Rbb_97_57 bitb_97_57 bitb_97_58 R_bl
Cb_97_57 bit_97_57 gnd C_bl
Cbb_97_57 bitb_97_57 gnd C_bl
Rb_97_58 bit_97_58 bit_97_59 R_bl
Rbb_97_58 bitb_97_58 bitb_97_59 R_bl
Cb_97_58 bit_97_58 gnd C_bl
Cbb_97_58 bitb_97_58 gnd C_bl
Rb_97_59 bit_97_59 bit_97_60 R_bl
Rbb_97_59 bitb_97_59 bitb_97_60 R_bl
Cb_97_59 bit_97_59 gnd C_bl
Cbb_97_59 bitb_97_59 gnd C_bl
Rb_97_60 bit_97_60 bit_97_61 R_bl
Rbb_97_60 bitb_97_60 bitb_97_61 R_bl
Cb_97_60 bit_97_60 gnd C_bl
Cbb_97_60 bitb_97_60 gnd C_bl
Rb_97_61 bit_97_61 bit_97_62 R_bl
Rbb_97_61 bitb_97_61 bitb_97_62 R_bl
Cb_97_61 bit_97_61 gnd C_bl
Cbb_97_61 bitb_97_61 gnd C_bl
Rb_97_62 bit_97_62 bit_97_63 R_bl
Rbb_97_62 bitb_97_62 bitb_97_63 R_bl
Cb_97_62 bit_97_62 gnd C_bl
Cbb_97_62 bitb_97_62 gnd C_bl
Rb_97_63 bit_97_63 bit_97_64 R_bl
Rbb_97_63 bitb_97_63 bitb_97_64 R_bl
Cb_97_63 bit_97_63 gnd C_bl
Cbb_97_63 bitb_97_63 gnd C_bl
Rb_97_64 bit_97_64 bit_97_65 R_bl
Rbb_97_64 bitb_97_64 bitb_97_65 R_bl
Cb_97_64 bit_97_64 gnd C_bl
Cbb_97_64 bitb_97_64 gnd C_bl
Rb_97_65 bit_97_65 bit_97_66 R_bl
Rbb_97_65 bitb_97_65 bitb_97_66 R_bl
Cb_97_65 bit_97_65 gnd C_bl
Cbb_97_65 bitb_97_65 gnd C_bl
Rb_97_66 bit_97_66 bit_97_67 R_bl
Rbb_97_66 bitb_97_66 bitb_97_67 R_bl
Cb_97_66 bit_97_66 gnd C_bl
Cbb_97_66 bitb_97_66 gnd C_bl
Rb_97_67 bit_97_67 bit_97_68 R_bl
Rbb_97_67 bitb_97_67 bitb_97_68 R_bl
Cb_97_67 bit_97_67 gnd C_bl
Cbb_97_67 bitb_97_67 gnd C_bl
Rb_97_68 bit_97_68 bit_97_69 R_bl
Rbb_97_68 bitb_97_68 bitb_97_69 R_bl
Cb_97_68 bit_97_68 gnd C_bl
Cbb_97_68 bitb_97_68 gnd C_bl
Rb_97_69 bit_97_69 bit_97_70 R_bl
Rbb_97_69 bitb_97_69 bitb_97_70 R_bl
Cb_97_69 bit_97_69 gnd C_bl
Cbb_97_69 bitb_97_69 gnd C_bl
Rb_97_70 bit_97_70 bit_97_71 R_bl
Rbb_97_70 bitb_97_70 bitb_97_71 R_bl
Cb_97_70 bit_97_70 gnd C_bl
Cbb_97_70 bitb_97_70 gnd C_bl
Rb_97_71 bit_97_71 bit_97_72 R_bl
Rbb_97_71 bitb_97_71 bitb_97_72 R_bl
Cb_97_71 bit_97_71 gnd C_bl
Cbb_97_71 bitb_97_71 gnd C_bl
Rb_97_72 bit_97_72 bit_97_73 R_bl
Rbb_97_72 bitb_97_72 bitb_97_73 R_bl
Cb_97_72 bit_97_72 gnd C_bl
Cbb_97_72 bitb_97_72 gnd C_bl
Rb_97_73 bit_97_73 bit_97_74 R_bl
Rbb_97_73 bitb_97_73 bitb_97_74 R_bl
Cb_97_73 bit_97_73 gnd C_bl
Cbb_97_73 bitb_97_73 gnd C_bl
Rb_97_74 bit_97_74 bit_97_75 R_bl
Rbb_97_74 bitb_97_74 bitb_97_75 R_bl
Cb_97_74 bit_97_74 gnd C_bl
Cbb_97_74 bitb_97_74 gnd C_bl
Rb_97_75 bit_97_75 bit_97_76 R_bl
Rbb_97_75 bitb_97_75 bitb_97_76 R_bl
Cb_97_75 bit_97_75 gnd C_bl
Cbb_97_75 bitb_97_75 gnd C_bl
Rb_97_76 bit_97_76 bit_97_77 R_bl
Rbb_97_76 bitb_97_76 bitb_97_77 R_bl
Cb_97_76 bit_97_76 gnd C_bl
Cbb_97_76 bitb_97_76 gnd C_bl
Rb_97_77 bit_97_77 bit_97_78 R_bl
Rbb_97_77 bitb_97_77 bitb_97_78 R_bl
Cb_97_77 bit_97_77 gnd C_bl
Cbb_97_77 bitb_97_77 gnd C_bl
Rb_97_78 bit_97_78 bit_97_79 R_bl
Rbb_97_78 bitb_97_78 bitb_97_79 R_bl
Cb_97_78 bit_97_78 gnd C_bl
Cbb_97_78 bitb_97_78 gnd C_bl
Rb_97_79 bit_97_79 bit_97_80 R_bl
Rbb_97_79 bitb_97_79 bitb_97_80 R_bl
Cb_97_79 bit_97_79 gnd C_bl
Cbb_97_79 bitb_97_79 gnd C_bl
Rb_97_80 bit_97_80 bit_97_81 R_bl
Rbb_97_80 bitb_97_80 bitb_97_81 R_bl
Cb_97_80 bit_97_80 gnd C_bl
Cbb_97_80 bitb_97_80 gnd C_bl
Rb_97_81 bit_97_81 bit_97_82 R_bl
Rbb_97_81 bitb_97_81 bitb_97_82 R_bl
Cb_97_81 bit_97_81 gnd C_bl
Cbb_97_81 bitb_97_81 gnd C_bl
Rb_97_82 bit_97_82 bit_97_83 R_bl
Rbb_97_82 bitb_97_82 bitb_97_83 R_bl
Cb_97_82 bit_97_82 gnd C_bl
Cbb_97_82 bitb_97_82 gnd C_bl
Rb_97_83 bit_97_83 bit_97_84 R_bl
Rbb_97_83 bitb_97_83 bitb_97_84 R_bl
Cb_97_83 bit_97_83 gnd C_bl
Cbb_97_83 bitb_97_83 gnd C_bl
Rb_97_84 bit_97_84 bit_97_85 R_bl
Rbb_97_84 bitb_97_84 bitb_97_85 R_bl
Cb_97_84 bit_97_84 gnd C_bl
Cbb_97_84 bitb_97_84 gnd C_bl
Rb_97_85 bit_97_85 bit_97_86 R_bl
Rbb_97_85 bitb_97_85 bitb_97_86 R_bl
Cb_97_85 bit_97_85 gnd C_bl
Cbb_97_85 bitb_97_85 gnd C_bl
Rb_97_86 bit_97_86 bit_97_87 R_bl
Rbb_97_86 bitb_97_86 bitb_97_87 R_bl
Cb_97_86 bit_97_86 gnd C_bl
Cbb_97_86 bitb_97_86 gnd C_bl
Rb_97_87 bit_97_87 bit_97_88 R_bl
Rbb_97_87 bitb_97_87 bitb_97_88 R_bl
Cb_97_87 bit_97_87 gnd C_bl
Cbb_97_87 bitb_97_87 gnd C_bl
Rb_97_88 bit_97_88 bit_97_89 R_bl
Rbb_97_88 bitb_97_88 bitb_97_89 R_bl
Cb_97_88 bit_97_88 gnd C_bl
Cbb_97_88 bitb_97_88 gnd C_bl
Rb_97_89 bit_97_89 bit_97_90 R_bl
Rbb_97_89 bitb_97_89 bitb_97_90 R_bl
Cb_97_89 bit_97_89 gnd C_bl
Cbb_97_89 bitb_97_89 gnd C_bl
Rb_97_90 bit_97_90 bit_97_91 R_bl
Rbb_97_90 bitb_97_90 bitb_97_91 R_bl
Cb_97_90 bit_97_90 gnd C_bl
Cbb_97_90 bitb_97_90 gnd C_bl
Rb_97_91 bit_97_91 bit_97_92 R_bl
Rbb_97_91 bitb_97_91 bitb_97_92 R_bl
Cb_97_91 bit_97_91 gnd C_bl
Cbb_97_91 bitb_97_91 gnd C_bl
Rb_97_92 bit_97_92 bit_97_93 R_bl
Rbb_97_92 bitb_97_92 bitb_97_93 R_bl
Cb_97_92 bit_97_92 gnd C_bl
Cbb_97_92 bitb_97_92 gnd C_bl
Rb_97_93 bit_97_93 bit_97_94 R_bl
Rbb_97_93 bitb_97_93 bitb_97_94 R_bl
Cb_97_93 bit_97_93 gnd C_bl
Cbb_97_93 bitb_97_93 gnd C_bl
Rb_97_94 bit_97_94 bit_97_95 R_bl
Rbb_97_94 bitb_97_94 bitb_97_95 R_bl
Cb_97_94 bit_97_94 gnd C_bl
Cbb_97_94 bitb_97_94 gnd C_bl
Rb_97_95 bit_97_95 bit_97_96 R_bl
Rbb_97_95 bitb_97_95 bitb_97_96 R_bl
Cb_97_95 bit_97_95 gnd C_bl
Cbb_97_95 bitb_97_95 gnd C_bl
Rb_97_96 bit_97_96 bit_97_97 R_bl
Rbb_97_96 bitb_97_96 bitb_97_97 R_bl
Cb_97_96 bit_97_96 gnd C_bl
Cbb_97_96 bitb_97_96 gnd C_bl
Rb_97_97 bit_97_97 bit_97_98 R_bl
Rbb_97_97 bitb_97_97 bitb_97_98 R_bl
Cb_97_97 bit_97_97 gnd C_bl
Cbb_97_97 bitb_97_97 gnd C_bl
Rb_97_98 bit_97_98 bit_97_99 R_bl
Rbb_97_98 bitb_97_98 bitb_97_99 R_bl
Cb_97_98 bit_97_98 gnd C_bl
Cbb_97_98 bitb_97_98 gnd C_bl
Rb_97_99 bit_97_99 bit_97_100 R_bl
Rbb_97_99 bitb_97_99 bitb_97_100 R_bl
Cb_97_99 bit_97_99 gnd C_bl
Cbb_97_99 bitb_97_99 gnd C_bl
Rb_98_0 bit_98_0 bit_98_1 R_bl
Rbb_98_0 bitb_98_0 bitb_98_1 R_bl
Cb_98_0 bit_98_0 gnd C_bl
Cbb_98_0 bitb_98_0 gnd C_bl
Rb_98_1 bit_98_1 bit_98_2 R_bl
Rbb_98_1 bitb_98_1 bitb_98_2 R_bl
Cb_98_1 bit_98_1 gnd C_bl
Cbb_98_1 bitb_98_1 gnd C_bl
Rb_98_2 bit_98_2 bit_98_3 R_bl
Rbb_98_2 bitb_98_2 bitb_98_3 R_bl
Cb_98_2 bit_98_2 gnd C_bl
Cbb_98_2 bitb_98_2 gnd C_bl
Rb_98_3 bit_98_3 bit_98_4 R_bl
Rbb_98_3 bitb_98_3 bitb_98_4 R_bl
Cb_98_3 bit_98_3 gnd C_bl
Cbb_98_3 bitb_98_3 gnd C_bl
Rb_98_4 bit_98_4 bit_98_5 R_bl
Rbb_98_4 bitb_98_4 bitb_98_5 R_bl
Cb_98_4 bit_98_4 gnd C_bl
Cbb_98_4 bitb_98_4 gnd C_bl
Rb_98_5 bit_98_5 bit_98_6 R_bl
Rbb_98_5 bitb_98_5 bitb_98_6 R_bl
Cb_98_5 bit_98_5 gnd C_bl
Cbb_98_5 bitb_98_5 gnd C_bl
Rb_98_6 bit_98_6 bit_98_7 R_bl
Rbb_98_6 bitb_98_6 bitb_98_7 R_bl
Cb_98_6 bit_98_6 gnd C_bl
Cbb_98_6 bitb_98_6 gnd C_bl
Rb_98_7 bit_98_7 bit_98_8 R_bl
Rbb_98_7 bitb_98_7 bitb_98_8 R_bl
Cb_98_7 bit_98_7 gnd C_bl
Cbb_98_7 bitb_98_7 gnd C_bl
Rb_98_8 bit_98_8 bit_98_9 R_bl
Rbb_98_8 bitb_98_8 bitb_98_9 R_bl
Cb_98_8 bit_98_8 gnd C_bl
Cbb_98_8 bitb_98_8 gnd C_bl
Rb_98_9 bit_98_9 bit_98_10 R_bl
Rbb_98_9 bitb_98_9 bitb_98_10 R_bl
Cb_98_9 bit_98_9 gnd C_bl
Cbb_98_9 bitb_98_9 gnd C_bl
Rb_98_10 bit_98_10 bit_98_11 R_bl
Rbb_98_10 bitb_98_10 bitb_98_11 R_bl
Cb_98_10 bit_98_10 gnd C_bl
Cbb_98_10 bitb_98_10 gnd C_bl
Rb_98_11 bit_98_11 bit_98_12 R_bl
Rbb_98_11 bitb_98_11 bitb_98_12 R_bl
Cb_98_11 bit_98_11 gnd C_bl
Cbb_98_11 bitb_98_11 gnd C_bl
Rb_98_12 bit_98_12 bit_98_13 R_bl
Rbb_98_12 bitb_98_12 bitb_98_13 R_bl
Cb_98_12 bit_98_12 gnd C_bl
Cbb_98_12 bitb_98_12 gnd C_bl
Rb_98_13 bit_98_13 bit_98_14 R_bl
Rbb_98_13 bitb_98_13 bitb_98_14 R_bl
Cb_98_13 bit_98_13 gnd C_bl
Cbb_98_13 bitb_98_13 gnd C_bl
Rb_98_14 bit_98_14 bit_98_15 R_bl
Rbb_98_14 bitb_98_14 bitb_98_15 R_bl
Cb_98_14 bit_98_14 gnd C_bl
Cbb_98_14 bitb_98_14 gnd C_bl
Rb_98_15 bit_98_15 bit_98_16 R_bl
Rbb_98_15 bitb_98_15 bitb_98_16 R_bl
Cb_98_15 bit_98_15 gnd C_bl
Cbb_98_15 bitb_98_15 gnd C_bl
Rb_98_16 bit_98_16 bit_98_17 R_bl
Rbb_98_16 bitb_98_16 bitb_98_17 R_bl
Cb_98_16 bit_98_16 gnd C_bl
Cbb_98_16 bitb_98_16 gnd C_bl
Rb_98_17 bit_98_17 bit_98_18 R_bl
Rbb_98_17 bitb_98_17 bitb_98_18 R_bl
Cb_98_17 bit_98_17 gnd C_bl
Cbb_98_17 bitb_98_17 gnd C_bl
Rb_98_18 bit_98_18 bit_98_19 R_bl
Rbb_98_18 bitb_98_18 bitb_98_19 R_bl
Cb_98_18 bit_98_18 gnd C_bl
Cbb_98_18 bitb_98_18 gnd C_bl
Rb_98_19 bit_98_19 bit_98_20 R_bl
Rbb_98_19 bitb_98_19 bitb_98_20 R_bl
Cb_98_19 bit_98_19 gnd C_bl
Cbb_98_19 bitb_98_19 gnd C_bl
Rb_98_20 bit_98_20 bit_98_21 R_bl
Rbb_98_20 bitb_98_20 bitb_98_21 R_bl
Cb_98_20 bit_98_20 gnd C_bl
Cbb_98_20 bitb_98_20 gnd C_bl
Rb_98_21 bit_98_21 bit_98_22 R_bl
Rbb_98_21 bitb_98_21 bitb_98_22 R_bl
Cb_98_21 bit_98_21 gnd C_bl
Cbb_98_21 bitb_98_21 gnd C_bl
Rb_98_22 bit_98_22 bit_98_23 R_bl
Rbb_98_22 bitb_98_22 bitb_98_23 R_bl
Cb_98_22 bit_98_22 gnd C_bl
Cbb_98_22 bitb_98_22 gnd C_bl
Rb_98_23 bit_98_23 bit_98_24 R_bl
Rbb_98_23 bitb_98_23 bitb_98_24 R_bl
Cb_98_23 bit_98_23 gnd C_bl
Cbb_98_23 bitb_98_23 gnd C_bl
Rb_98_24 bit_98_24 bit_98_25 R_bl
Rbb_98_24 bitb_98_24 bitb_98_25 R_bl
Cb_98_24 bit_98_24 gnd C_bl
Cbb_98_24 bitb_98_24 gnd C_bl
Rb_98_25 bit_98_25 bit_98_26 R_bl
Rbb_98_25 bitb_98_25 bitb_98_26 R_bl
Cb_98_25 bit_98_25 gnd C_bl
Cbb_98_25 bitb_98_25 gnd C_bl
Rb_98_26 bit_98_26 bit_98_27 R_bl
Rbb_98_26 bitb_98_26 bitb_98_27 R_bl
Cb_98_26 bit_98_26 gnd C_bl
Cbb_98_26 bitb_98_26 gnd C_bl
Rb_98_27 bit_98_27 bit_98_28 R_bl
Rbb_98_27 bitb_98_27 bitb_98_28 R_bl
Cb_98_27 bit_98_27 gnd C_bl
Cbb_98_27 bitb_98_27 gnd C_bl
Rb_98_28 bit_98_28 bit_98_29 R_bl
Rbb_98_28 bitb_98_28 bitb_98_29 R_bl
Cb_98_28 bit_98_28 gnd C_bl
Cbb_98_28 bitb_98_28 gnd C_bl
Rb_98_29 bit_98_29 bit_98_30 R_bl
Rbb_98_29 bitb_98_29 bitb_98_30 R_bl
Cb_98_29 bit_98_29 gnd C_bl
Cbb_98_29 bitb_98_29 gnd C_bl
Rb_98_30 bit_98_30 bit_98_31 R_bl
Rbb_98_30 bitb_98_30 bitb_98_31 R_bl
Cb_98_30 bit_98_30 gnd C_bl
Cbb_98_30 bitb_98_30 gnd C_bl
Rb_98_31 bit_98_31 bit_98_32 R_bl
Rbb_98_31 bitb_98_31 bitb_98_32 R_bl
Cb_98_31 bit_98_31 gnd C_bl
Cbb_98_31 bitb_98_31 gnd C_bl
Rb_98_32 bit_98_32 bit_98_33 R_bl
Rbb_98_32 bitb_98_32 bitb_98_33 R_bl
Cb_98_32 bit_98_32 gnd C_bl
Cbb_98_32 bitb_98_32 gnd C_bl
Rb_98_33 bit_98_33 bit_98_34 R_bl
Rbb_98_33 bitb_98_33 bitb_98_34 R_bl
Cb_98_33 bit_98_33 gnd C_bl
Cbb_98_33 bitb_98_33 gnd C_bl
Rb_98_34 bit_98_34 bit_98_35 R_bl
Rbb_98_34 bitb_98_34 bitb_98_35 R_bl
Cb_98_34 bit_98_34 gnd C_bl
Cbb_98_34 bitb_98_34 gnd C_bl
Rb_98_35 bit_98_35 bit_98_36 R_bl
Rbb_98_35 bitb_98_35 bitb_98_36 R_bl
Cb_98_35 bit_98_35 gnd C_bl
Cbb_98_35 bitb_98_35 gnd C_bl
Rb_98_36 bit_98_36 bit_98_37 R_bl
Rbb_98_36 bitb_98_36 bitb_98_37 R_bl
Cb_98_36 bit_98_36 gnd C_bl
Cbb_98_36 bitb_98_36 gnd C_bl
Rb_98_37 bit_98_37 bit_98_38 R_bl
Rbb_98_37 bitb_98_37 bitb_98_38 R_bl
Cb_98_37 bit_98_37 gnd C_bl
Cbb_98_37 bitb_98_37 gnd C_bl
Rb_98_38 bit_98_38 bit_98_39 R_bl
Rbb_98_38 bitb_98_38 bitb_98_39 R_bl
Cb_98_38 bit_98_38 gnd C_bl
Cbb_98_38 bitb_98_38 gnd C_bl
Rb_98_39 bit_98_39 bit_98_40 R_bl
Rbb_98_39 bitb_98_39 bitb_98_40 R_bl
Cb_98_39 bit_98_39 gnd C_bl
Cbb_98_39 bitb_98_39 gnd C_bl
Rb_98_40 bit_98_40 bit_98_41 R_bl
Rbb_98_40 bitb_98_40 bitb_98_41 R_bl
Cb_98_40 bit_98_40 gnd C_bl
Cbb_98_40 bitb_98_40 gnd C_bl
Rb_98_41 bit_98_41 bit_98_42 R_bl
Rbb_98_41 bitb_98_41 bitb_98_42 R_bl
Cb_98_41 bit_98_41 gnd C_bl
Cbb_98_41 bitb_98_41 gnd C_bl
Rb_98_42 bit_98_42 bit_98_43 R_bl
Rbb_98_42 bitb_98_42 bitb_98_43 R_bl
Cb_98_42 bit_98_42 gnd C_bl
Cbb_98_42 bitb_98_42 gnd C_bl
Rb_98_43 bit_98_43 bit_98_44 R_bl
Rbb_98_43 bitb_98_43 bitb_98_44 R_bl
Cb_98_43 bit_98_43 gnd C_bl
Cbb_98_43 bitb_98_43 gnd C_bl
Rb_98_44 bit_98_44 bit_98_45 R_bl
Rbb_98_44 bitb_98_44 bitb_98_45 R_bl
Cb_98_44 bit_98_44 gnd C_bl
Cbb_98_44 bitb_98_44 gnd C_bl
Rb_98_45 bit_98_45 bit_98_46 R_bl
Rbb_98_45 bitb_98_45 bitb_98_46 R_bl
Cb_98_45 bit_98_45 gnd C_bl
Cbb_98_45 bitb_98_45 gnd C_bl
Rb_98_46 bit_98_46 bit_98_47 R_bl
Rbb_98_46 bitb_98_46 bitb_98_47 R_bl
Cb_98_46 bit_98_46 gnd C_bl
Cbb_98_46 bitb_98_46 gnd C_bl
Rb_98_47 bit_98_47 bit_98_48 R_bl
Rbb_98_47 bitb_98_47 bitb_98_48 R_bl
Cb_98_47 bit_98_47 gnd C_bl
Cbb_98_47 bitb_98_47 gnd C_bl
Rb_98_48 bit_98_48 bit_98_49 R_bl
Rbb_98_48 bitb_98_48 bitb_98_49 R_bl
Cb_98_48 bit_98_48 gnd C_bl
Cbb_98_48 bitb_98_48 gnd C_bl
Rb_98_49 bit_98_49 bit_98_50 R_bl
Rbb_98_49 bitb_98_49 bitb_98_50 R_bl
Cb_98_49 bit_98_49 gnd C_bl
Cbb_98_49 bitb_98_49 gnd C_bl
Rb_98_50 bit_98_50 bit_98_51 R_bl
Rbb_98_50 bitb_98_50 bitb_98_51 R_bl
Cb_98_50 bit_98_50 gnd C_bl
Cbb_98_50 bitb_98_50 gnd C_bl
Rb_98_51 bit_98_51 bit_98_52 R_bl
Rbb_98_51 bitb_98_51 bitb_98_52 R_bl
Cb_98_51 bit_98_51 gnd C_bl
Cbb_98_51 bitb_98_51 gnd C_bl
Rb_98_52 bit_98_52 bit_98_53 R_bl
Rbb_98_52 bitb_98_52 bitb_98_53 R_bl
Cb_98_52 bit_98_52 gnd C_bl
Cbb_98_52 bitb_98_52 gnd C_bl
Rb_98_53 bit_98_53 bit_98_54 R_bl
Rbb_98_53 bitb_98_53 bitb_98_54 R_bl
Cb_98_53 bit_98_53 gnd C_bl
Cbb_98_53 bitb_98_53 gnd C_bl
Rb_98_54 bit_98_54 bit_98_55 R_bl
Rbb_98_54 bitb_98_54 bitb_98_55 R_bl
Cb_98_54 bit_98_54 gnd C_bl
Cbb_98_54 bitb_98_54 gnd C_bl
Rb_98_55 bit_98_55 bit_98_56 R_bl
Rbb_98_55 bitb_98_55 bitb_98_56 R_bl
Cb_98_55 bit_98_55 gnd C_bl
Cbb_98_55 bitb_98_55 gnd C_bl
Rb_98_56 bit_98_56 bit_98_57 R_bl
Rbb_98_56 bitb_98_56 bitb_98_57 R_bl
Cb_98_56 bit_98_56 gnd C_bl
Cbb_98_56 bitb_98_56 gnd C_bl
Rb_98_57 bit_98_57 bit_98_58 R_bl
Rbb_98_57 bitb_98_57 bitb_98_58 R_bl
Cb_98_57 bit_98_57 gnd C_bl
Cbb_98_57 bitb_98_57 gnd C_bl
Rb_98_58 bit_98_58 bit_98_59 R_bl
Rbb_98_58 bitb_98_58 bitb_98_59 R_bl
Cb_98_58 bit_98_58 gnd C_bl
Cbb_98_58 bitb_98_58 gnd C_bl
Rb_98_59 bit_98_59 bit_98_60 R_bl
Rbb_98_59 bitb_98_59 bitb_98_60 R_bl
Cb_98_59 bit_98_59 gnd C_bl
Cbb_98_59 bitb_98_59 gnd C_bl
Rb_98_60 bit_98_60 bit_98_61 R_bl
Rbb_98_60 bitb_98_60 bitb_98_61 R_bl
Cb_98_60 bit_98_60 gnd C_bl
Cbb_98_60 bitb_98_60 gnd C_bl
Rb_98_61 bit_98_61 bit_98_62 R_bl
Rbb_98_61 bitb_98_61 bitb_98_62 R_bl
Cb_98_61 bit_98_61 gnd C_bl
Cbb_98_61 bitb_98_61 gnd C_bl
Rb_98_62 bit_98_62 bit_98_63 R_bl
Rbb_98_62 bitb_98_62 bitb_98_63 R_bl
Cb_98_62 bit_98_62 gnd C_bl
Cbb_98_62 bitb_98_62 gnd C_bl
Rb_98_63 bit_98_63 bit_98_64 R_bl
Rbb_98_63 bitb_98_63 bitb_98_64 R_bl
Cb_98_63 bit_98_63 gnd C_bl
Cbb_98_63 bitb_98_63 gnd C_bl
Rb_98_64 bit_98_64 bit_98_65 R_bl
Rbb_98_64 bitb_98_64 bitb_98_65 R_bl
Cb_98_64 bit_98_64 gnd C_bl
Cbb_98_64 bitb_98_64 gnd C_bl
Rb_98_65 bit_98_65 bit_98_66 R_bl
Rbb_98_65 bitb_98_65 bitb_98_66 R_bl
Cb_98_65 bit_98_65 gnd C_bl
Cbb_98_65 bitb_98_65 gnd C_bl
Rb_98_66 bit_98_66 bit_98_67 R_bl
Rbb_98_66 bitb_98_66 bitb_98_67 R_bl
Cb_98_66 bit_98_66 gnd C_bl
Cbb_98_66 bitb_98_66 gnd C_bl
Rb_98_67 bit_98_67 bit_98_68 R_bl
Rbb_98_67 bitb_98_67 bitb_98_68 R_bl
Cb_98_67 bit_98_67 gnd C_bl
Cbb_98_67 bitb_98_67 gnd C_bl
Rb_98_68 bit_98_68 bit_98_69 R_bl
Rbb_98_68 bitb_98_68 bitb_98_69 R_bl
Cb_98_68 bit_98_68 gnd C_bl
Cbb_98_68 bitb_98_68 gnd C_bl
Rb_98_69 bit_98_69 bit_98_70 R_bl
Rbb_98_69 bitb_98_69 bitb_98_70 R_bl
Cb_98_69 bit_98_69 gnd C_bl
Cbb_98_69 bitb_98_69 gnd C_bl
Rb_98_70 bit_98_70 bit_98_71 R_bl
Rbb_98_70 bitb_98_70 bitb_98_71 R_bl
Cb_98_70 bit_98_70 gnd C_bl
Cbb_98_70 bitb_98_70 gnd C_bl
Rb_98_71 bit_98_71 bit_98_72 R_bl
Rbb_98_71 bitb_98_71 bitb_98_72 R_bl
Cb_98_71 bit_98_71 gnd C_bl
Cbb_98_71 bitb_98_71 gnd C_bl
Rb_98_72 bit_98_72 bit_98_73 R_bl
Rbb_98_72 bitb_98_72 bitb_98_73 R_bl
Cb_98_72 bit_98_72 gnd C_bl
Cbb_98_72 bitb_98_72 gnd C_bl
Rb_98_73 bit_98_73 bit_98_74 R_bl
Rbb_98_73 bitb_98_73 bitb_98_74 R_bl
Cb_98_73 bit_98_73 gnd C_bl
Cbb_98_73 bitb_98_73 gnd C_bl
Rb_98_74 bit_98_74 bit_98_75 R_bl
Rbb_98_74 bitb_98_74 bitb_98_75 R_bl
Cb_98_74 bit_98_74 gnd C_bl
Cbb_98_74 bitb_98_74 gnd C_bl
Rb_98_75 bit_98_75 bit_98_76 R_bl
Rbb_98_75 bitb_98_75 bitb_98_76 R_bl
Cb_98_75 bit_98_75 gnd C_bl
Cbb_98_75 bitb_98_75 gnd C_bl
Rb_98_76 bit_98_76 bit_98_77 R_bl
Rbb_98_76 bitb_98_76 bitb_98_77 R_bl
Cb_98_76 bit_98_76 gnd C_bl
Cbb_98_76 bitb_98_76 gnd C_bl
Rb_98_77 bit_98_77 bit_98_78 R_bl
Rbb_98_77 bitb_98_77 bitb_98_78 R_bl
Cb_98_77 bit_98_77 gnd C_bl
Cbb_98_77 bitb_98_77 gnd C_bl
Rb_98_78 bit_98_78 bit_98_79 R_bl
Rbb_98_78 bitb_98_78 bitb_98_79 R_bl
Cb_98_78 bit_98_78 gnd C_bl
Cbb_98_78 bitb_98_78 gnd C_bl
Rb_98_79 bit_98_79 bit_98_80 R_bl
Rbb_98_79 bitb_98_79 bitb_98_80 R_bl
Cb_98_79 bit_98_79 gnd C_bl
Cbb_98_79 bitb_98_79 gnd C_bl
Rb_98_80 bit_98_80 bit_98_81 R_bl
Rbb_98_80 bitb_98_80 bitb_98_81 R_bl
Cb_98_80 bit_98_80 gnd C_bl
Cbb_98_80 bitb_98_80 gnd C_bl
Rb_98_81 bit_98_81 bit_98_82 R_bl
Rbb_98_81 bitb_98_81 bitb_98_82 R_bl
Cb_98_81 bit_98_81 gnd C_bl
Cbb_98_81 bitb_98_81 gnd C_bl
Rb_98_82 bit_98_82 bit_98_83 R_bl
Rbb_98_82 bitb_98_82 bitb_98_83 R_bl
Cb_98_82 bit_98_82 gnd C_bl
Cbb_98_82 bitb_98_82 gnd C_bl
Rb_98_83 bit_98_83 bit_98_84 R_bl
Rbb_98_83 bitb_98_83 bitb_98_84 R_bl
Cb_98_83 bit_98_83 gnd C_bl
Cbb_98_83 bitb_98_83 gnd C_bl
Rb_98_84 bit_98_84 bit_98_85 R_bl
Rbb_98_84 bitb_98_84 bitb_98_85 R_bl
Cb_98_84 bit_98_84 gnd C_bl
Cbb_98_84 bitb_98_84 gnd C_bl
Rb_98_85 bit_98_85 bit_98_86 R_bl
Rbb_98_85 bitb_98_85 bitb_98_86 R_bl
Cb_98_85 bit_98_85 gnd C_bl
Cbb_98_85 bitb_98_85 gnd C_bl
Rb_98_86 bit_98_86 bit_98_87 R_bl
Rbb_98_86 bitb_98_86 bitb_98_87 R_bl
Cb_98_86 bit_98_86 gnd C_bl
Cbb_98_86 bitb_98_86 gnd C_bl
Rb_98_87 bit_98_87 bit_98_88 R_bl
Rbb_98_87 bitb_98_87 bitb_98_88 R_bl
Cb_98_87 bit_98_87 gnd C_bl
Cbb_98_87 bitb_98_87 gnd C_bl
Rb_98_88 bit_98_88 bit_98_89 R_bl
Rbb_98_88 bitb_98_88 bitb_98_89 R_bl
Cb_98_88 bit_98_88 gnd C_bl
Cbb_98_88 bitb_98_88 gnd C_bl
Rb_98_89 bit_98_89 bit_98_90 R_bl
Rbb_98_89 bitb_98_89 bitb_98_90 R_bl
Cb_98_89 bit_98_89 gnd C_bl
Cbb_98_89 bitb_98_89 gnd C_bl
Rb_98_90 bit_98_90 bit_98_91 R_bl
Rbb_98_90 bitb_98_90 bitb_98_91 R_bl
Cb_98_90 bit_98_90 gnd C_bl
Cbb_98_90 bitb_98_90 gnd C_bl
Rb_98_91 bit_98_91 bit_98_92 R_bl
Rbb_98_91 bitb_98_91 bitb_98_92 R_bl
Cb_98_91 bit_98_91 gnd C_bl
Cbb_98_91 bitb_98_91 gnd C_bl
Rb_98_92 bit_98_92 bit_98_93 R_bl
Rbb_98_92 bitb_98_92 bitb_98_93 R_bl
Cb_98_92 bit_98_92 gnd C_bl
Cbb_98_92 bitb_98_92 gnd C_bl
Rb_98_93 bit_98_93 bit_98_94 R_bl
Rbb_98_93 bitb_98_93 bitb_98_94 R_bl
Cb_98_93 bit_98_93 gnd C_bl
Cbb_98_93 bitb_98_93 gnd C_bl
Rb_98_94 bit_98_94 bit_98_95 R_bl
Rbb_98_94 bitb_98_94 bitb_98_95 R_bl
Cb_98_94 bit_98_94 gnd C_bl
Cbb_98_94 bitb_98_94 gnd C_bl
Rb_98_95 bit_98_95 bit_98_96 R_bl
Rbb_98_95 bitb_98_95 bitb_98_96 R_bl
Cb_98_95 bit_98_95 gnd C_bl
Cbb_98_95 bitb_98_95 gnd C_bl
Rb_98_96 bit_98_96 bit_98_97 R_bl
Rbb_98_96 bitb_98_96 bitb_98_97 R_bl
Cb_98_96 bit_98_96 gnd C_bl
Cbb_98_96 bitb_98_96 gnd C_bl
Rb_98_97 bit_98_97 bit_98_98 R_bl
Rbb_98_97 bitb_98_97 bitb_98_98 R_bl
Cb_98_97 bit_98_97 gnd C_bl
Cbb_98_97 bitb_98_97 gnd C_bl
Rb_98_98 bit_98_98 bit_98_99 R_bl
Rbb_98_98 bitb_98_98 bitb_98_99 R_bl
Cb_98_98 bit_98_98 gnd C_bl
Cbb_98_98 bitb_98_98 gnd C_bl
Rb_98_99 bit_98_99 bit_98_100 R_bl
Rbb_98_99 bitb_98_99 bitb_98_100 R_bl
Cb_98_99 bit_98_99 gnd C_bl
Cbb_98_99 bitb_98_99 gnd C_bl
Rb_99_0 bit_99_0 bit_99_1 R_bl
Rbb_99_0 bitb_99_0 bitb_99_1 R_bl
Cb_99_0 bit_99_0 gnd C_bl
Cbb_99_0 bitb_99_0 gnd C_bl
Rb_99_1 bit_99_1 bit_99_2 R_bl
Rbb_99_1 bitb_99_1 bitb_99_2 R_bl
Cb_99_1 bit_99_1 gnd C_bl
Cbb_99_1 bitb_99_1 gnd C_bl
Rb_99_2 bit_99_2 bit_99_3 R_bl
Rbb_99_2 bitb_99_2 bitb_99_3 R_bl
Cb_99_2 bit_99_2 gnd C_bl
Cbb_99_2 bitb_99_2 gnd C_bl
Rb_99_3 bit_99_3 bit_99_4 R_bl
Rbb_99_3 bitb_99_3 bitb_99_4 R_bl
Cb_99_3 bit_99_3 gnd C_bl
Cbb_99_3 bitb_99_3 gnd C_bl
Rb_99_4 bit_99_4 bit_99_5 R_bl
Rbb_99_4 bitb_99_4 bitb_99_5 R_bl
Cb_99_4 bit_99_4 gnd C_bl
Cbb_99_4 bitb_99_4 gnd C_bl
Rb_99_5 bit_99_5 bit_99_6 R_bl
Rbb_99_5 bitb_99_5 bitb_99_6 R_bl
Cb_99_5 bit_99_5 gnd C_bl
Cbb_99_5 bitb_99_5 gnd C_bl
Rb_99_6 bit_99_6 bit_99_7 R_bl
Rbb_99_6 bitb_99_6 bitb_99_7 R_bl
Cb_99_6 bit_99_6 gnd C_bl
Cbb_99_6 bitb_99_6 gnd C_bl
Rb_99_7 bit_99_7 bit_99_8 R_bl
Rbb_99_7 bitb_99_7 bitb_99_8 R_bl
Cb_99_7 bit_99_7 gnd C_bl
Cbb_99_7 bitb_99_7 gnd C_bl
Rb_99_8 bit_99_8 bit_99_9 R_bl
Rbb_99_8 bitb_99_8 bitb_99_9 R_bl
Cb_99_8 bit_99_8 gnd C_bl
Cbb_99_8 bitb_99_8 gnd C_bl
Rb_99_9 bit_99_9 bit_99_10 R_bl
Rbb_99_9 bitb_99_9 bitb_99_10 R_bl
Cb_99_9 bit_99_9 gnd C_bl
Cbb_99_9 bitb_99_9 gnd C_bl
Rb_99_10 bit_99_10 bit_99_11 R_bl
Rbb_99_10 bitb_99_10 bitb_99_11 R_bl
Cb_99_10 bit_99_10 gnd C_bl
Cbb_99_10 bitb_99_10 gnd C_bl
Rb_99_11 bit_99_11 bit_99_12 R_bl
Rbb_99_11 bitb_99_11 bitb_99_12 R_bl
Cb_99_11 bit_99_11 gnd C_bl
Cbb_99_11 bitb_99_11 gnd C_bl
Rb_99_12 bit_99_12 bit_99_13 R_bl
Rbb_99_12 bitb_99_12 bitb_99_13 R_bl
Cb_99_12 bit_99_12 gnd C_bl
Cbb_99_12 bitb_99_12 gnd C_bl
Rb_99_13 bit_99_13 bit_99_14 R_bl
Rbb_99_13 bitb_99_13 bitb_99_14 R_bl
Cb_99_13 bit_99_13 gnd C_bl
Cbb_99_13 bitb_99_13 gnd C_bl
Rb_99_14 bit_99_14 bit_99_15 R_bl
Rbb_99_14 bitb_99_14 bitb_99_15 R_bl
Cb_99_14 bit_99_14 gnd C_bl
Cbb_99_14 bitb_99_14 gnd C_bl
Rb_99_15 bit_99_15 bit_99_16 R_bl
Rbb_99_15 bitb_99_15 bitb_99_16 R_bl
Cb_99_15 bit_99_15 gnd C_bl
Cbb_99_15 bitb_99_15 gnd C_bl
Rb_99_16 bit_99_16 bit_99_17 R_bl
Rbb_99_16 bitb_99_16 bitb_99_17 R_bl
Cb_99_16 bit_99_16 gnd C_bl
Cbb_99_16 bitb_99_16 gnd C_bl
Rb_99_17 bit_99_17 bit_99_18 R_bl
Rbb_99_17 bitb_99_17 bitb_99_18 R_bl
Cb_99_17 bit_99_17 gnd C_bl
Cbb_99_17 bitb_99_17 gnd C_bl
Rb_99_18 bit_99_18 bit_99_19 R_bl
Rbb_99_18 bitb_99_18 bitb_99_19 R_bl
Cb_99_18 bit_99_18 gnd C_bl
Cbb_99_18 bitb_99_18 gnd C_bl
Rb_99_19 bit_99_19 bit_99_20 R_bl
Rbb_99_19 bitb_99_19 bitb_99_20 R_bl
Cb_99_19 bit_99_19 gnd C_bl
Cbb_99_19 bitb_99_19 gnd C_bl
Rb_99_20 bit_99_20 bit_99_21 R_bl
Rbb_99_20 bitb_99_20 bitb_99_21 R_bl
Cb_99_20 bit_99_20 gnd C_bl
Cbb_99_20 bitb_99_20 gnd C_bl
Rb_99_21 bit_99_21 bit_99_22 R_bl
Rbb_99_21 bitb_99_21 bitb_99_22 R_bl
Cb_99_21 bit_99_21 gnd C_bl
Cbb_99_21 bitb_99_21 gnd C_bl
Rb_99_22 bit_99_22 bit_99_23 R_bl
Rbb_99_22 bitb_99_22 bitb_99_23 R_bl
Cb_99_22 bit_99_22 gnd C_bl
Cbb_99_22 bitb_99_22 gnd C_bl
Rb_99_23 bit_99_23 bit_99_24 R_bl
Rbb_99_23 bitb_99_23 bitb_99_24 R_bl
Cb_99_23 bit_99_23 gnd C_bl
Cbb_99_23 bitb_99_23 gnd C_bl
Rb_99_24 bit_99_24 bit_99_25 R_bl
Rbb_99_24 bitb_99_24 bitb_99_25 R_bl
Cb_99_24 bit_99_24 gnd C_bl
Cbb_99_24 bitb_99_24 gnd C_bl
Rb_99_25 bit_99_25 bit_99_26 R_bl
Rbb_99_25 bitb_99_25 bitb_99_26 R_bl
Cb_99_25 bit_99_25 gnd C_bl
Cbb_99_25 bitb_99_25 gnd C_bl
Rb_99_26 bit_99_26 bit_99_27 R_bl
Rbb_99_26 bitb_99_26 bitb_99_27 R_bl
Cb_99_26 bit_99_26 gnd C_bl
Cbb_99_26 bitb_99_26 gnd C_bl
Rb_99_27 bit_99_27 bit_99_28 R_bl
Rbb_99_27 bitb_99_27 bitb_99_28 R_bl
Cb_99_27 bit_99_27 gnd C_bl
Cbb_99_27 bitb_99_27 gnd C_bl
Rb_99_28 bit_99_28 bit_99_29 R_bl
Rbb_99_28 bitb_99_28 bitb_99_29 R_bl
Cb_99_28 bit_99_28 gnd C_bl
Cbb_99_28 bitb_99_28 gnd C_bl
Rb_99_29 bit_99_29 bit_99_30 R_bl
Rbb_99_29 bitb_99_29 bitb_99_30 R_bl
Cb_99_29 bit_99_29 gnd C_bl
Cbb_99_29 bitb_99_29 gnd C_bl
Rb_99_30 bit_99_30 bit_99_31 R_bl
Rbb_99_30 bitb_99_30 bitb_99_31 R_bl
Cb_99_30 bit_99_30 gnd C_bl
Cbb_99_30 bitb_99_30 gnd C_bl
Rb_99_31 bit_99_31 bit_99_32 R_bl
Rbb_99_31 bitb_99_31 bitb_99_32 R_bl
Cb_99_31 bit_99_31 gnd C_bl
Cbb_99_31 bitb_99_31 gnd C_bl
Rb_99_32 bit_99_32 bit_99_33 R_bl
Rbb_99_32 bitb_99_32 bitb_99_33 R_bl
Cb_99_32 bit_99_32 gnd C_bl
Cbb_99_32 bitb_99_32 gnd C_bl
Rb_99_33 bit_99_33 bit_99_34 R_bl
Rbb_99_33 bitb_99_33 bitb_99_34 R_bl
Cb_99_33 bit_99_33 gnd C_bl
Cbb_99_33 bitb_99_33 gnd C_bl
Rb_99_34 bit_99_34 bit_99_35 R_bl
Rbb_99_34 bitb_99_34 bitb_99_35 R_bl
Cb_99_34 bit_99_34 gnd C_bl
Cbb_99_34 bitb_99_34 gnd C_bl
Rb_99_35 bit_99_35 bit_99_36 R_bl
Rbb_99_35 bitb_99_35 bitb_99_36 R_bl
Cb_99_35 bit_99_35 gnd C_bl
Cbb_99_35 bitb_99_35 gnd C_bl
Rb_99_36 bit_99_36 bit_99_37 R_bl
Rbb_99_36 bitb_99_36 bitb_99_37 R_bl
Cb_99_36 bit_99_36 gnd C_bl
Cbb_99_36 bitb_99_36 gnd C_bl
Rb_99_37 bit_99_37 bit_99_38 R_bl
Rbb_99_37 bitb_99_37 bitb_99_38 R_bl
Cb_99_37 bit_99_37 gnd C_bl
Cbb_99_37 bitb_99_37 gnd C_bl
Rb_99_38 bit_99_38 bit_99_39 R_bl
Rbb_99_38 bitb_99_38 bitb_99_39 R_bl
Cb_99_38 bit_99_38 gnd C_bl
Cbb_99_38 bitb_99_38 gnd C_bl
Rb_99_39 bit_99_39 bit_99_40 R_bl
Rbb_99_39 bitb_99_39 bitb_99_40 R_bl
Cb_99_39 bit_99_39 gnd C_bl
Cbb_99_39 bitb_99_39 gnd C_bl
Rb_99_40 bit_99_40 bit_99_41 R_bl
Rbb_99_40 bitb_99_40 bitb_99_41 R_bl
Cb_99_40 bit_99_40 gnd C_bl
Cbb_99_40 bitb_99_40 gnd C_bl
Rb_99_41 bit_99_41 bit_99_42 R_bl
Rbb_99_41 bitb_99_41 bitb_99_42 R_bl
Cb_99_41 bit_99_41 gnd C_bl
Cbb_99_41 bitb_99_41 gnd C_bl
Rb_99_42 bit_99_42 bit_99_43 R_bl
Rbb_99_42 bitb_99_42 bitb_99_43 R_bl
Cb_99_42 bit_99_42 gnd C_bl
Cbb_99_42 bitb_99_42 gnd C_bl
Rb_99_43 bit_99_43 bit_99_44 R_bl
Rbb_99_43 bitb_99_43 bitb_99_44 R_bl
Cb_99_43 bit_99_43 gnd C_bl
Cbb_99_43 bitb_99_43 gnd C_bl
Rb_99_44 bit_99_44 bit_99_45 R_bl
Rbb_99_44 bitb_99_44 bitb_99_45 R_bl
Cb_99_44 bit_99_44 gnd C_bl
Cbb_99_44 bitb_99_44 gnd C_bl
Rb_99_45 bit_99_45 bit_99_46 R_bl
Rbb_99_45 bitb_99_45 bitb_99_46 R_bl
Cb_99_45 bit_99_45 gnd C_bl
Cbb_99_45 bitb_99_45 gnd C_bl
Rb_99_46 bit_99_46 bit_99_47 R_bl
Rbb_99_46 bitb_99_46 bitb_99_47 R_bl
Cb_99_46 bit_99_46 gnd C_bl
Cbb_99_46 bitb_99_46 gnd C_bl
Rb_99_47 bit_99_47 bit_99_48 R_bl
Rbb_99_47 bitb_99_47 bitb_99_48 R_bl
Cb_99_47 bit_99_47 gnd C_bl
Cbb_99_47 bitb_99_47 gnd C_bl
Rb_99_48 bit_99_48 bit_99_49 R_bl
Rbb_99_48 bitb_99_48 bitb_99_49 R_bl
Cb_99_48 bit_99_48 gnd C_bl
Cbb_99_48 bitb_99_48 gnd C_bl
Rb_99_49 bit_99_49 bit_99_50 R_bl
Rbb_99_49 bitb_99_49 bitb_99_50 R_bl
Cb_99_49 bit_99_49 gnd C_bl
Cbb_99_49 bitb_99_49 gnd C_bl
Rb_99_50 bit_99_50 bit_99_51 R_bl
Rbb_99_50 bitb_99_50 bitb_99_51 R_bl
Cb_99_50 bit_99_50 gnd C_bl
Cbb_99_50 bitb_99_50 gnd C_bl
Rb_99_51 bit_99_51 bit_99_52 R_bl
Rbb_99_51 bitb_99_51 bitb_99_52 R_bl
Cb_99_51 bit_99_51 gnd C_bl
Cbb_99_51 bitb_99_51 gnd C_bl
Rb_99_52 bit_99_52 bit_99_53 R_bl
Rbb_99_52 bitb_99_52 bitb_99_53 R_bl
Cb_99_52 bit_99_52 gnd C_bl
Cbb_99_52 bitb_99_52 gnd C_bl
Rb_99_53 bit_99_53 bit_99_54 R_bl
Rbb_99_53 bitb_99_53 bitb_99_54 R_bl
Cb_99_53 bit_99_53 gnd C_bl
Cbb_99_53 bitb_99_53 gnd C_bl
Rb_99_54 bit_99_54 bit_99_55 R_bl
Rbb_99_54 bitb_99_54 bitb_99_55 R_bl
Cb_99_54 bit_99_54 gnd C_bl
Cbb_99_54 bitb_99_54 gnd C_bl
Rb_99_55 bit_99_55 bit_99_56 R_bl
Rbb_99_55 bitb_99_55 bitb_99_56 R_bl
Cb_99_55 bit_99_55 gnd C_bl
Cbb_99_55 bitb_99_55 gnd C_bl
Rb_99_56 bit_99_56 bit_99_57 R_bl
Rbb_99_56 bitb_99_56 bitb_99_57 R_bl
Cb_99_56 bit_99_56 gnd C_bl
Cbb_99_56 bitb_99_56 gnd C_bl
Rb_99_57 bit_99_57 bit_99_58 R_bl
Rbb_99_57 bitb_99_57 bitb_99_58 R_bl
Cb_99_57 bit_99_57 gnd C_bl
Cbb_99_57 bitb_99_57 gnd C_bl
Rb_99_58 bit_99_58 bit_99_59 R_bl
Rbb_99_58 bitb_99_58 bitb_99_59 R_bl
Cb_99_58 bit_99_58 gnd C_bl
Cbb_99_58 bitb_99_58 gnd C_bl
Rb_99_59 bit_99_59 bit_99_60 R_bl
Rbb_99_59 bitb_99_59 bitb_99_60 R_bl
Cb_99_59 bit_99_59 gnd C_bl
Cbb_99_59 bitb_99_59 gnd C_bl
Rb_99_60 bit_99_60 bit_99_61 R_bl
Rbb_99_60 bitb_99_60 bitb_99_61 R_bl
Cb_99_60 bit_99_60 gnd C_bl
Cbb_99_60 bitb_99_60 gnd C_bl
Rb_99_61 bit_99_61 bit_99_62 R_bl
Rbb_99_61 bitb_99_61 bitb_99_62 R_bl
Cb_99_61 bit_99_61 gnd C_bl
Cbb_99_61 bitb_99_61 gnd C_bl
Rb_99_62 bit_99_62 bit_99_63 R_bl
Rbb_99_62 bitb_99_62 bitb_99_63 R_bl
Cb_99_62 bit_99_62 gnd C_bl
Cbb_99_62 bitb_99_62 gnd C_bl
Rb_99_63 bit_99_63 bit_99_64 R_bl
Rbb_99_63 bitb_99_63 bitb_99_64 R_bl
Cb_99_63 bit_99_63 gnd C_bl
Cbb_99_63 bitb_99_63 gnd C_bl
Rb_99_64 bit_99_64 bit_99_65 R_bl
Rbb_99_64 bitb_99_64 bitb_99_65 R_bl
Cb_99_64 bit_99_64 gnd C_bl
Cbb_99_64 bitb_99_64 gnd C_bl
Rb_99_65 bit_99_65 bit_99_66 R_bl
Rbb_99_65 bitb_99_65 bitb_99_66 R_bl
Cb_99_65 bit_99_65 gnd C_bl
Cbb_99_65 bitb_99_65 gnd C_bl
Rb_99_66 bit_99_66 bit_99_67 R_bl
Rbb_99_66 bitb_99_66 bitb_99_67 R_bl
Cb_99_66 bit_99_66 gnd C_bl
Cbb_99_66 bitb_99_66 gnd C_bl
Rb_99_67 bit_99_67 bit_99_68 R_bl
Rbb_99_67 bitb_99_67 bitb_99_68 R_bl
Cb_99_67 bit_99_67 gnd C_bl
Cbb_99_67 bitb_99_67 gnd C_bl
Rb_99_68 bit_99_68 bit_99_69 R_bl
Rbb_99_68 bitb_99_68 bitb_99_69 R_bl
Cb_99_68 bit_99_68 gnd C_bl
Cbb_99_68 bitb_99_68 gnd C_bl
Rb_99_69 bit_99_69 bit_99_70 R_bl
Rbb_99_69 bitb_99_69 bitb_99_70 R_bl
Cb_99_69 bit_99_69 gnd C_bl
Cbb_99_69 bitb_99_69 gnd C_bl
Rb_99_70 bit_99_70 bit_99_71 R_bl
Rbb_99_70 bitb_99_70 bitb_99_71 R_bl
Cb_99_70 bit_99_70 gnd C_bl
Cbb_99_70 bitb_99_70 gnd C_bl
Rb_99_71 bit_99_71 bit_99_72 R_bl
Rbb_99_71 bitb_99_71 bitb_99_72 R_bl
Cb_99_71 bit_99_71 gnd C_bl
Cbb_99_71 bitb_99_71 gnd C_bl
Rb_99_72 bit_99_72 bit_99_73 R_bl
Rbb_99_72 bitb_99_72 bitb_99_73 R_bl
Cb_99_72 bit_99_72 gnd C_bl
Cbb_99_72 bitb_99_72 gnd C_bl
Rb_99_73 bit_99_73 bit_99_74 R_bl
Rbb_99_73 bitb_99_73 bitb_99_74 R_bl
Cb_99_73 bit_99_73 gnd C_bl
Cbb_99_73 bitb_99_73 gnd C_bl
Rb_99_74 bit_99_74 bit_99_75 R_bl
Rbb_99_74 bitb_99_74 bitb_99_75 R_bl
Cb_99_74 bit_99_74 gnd C_bl
Cbb_99_74 bitb_99_74 gnd C_bl
Rb_99_75 bit_99_75 bit_99_76 R_bl
Rbb_99_75 bitb_99_75 bitb_99_76 R_bl
Cb_99_75 bit_99_75 gnd C_bl
Cbb_99_75 bitb_99_75 gnd C_bl
Rb_99_76 bit_99_76 bit_99_77 R_bl
Rbb_99_76 bitb_99_76 bitb_99_77 R_bl
Cb_99_76 bit_99_76 gnd C_bl
Cbb_99_76 bitb_99_76 gnd C_bl
Rb_99_77 bit_99_77 bit_99_78 R_bl
Rbb_99_77 bitb_99_77 bitb_99_78 R_bl
Cb_99_77 bit_99_77 gnd C_bl
Cbb_99_77 bitb_99_77 gnd C_bl
Rb_99_78 bit_99_78 bit_99_79 R_bl
Rbb_99_78 bitb_99_78 bitb_99_79 R_bl
Cb_99_78 bit_99_78 gnd C_bl
Cbb_99_78 bitb_99_78 gnd C_bl
Rb_99_79 bit_99_79 bit_99_80 R_bl
Rbb_99_79 bitb_99_79 bitb_99_80 R_bl
Cb_99_79 bit_99_79 gnd C_bl
Cbb_99_79 bitb_99_79 gnd C_bl
Rb_99_80 bit_99_80 bit_99_81 R_bl
Rbb_99_80 bitb_99_80 bitb_99_81 R_bl
Cb_99_80 bit_99_80 gnd C_bl
Cbb_99_80 bitb_99_80 gnd C_bl
Rb_99_81 bit_99_81 bit_99_82 R_bl
Rbb_99_81 bitb_99_81 bitb_99_82 R_bl
Cb_99_81 bit_99_81 gnd C_bl
Cbb_99_81 bitb_99_81 gnd C_bl
Rb_99_82 bit_99_82 bit_99_83 R_bl
Rbb_99_82 bitb_99_82 bitb_99_83 R_bl
Cb_99_82 bit_99_82 gnd C_bl
Cbb_99_82 bitb_99_82 gnd C_bl
Rb_99_83 bit_99_83 bit_99_84 R_bl
Rbb_99_83 bitb_99_83 bitb_99_84 R_bl
Cb_99_83 bit_99_83 gnd C_bl
Cbb_99_83 bitb_99_83 gnd C_bl
Rb_99_84 bit_99_84 bit_99_85 R_bl
Rbb_99_84 bitb_99_84 bitb_99_85 R_bl
Cb_99_84 bit_99_84 gnd C_bl
Cbb_99_84 bitb_99_84 gnd C_bl
Rb_99_85 bit_99_85 bit_99_86 R_bl
Rbb_99_85 bitb_99_85 bitb_99_86 R_bl
Cb_99_85 bit_99_85 gnd C_bl
Cbb_99_85 bitb_99_85 gnd C_bl
Rb_99_86 bit_99_86 bit_99_87 R_bl
Rbb_99_86 bitb_99_86 bitb_99_87 R_bl
Cb_99_86 bit_99_86 gnd C_bl
Cbb_99_86 bitb_99_86 gnd C_bl
Rb_99_87 bit_99_87 bit_99_88 R_bl
Rbb_99_87 bitb_99_87 bitb_99_88 R_bl
Cb_99_87 bit_99_87 gnd C_bl
Cbb_99_87 bitb_99_87 gnd C_bl
Rb_99_88 bit_99_88 bit_99_89 R_bl
Rbb_99_88 bitb_99_88 bitb_99_89 R_bl
Cb_99_88 bit_99_88 gnd C_bl
Cbb_99_88 bitb_99_88 gnd C_bl
Rb_99_89 bit_99_89 bit_99_90 R_bl
Rbb_99_89 bitb_99_89 bitb_99_90 R_bl
Cb_99_89 bit_99_89 gnd C_bl
Cbb_99_89 bitb_99_89 gnd C_bl
Rb_99_90 bit_99_90 bit_99_91 R_bl
Rbb_99_90 bitb_99_90 bitb_99_91 R_bl
Cb_99_90 bit_99_90 gnd C_bl
Cbb_99_90 bitb_99_90 gnd C_bl
Rb_99_91 bit_99_91 bit_99_92 R_bl
Rbb_99_91 bitb_99_91 bitb_99_92 R_bl
Cb_99_91 bit_99_91 gnd C_bl
Cbb_99_91 bitb_99_91 gnd C_bl
Rb_99_92 bit_99_92 bit_99_93 R_bl
Rbb_99_92 bitb_99_92 bitb_99_93 R_bl
Cb_99_92 bit_99_92 gnd C_bl
Cbb_99_92 bitb_99_92 gnd C_bl
Rb_99_93 bit_99_93 bit_99_94 R_bl
Rbb_99_93 bitb_99_93 bitb_99_94 R_bl
Cb_99_93 bit_99_93 gnd C_bl
Cbb_99_93 bitb_99_93 gnd C_bl
Rb_99_94 bit_99_94 bit_99_95 R_bl
Rbb_99_94 bitb_99_94 bitb_99_95 R_bl
Cb_99_94 bit_99_94 gnd C_bl
Cbb_99_94 bitb_99_94 gnd C_bl
Rb_99_95 bit_99_95 bit_99_96 R_bl
Rbb_99_95 bitb_99_95 bitb_99_96 R_bl
Cb_99_95 bit_99_95 gnd C_bl
Cbb_99_95 bitb_99_95 gnd C_bl
Rb_99_96 bit_99_96 bit_99_97 R_bl
Rbb_99_96 bitb_99_96 bitb_99_97 R_bl
Cb_99_96 bit_99_96 gnd C_bl
Cbb_99_96 bitb_99_96 gnd C_bl
Rb_99_97 bit_99_97 bit_99_98 R_bl
Rbb_99_97 bitb_99_97 bitb_99_98 R_bl
Cb_99_97 bit_99_97 gnd C_bl
Cbb_99_97 bitb_99_97 gnd C_bl
Rb_99_98 bit_99_98 bit_99_99 R_bl
Rbb_99_98 bitb_99_98 bitb_99_99 R_bl
Cb_99_98 bit_99_98 gnd C_bl
Cbb_99_98 bitb_99_98 gnd C_bl
Rb_99_99 bit_99_99 bit_99_100 R_bl
Rbb_99_99 bitb_99_99 bitb_99_100 R_bl
Cb_99_99 bit_99_99 gnd C_bl
Cbb_99_99 bitb_99_99 gnd C_bl
Vwrite_0 write_0 gnd dc 0
Vwrite_1 write_1 gnd dc 0
Vwrite_2 write_2 gnd dc 0
Vwrite_3 write_3 gnd dc 0
Vwrite_4 write_4 gnd dc 0
Vwrite_5 write_5 gnd dc 0
Vwrite_6 write_6 gnd dc 0
Vwrite_7 write_7 gnd dc 0
Vwrite_8 write_8 gnd dc 0
Vwrite_9 write_9 gnd dc 0
Vwrite_10 write_10 gnd dc 0
Vwrite_11 write_11 gnd dc 0
Vwrite_12 write_12 gnd dc 0
Vwrite_13 write_13 gnd dc 0
Vwrite_14 write_14 gnd dc 0
Vwrite_15 write_15 gnd dc 0
Vwrite_16 write_16 gnd dc 0
Vwrite_17 write_17 gnd dc 0
Vwrite_18 write_18 gnd dc 0
Vwrite_19 write_19 gnd dc 0
Vwrite_20 write_20 gnd dc 0
Vwrite_21 write_21 gnd dc 0
Vwrite_22 write_22 gnd dc 0
Vwrite_23 write_23 gnd dc 0
Vwrite_24 write_24 gnd dc 0
Vwrite_25 write_25 gnd dc 0
Vwrite_26 write_26 gnd dc 0
Vwrite_27 write_27 gnd dc 0
Vwrite_28 write_28 gnd dc 0
Vwrite_29 write_29 gnd dc 0
Vwrite_30 write_30 gnd dc 0
Vwrite_31 write_31 gnd dc 0
Vwrite_32 write_32 gnd dc 0
Vwrite_33 write_33 gnd dc 0
Vwrite_34 write_34 gnd dc 0
Vwrite_35 write_35 gnd dc 0
Vwrite_36 write_36 gnd dc 0
Vwrite_37 write_37 gnd dc 0
Vwrite_38 write_38 gnd dc 0
Vwrite_39 write_39 gnd dc 0
Vwrite_40 write_40 gnd dc 0
Vwrite_41 write_41 gnd dc 0
Vwrite_42 write_42 gnd dc 0
Vwrite_43 write_43 gnd dc 0
Vwrite_44 write_44 gnd dc 0
Vwrite_45 write_45 gnd dc 0
Vwrite_46 write_46 gnd dc 0
Vwrite_47 write_47 gnd dc 0
Vwrite_48 write_48 gnd dc 0
Vwrite_49 write_49 gnd dc 0
Vwrite_50 write_50 gnd dc 0
Vwrite_51 write_51 gnd dc 0
Vwrite_52 write_52 gnd dc 0
Vwrite_53 write_53 gnd dc 0
Vwrite_54 write_54 gnd dc 0
Vwrite_55 write_55 gnd dc 0
Vwrite_56 write_56 gnd dc 0
Vwrite_57 write_57 gnd dc 0
Vwrite_58 write_58 gnd dc 0
Vwrite_59 write_59 gnd dc 0
Vwrite_60 write_60 gnd dc 0
Vwrite_61 write_61 gnd dc 0
Vwrite_62 write_62 gnd dc 0
Vwrite_63 write_63 gnd dc 0
Vwrite_64 write_64 gnd dc 0
Vwrite_65 write_65 gnd dc 0
Vwrite_66 write_66 gnd dc 0
Vwrite_67 write_67 gnd dc 0
Vwrite_68 write_68 gnd dc 0
Vwrite_69 write_69 gnd dc 0
Vwrite_70 write_70 gnd dc 0
Vwrite_71 write_71 gnd dc 0
Vwrite_72 write_72 gnd dc 0
Vwrite_73 write_73 gnd dc 0
Vwrite_74 write_74 gnd dc 0
Vwrite_75 write_75 gnd dc 0
Vwrite_76 write_76 gnd dc 0
Vwrite_77 write_77 gnd dc 0
Vwrite_78 write_78 gnd dc 0
Vwrite_79 write_79 gnd dc 0
Vwrite_80 write_80 gnd dc 0
Vwrite_81 write_81 gnd dc 0
Vwrite_82 write_82 gnd dc 0
Vwrite_83 write_83 gnd dc 0
Vwrite_84 write_84 gnd dc 0
Vwrite_85 write_85 gnd dc 0
Vwrite_86 write_86 gnd dc 0
Vwrite_87 write_87 gnd dc 0
Vwrite_88 write_88 gnd dc 0
Vwrite_89 write_89 gnd dc 0
Vwrite_90 write_90 gnd dc 0
Vwrite_91 write_91 gnd dc 0
Vwrite_92 write_92 gnd dc 0
Vwrite_93 write_93 gnd dc 0
Vwrite_94 write_94 gnd dc 0
Vwrite_95 write_95 gnd dc 0
Vwrite_96 write_96 gnd dc 0
Vwrite_97 write_97 gnd dc 0
Vwrite_98 write_98 gnd dc 0
Vwrite_99 write_99 gnd dc 0
Vdata_0 data_0 gnd dc 0 
Vdatab_0 datab_0 gnd dc 1.8
Vdata_1 data_1 gnd dc 0 
Vdatab_1 datab_1 gnd dc 1.8
Vdata_2 data_2 gnd dc 0 
Vdatab_2 datab_2 gnd dc 1.8
Vdata_3 data_3 gnd dc 0 
Vdatab_3 datab_3 gnd dc 1.8
Vdata_4 data_4 gnd dc 0 
Vdatab_4 datab_4 gnd dc 1.8
Vdata_5 data_5 gnd dc 0 
Vdatab_5 datab_5 gnd dc 1.8
Vdata_6 data_6 gnd dc 0 
Vdatab_6 datab_6 gnd dc 1.8
Vdata_7 data_7 gnd dc 0 
Vdatab_7 datab_7 gnd dc 1.8
Vdata_8 data_8 gnd dc 0 
Vdatab_8 datab_8 gnd dc 1.8
Vdata_9 data_9 gnd dc 0 
Vdatab_9 datab_9 gnd dc 1.8
Vdata_10 data_10 gnd dc 0 
Vdatab_10 datab_10 gnd dc 1.8
Vdata_11 data_11 gnd dc 0 
Vdatab_11 datab_11 gnd dc 1.8
Vdata_12 data_12 gnd dc 0 
Vdatab_12 datab_12 gnd dc 1.8
Vdata_13 data_13 gnd dc 0 
Vdatab_13 datab_13 gnd dc 1.8
Vdata_14 data_14 gnd dc 0 
Vdatab_14 datab_14 gnd dc 1.8
Vdata_15 data_15 gnd dc 0 
Vdatab_15 datab_15 gnd dc 1.8
Vdata_16 data_16 gnd dc 0 
Vdatab_16 datab_16 gnd dc 1.8
Vdata_17 data_17 gnd dc 0 
Vdatab_17 datab_17 gnd dc 1.8
Vdata_18 data_18 gnd dc 0 
Vdatab_18 datab_18 gnd dc 1.8
Vdata_19 data_19 gnd dc 0 
Vdatab_19 datab_19 gnd dc 1.8
Vdata_20 data_20 gnd dc 0 
Vdatab_20 datab_20 gnd dc 1.8
Vdata_21 data_21 gnd dc 0 
Vdatab_21 datab_21 gnd dc 1.8
Vdata_22 data_22 gnd dc 0 
Vdatab_22 datab_22 gnd dc 1.8
Vdata_23 data_23 gnd dc 0 
Vdatab_23 datab_23 gnd dc 1.8
Vdata_24 data_24 gnd dc 0 
Vdatab_24 datab_24 gnd dc 1.8
Vdata_25 data_25 gnd dc 0 
Vdatab_25 datab_25 gnd dc 1.8
Vdata_26 data_26 gnd dc 0 
Vdatab_26 datab_26 gnd dc 1.8
Vdata_27 data_27 gnd dc 0 
Vdatab_27 datab_27 gnd dc 1.8
Vdata_28 data_28 gnd dc 0 
Vdatab_28 datab_28 gnd dc 1.8
Vdata_29 data_29 gnd dc 0 
Vdatab_29 datab_29 gnd dc 1.8
Vdata_30 data_30 gnd dc 0 
Vdatab_30 datab_30 gnd dc 1.8
Vdata_31 data_31 gnd dc 0 
Vdatab_31 datab_31 gnd dc 1.8
Vdata_32 data_32 gnd dc 0 
Vdatab_32 datab_32 gnd dc 1.8
Vdata_33 data_33 gnd dc 0 
Vdatab_33 datab_33 gnd dc 1.8
Vdata_34 data_34 gnd dc 0 
Vdatab_34 datab_34 gnd dc 1.8
Vdata_35 data_35 gnd dc 0 
Vdatab_35 datab_35 gnd dc 1.8
Vdata_36 data_36 gnd dc 0 
Vdatab_36 datab_36 gnd dc 1.8
Vdata_37 data_37 gnd dc 0 
Vdatab_37 datab_37 gnd dc 1.8
Vdata_38 data_38 gnd dc 0 
Vdatab_38 datab_38 gnd dc 1.8
Vdata_39 data_39 gnd dc 0 
Vdatab_39 datab_39 gnd dc 1.8
Vdata_40 data_40 gnd dc 0 
Vdatab_40 datab_40 gnd dc 1.8
Vdata_41 data_41 gnd dc 0 
Vdatab_41 datab_41 gnd dc 1.8
Vdata_42 data_42 gnd dc 0 
Vdatab_42 datab_42 gnd dc 1.8
Vdata_43 data_43 gnd dc 0 
Vdatab_43 datab_43 gnd dc 1.8
Vdata_44 data_44 gnd dc 0 
Vdatab_44 datab_44 gnd dc 1.8
Vdata_45 data_45 gnd dc 0 
Vdatab_45 datab_45 gnd dc 1.8
Vdata_46 data_46 gnd dc 0 
Vdatab_46 datab_46 gnd dc 1.8
Vdata_47 data_47 gnd dc 0 
Vdatab_47 datab_47 gnd dc 1.8
Vdata_48 data_48 gnd dc 0 
Vdatab_48 datab_48 gnd dc 1.8
Vdata_49 data_49 gnd dc 0 
Vdatab_49 datab_49 gnd dc 1.8
Vdata_50 data_50 gnd dc 0 
Vdatab_50 datab_50 gnd dc 1.8
Vdata_51 data_51 gnd dc 0 
Vdatab_51 datab_51 gnd dc 1.8
Vdata_52 data_52 gnd dc 0 
Vdatab_52 datab_52 gnd dc 1.8
Vdata_53 data_53 gnd dc 0 
Vdatab_53 datab_53 gnd dc 1.8
Vdata_54 data_54 gnd dc 0 
Vdatab_54 datab_54 gnd dc 1.8
Vdata_55 data_55 gnd dc 0 
Vdatab_55 datab_55 gnd dc 1.8
Vdata_56 data_56 gnd dc 0 
Vdatab_56 datab_56 gnd dc 1.8
Vdata_57 data_57 gnd dc 0 
Vdatab_57 datab_57 gnd dc 1.8
Vdata_58 data_58 gnd dc 0 
Vdatab_58 datab_58 gnd dc 1.8
Vdata_59 data_59 gnd dc 0 
Vdatab_59 datab_59 gnd dc 1.8
Vdata_60 data_60 gnd dc 0 
Vdatab_60 datab_60 gnd dc 1.8
Vdata_61 data_61 gnd dc 0 
Vdatab_61 datab_61 gnd dc 1.8
Vdata_62 data_62 gnd dc 0 
Vdatab_62 datab_62 gnd dc 1.8
Vdata_63 data_63 gnd dc 0 
Vdatab_63 datab_63 gnd dc 1.8
Vdata_64 data_64 gnd dc 0 
Vdatab_64 datab_64 gnd dc 1.8
Vdata_65 data_65 gnd dc 0 
Vdatab_65 datab_65 gnd dc 1.8
Vdata_66 data_66 gnd dc 0 
Vdatab_66 datab_66 gnd dc 1.8
Vdata_67 data_67 gnd dc 0 
Vdatab_67 datab_67 gnd dc 1.8
Vdata_68 data_68 gnd dc 0 
Vdatab_68 datab_68 gnd dc 1.8
Vdata_69 data_69 gnd dc 0 
Vdatab_69 datab_69 gnd dc 1.8
Vdata_70 data_70 gnd dc 0 
Vdatab_70 datab_70 gnd dc 1.8
Vdata_71 data_71 gnd dc 0 
Vdatab_71 datab_71 gnd dc 1.8
Vdata_72 data_72 gnd dc 0 
Vdatab_72 datab_72 gnd dc 1.8
Vdata_73 data_73 gnd dc 0 
Vdatab_73 datab_73 gnd dc 1.8
Vdata_74 data_74 gnd dc 0 
Vdatab_74 datab_74 gnd dc 1.8
Vdata_75 data_75 gnd dc 0 
Vdatab_75 datab_75 gnd dc 1.8
Vdata_76 data_76 gnd dc 0 
Vdatab_76 datab_76 gnd dc 1.8
Vdata_77 data_77 gnd dc 0 
Vdatab_77 datab_77 gnd dc 1.8
Vdata_78 data_78 gnd dc 0 
Vdatab_78 datab_78 gnd dc 1.8
Vdata_79 data_79 gnd dc 0 
Vdatab_79 datab_79 gnd dc 1.8
Vdata_80 data_80 gnd dc 0 
Vdatab_80 datab_80 gnd dc 1.8
Vdata_81 data_81 gnd dc 0 
Vdatab_81 datab_81 gnd dc 1.8
Vdata_82 data_82 gnd dc 0 
Vdatab_82 datab_82 gnd dc 1.8
Vdata_83 data_83 gnd dc 0 
Vdatab_83 datab_83 gnd dc 1.8
Vdata_84 data_84 gnd dc 0 
Vdatab_84 datab_84 gnd dc 1.8
Vdata_85 data_85 gnd dc 0 
Vdatab_85 datab_85 gnd dc 1.8
Vdata_86 data_86 gnd dc 0 
Vdatab_86 datab_86 gnd dc 1.8
Vdata_87 data_87 gnd dc 0 
Vdatab_87 datab_87 gnd dc 1.8
Vdata_88 data_88 gnd dc 0 
Vdatab_88 datab_88 gnd dc 1.8
Vdata_89 data_89 gnd dc 0 
Vdatab_89 datab_89 gnd dc 1.8
Vdata_90 data_90 gnd dc 0 
Vdatab_90 datab_90 gnd dc 1.8
Vdata_91 data_91 gnd dc 0 
Vdatab_91 datab_91 gnd dc 1.8
Vdata_92 data_92 gnd dc 0 
Vdatab_92 datab_92 gnd dc 1.8
Vdata_93 data_93 gnd dc 0 
Vdatab_93 datab_93 gnd dc 1.8
Vdata_94 data_94 gnd dc 0 
Vdatab_94 datab_94 gnd dc 1.8
Vdata_95 data_95 gnd dc 0 
Vdatab_95 datab_95 gnd dc 1.8
Vdata_96 data_96 gnd dc 0 
Vdatab_96 datab_96 gnd dc 1.8
Vdata_97 data_97 gnd dc 0 
Vdatab_97 datab_97 gnd dc 1.8
Vdata_98 data_98 gnd dc 0 
Vdatab_98 datab_98 gnd dc 1.8
Vdata_99 data_99 gnd dc 0 
Vdatab_99 datab_99 gnd dc 1.8
.ic q_0_0=0
.ic qb_0_0=1.8
.ic q_1_0=0
.ic qb_1_0=1.8
.ic q_2_0=0
.ic qb_2_0=1.8
.ic q_3_0=0
.ic qb_3_0=1.8
.ic q_4_0=0
.ic qb_4_0=1.8
.ic q_5_0=0
.ic qb_5_0=1.8
.ic q_6_0=0
.ic qb_6_0=1.8
.ic q_7_0=0
.ic qb_7_0=1.8
.ic q_8_0=0
.ic qb_8_0=1.8
.ic q_9_0=0
.ic qb_9_0=1.8
.ic q_10_0=0
.ic qb_10_0=1.8
.ic q_11_0=0
.ic qb_11_0=1.8
.ic q_12_0=0
.ic qb_12_0=1.8
.ic q_13_0=0
.ic qb_13_0=1.8
.ic q_14_0=0
.ic qb_14_0=1.8
.ic q_15_0=0
.ic qb_15_0=1.8
.ic q_16_0=0
.ic qb_16_0=1.8
.ic q_17_0=0
.ic qb_17_0=1.8
.ic q_18_0=0
.ic qb_18_0=1.8
.ic q_19_0=0
.ic qb_19_0=1.8
.ic q_20_0=0
.ic qb_20_0=1.8
.ic q_21_0=0
.ic qb_21_0=1.8
.ic q_22_0=0
.ic qb_22_0=1.8
.ic q_23_0=0
.ic qb_23_0=1.8
.ic q_24_0=0
.ic qb_24_0=1.8
.ic q_25_0=0
.ic qb_25_0=1.8
.ic q_26_0=0
.ic qb_26_0=1.8
.ic q_27_0=0
.ic qb_27_0=1.8
.ic q_28_0=0
.ic qb_28_0=1.8
.ic q_29_0=0
.ic qb_29_0=1.8
.ic q_30_0=0
.ic qb_30_0=1.8
.ic q_31_0=0
.ic qb_31_0=1.8
.ic q_32_0=0
.ic qb_32_0=1.8
.ic q_33_0=0
.ic qb_33_0=1.8
.ic q_34_0=0
.ic qb_34_0=1.8
.ic q_35_0=0
.ic qb_35_0=1.8
.ic q_36_0=0
.ic qb_36_0=1.8
.ic q_37_0=0
.ic qb_37_0=1.8
.ic q_38_0=0
.ic qb_38_0=1.8
.ic q_39_0=0
.ic qb_39_0=1.8
.ic q_40_0=0
.ic qb_40_0=1.8
.ic q_41_0=0
.ic qb_41_0=1.8
.ic q_42_0=0
.ic qb_42_0=1.8
.ic q_43_0=0
.ic qb_43_0=1.8
.ic q_44_0=0
.ic qb_44_0=1.8
.ic q_45_0=0
.ic qb_45_0=1.8
.ic q_46_0=0
.ic qb_46_0=1.8
.ic q_47_0=0
.ic qb_47_0=1.8
.ic q_48_0=0
.ic qb_48_0=1.8
.ic q_49_0=0
.ic qb_49_0=1.8
.ic q_50_0=0
.ic qb_50_0=1.8
.ic q_51_0=0
.ic qb_51_0=1.8
.ic q_52_0=0
.ic qb_52_0=1.8
.ic q_53_0=0
.ic qb_53_0=1.8
.ic q_54_0=0
.ic qb_54_0=1.8
.ic q_55_0=0
.ic qb_55_0=1.8
.ic q_56_0=0
.ic qb_56_0=1.8
.ic q_57_0=0
.ic qb_57_0=1.8
.ic q_58_0=0
.ic qb_58_0=1.8
.ic q_59_0=0
.ic qb_59_0=1.8
.ic q_60_0=0
.ic qb_60_0=1.8
.ic q_61_0=0
.ic qb_61_0=1.8
.ic q_62_0=0
.ic qb_62_0=1.8
.ic q_63_0=0
.ic qb_63_0=1.8
.ic q_64_0=0
.ic qb_64_0=1.8
.ic q_65_0=0
.ic qb_65_0=1.8
.ic q_66_0=0
.ic qb_66_0=1.8
.ic q_67_0=0
.ic qb_67_0=1.8
.ic q_68_0=0
.ic qb_68_0=1.8
.ic q_69_0=0
.ic qb_69_0=1.8
.ic q_70_0=0
.ic qb_70_0=1.8
.ic q_71_0=0
.ic qb_71_0=1.8
.ic q_72_0=0
.ic qb_72_0=1.8
.ic q_73_0=0
.ic qb_73_0=1.8
.ic q_74_0=0
.ic qb_74_0=1.8
.ic q_75_0=0
.ic qb_75_0=1.8
.ic q_76_0=0
.ic qb_76_0=1.8
.ic q_77_0=0
.ic qb_77_0=1.8
.ic q_78_0=0
.ic qb_78_0=1.8
.ic q_79_0=0
.ic qb_79_0=1.8
.ic q_80_0=0
.ic qb_80_0=1.8
.ic q_81_0=0
.ic qb_81_0=1.8
.ic q_82_0=0
.ic qb_82_0=1.8
.ic q_83_0=0
.ic qb_83_0=1.8
.ic q_84_0=0
.ic qb_84_0=1.8
.ic q_85_0=0
.ic qb_85_0=1.8
.ic q_86_0=0
.ic qb_86_0=1.8
.ic q_87_0=0
.ic qb_87_0=1.8
.ic q_88_0=0
.ic qb_88_0=1.8
.ic q_89_0=0
.ic qb_89_0=1.8
.ic q_90_0=0
.ic qb_90_0=1.8
.ic q_91_0=0
.ic qb_91_0=1.8
.ic q_92_0=0
.ic qb_92_0=1.8
.ic q_93_0=0
.ic qb_93_0=1.8
.ic q_94_0=0
.ic qb_94_0=1.8
.ic q_95_0=0
.ic qb_95_0=1.8
.ic q_96_0=0
.ic qb_96_0=1.8
.ic q_97_0=0
.ic qb_97_0=1.8
.ic q_98_0=0
.ic qb_98_0=1.8
.ic q_99_0=0
.ic qb_99_0=1.8
.ic q_0_1=0
.ic qb_0_1=1.8
.ic q_1_1=0
.ic qb_1_1=1.8
.ic q_2_1=0
.ic qb_2_1=1.8
.ic q_3_1=0
.ic qb_3_1=1.8
.ic q_4_1=0
.ic qb_4_1=1.8
.ic q_5_1=0
.ic qb_5_1=1.8
.ic q_6_1=0
.ic qb_6_1=1.8
.ic q_7_1=0
.ic qb_7_1=1.8
.ic q_8_1=0
.ic qb_8_1=1.8
.ic q_9_1=0
.ic qb_9_1=1.8
.ic q_10_1=0
.ic qb_10_1=1.8
.ic q_11_1=0
.ic qb_11_1=1.8
.ic q_12_1=0
.ic qb_12_1=1.8
.ic q_13_1=0
.ic qb_13_1=1.8
.ic q_14_1=0
.ic qb_14_1=1.8
.ic q_15_1=0
.ic qb_15_1=1.8
.ic q_16_1=0
.ic qb_16_1=1.8
.ic q_17_1=0
.ic qb_17_1=1.8
.ic q_18_1=0
.ic qb_18_1=1.8
.ic q_19_1=0
.ic qb_19_1=1.8
.ic q_20_1=0
.ic qb_20_1=1.8
.ic q_21_1=0
.ic qb_21_1=1.8
.ic q_22_1=0
.ic qb_22_1=1.8
.ic q_23_1=0
.ic qb_23_1=1.8
.ic q_24_1=0
.ic qb_24_1=1.8
.ic q_25_1=0
.ic qb_25_1=1.8
.ic q_26_1=0
.ic qb_26_1=1.8
.ic q_27_1=0
.ic qb_27_1=1.8
.ic q_28_1=0
.ic qb_28_1=1.8
.ic q_29_1=0
.ic qb_29_1=1.8
.ic q_30_1=0
.ic qb_30_1=1.8
.ic q_31_1=0
.ic qb_31_1=1.8
.ic q_32_1=0
.ic qb_32_1=1.8
.ic q_33_1=0
.ic qb_33_1=1.8
.ic q_34_1=0
.ic qb_34_1=1.8
.ic q_35_1=0
.ic qb_35_1=1.8
.ic q_36_1=0
.ic qb_36_1=1.8
.ic q_37_1=0
.ic qb_37_1=1.8
.ic q_38_1=0
.ic qb_38_1=1.8
.ic q_39_1=0
.ic qb_39_1=1.8
.ic q_40_1=0
.ic qb_40_1=1.8
.ic q_41_1=0
.ic qb_41_1=1.8
.ic q_42_1=0
.ic qb_42_1=1.8
.ic q_43_1=0
.ic qb_43_1=1.8
.ic q_44_1=0
.ic qb_44_1=1.8
.ic q_45_1=0
.ic qb_45_1=1.8
.ic q_46_1=0
.ic qb_46_1=1.8
.ic q_47_1=0
.ic qb_47_1=1.8
.ic q_48_1=0
.ic qb_48_1=1.8
.ic q_49_1=0
.ic qb_49_1=1.8
.ic q_50_1=0
.ic qb_50_1=1.8
.ic q_51_1=0
.ic qb_51_1=1.8
.ic q_52_1=0
.ic qb_52_1=1.8
.ic q_53_1=0
.ic qb_53_1=1.8
.ic q_54_1=0
.ic qb_54_1=1.8
.ic q_55_1=0
.ic qb_55_1=1.8
.ic q_56_1=0
.ic qb_56_1=1.8
.ic q_57_1=0
.ic qb_57_1=1.8
.ic q_58_1=0
.ic qb_58_1=1.8
.ic q_59_1=0
.ic qb_59_1=1.8
.ic q_60_1=0
.ic qb_60_1=1.8
.ic q_61_1=0
.ic qb_61_1=1.8
.ic q_62_1=0
.ic qb_62_1=1.8
.ic q_63_1=0
.ic qb_63_1=1.8
.ic q_64_1=0
.ic qb_64_1=1.8
.ic q_65_1=0
.ic qb_65_1=1.8
.ic q_66_1=0
.ic qb_66_1=1.8
.ic q_67_1=0
.ic qb_67_1=1.8
.ic q_68_1=0
.ic qb_68_1=1.8
.ic q_69_1=0
.ic qb_69_1=1.8
.ic q_70_1=0
.ic qb_70_1=1.8
.ic q_71_1=0
.ic qb_71_1=1.8
.ic q_72_1=0
.ic qb_72_1=1.8
.ic q_73_1=0
.ic qb_73_1=1.8
.ic q_74_1=0
.ic qb_74_1=1.8
.ic q_75_1=0
.ic qb_75_1=1.8
.ic q_76_1=0
.ic qb_76_1=1.8
.ic q_77_1=0
.ic qb_77_1=1.8
.ic q_78_1=0
.ic qb_78_1=1.8
.ic q_79_1=0
.ic qb_79_1=1.8
.ic q_80_1=0
.ic qb_80_1=1.8
.ic q_81_1=0
.ic qb_81_1=1.8
.ic q_82_1=0
.ic qb_82_1=1.8
.ic q_83_1=0
.ic qb_83_1=1.8
.ic q_84_1=0
.ic qb_84_1=1.8
.ic q_85_1=0
.ic qb_85_1=1.8
.ic q_86_1=0
.ic qb_86_1=1.8
.ic q_87_1=0
.ic qb_87_1=1.8
.ic q_88_1=0
.ic qb_88_1=1.8
.ic q_89_1=0
.ic qb_89_1=1.8
.ic q_90_1=0
.ic qb_90_1=1.8
.ic q_91_1=0
.ic qb_91_1=1.8
.ic q_92_1=0
.ic qb_92_1=1.8
.ic q_93_1=0
.ic qb_93_1=1.8
.ic q_94_1=0
.ic qb_94_1=1.8
.ic q_95_1=0
.ic qb_95_1=1.8
.ic q_96_1=0
.ic qb_96_1=1.8
.ic q_97_1=0
.ic qb_97_1=1.8
.ic q_98_1=0
.ic qb_98_1=1.8
.ic q_99_1=0
.ic qb_99_1=1.8
.ic q_0_2=0
.ic qb_0_2=1.8
.ic q_1_2=0
.ic qb_1_2=1.8
.ic q_2_2=0
.ic qb_2_2=1.8
.ic q_3_2=0
.ic qb_3_2=1.8
.ic q_4_2=0
.ic qb_4_2=1.8
.ic q_5_2=0
.ic qb_5_2=1.8
.ic q_6_2=0
.ic qb_6_2=1.8
.ic q_7_2=0
.ic qb_7_2=1.8
.ic q_8_2=0
.ic qb_8_2=1.8
.ic q_9_2=0
.ic qb_9_2=1.8
.ic q_10_2=0
.ic qb_10_2=1.8
.ic q_11_2=0
.ic qb_11_2=1.8
.ic q_12_2=0
.ic qb_12_2=1.8
.ic q_13_2=0
.ic qb_13_2=1.8
.ic q_14_2=0
.ic qb_14_2=1.8
.ic q_15_2=0
.ic qb_15_2=1.8
.ic q_16_2=0
.ic qb_16_2=1.8
.ic q_17_2=0
.ic qb_17_2=1.8
.ic q_18_2=0
.ic qb_18_2=1.8
.ic q_19_2=0
.ic qb_19_2=1.8
.ic q_20_2=0
.ic qb_20_2=1.8
.ic q_21_2=0
.ic qb_21_2=1.8
.ic q_22_2=0
.ic qb_22_2=1.8
.ic q_23_2=0
.ic qb_23_2=1.8
.ic q_24_2=0
.ic qb_24_2=1.8
.ic q_25_2=0
.ic qb_25_2=1.8
.ic q_26_2=0
.ic qb_26_2=1.8
.ic q_27_2=0
.ic qb_27_2=1.8
.ic q_28_2=0
.ic qb_28_2=1.8
.ic q_29_2=0
.ic qb_29_2=1.8
.ic q_30_2=0
.ic qb_30_2=1.8
.ic q_31_2=0
.ic qb_31_2=1.8
.ic q_32_2=0
.ic qb_32_2=1.8
.ic q_33_2=0
.ic qb_33_2=1.8
.ic q_34_2=0
.ic qb_34_2=1.8
.ic q_35_2=0
.ic qb_35_2=1.8
.ic q_36_2=0
.ic qb_36_2=1.8
.ic q_37_2=0
.ic qb_37_2=1.8
.ic q_38_2=0
.ic qb_38_2=1.8
.ic q_39_2=0
.ic qb_39_2=1.8
.ic q_40_2=0
.ic qb_40_2=1.8
.ic q_41_2=0
.ic qb_41_2=1.8
.ic q_42_2=0
.ic qb_42_2=1.8
.ic q_43_2=0
.ic qb_43_2=1.8
.ic q_44_2=0
.ic qb_44_2=1.8
.ic q_45_2=0
.ic qb_45_2=1.8
.ic q_46_2=0
.ic qb_46_2=1.8
.ic q_47_2=0
.ic qb_47_2=1.8
.ic q_48_2=0
.ic qb_48_2=1.8
.ic q_49_2=0
.ic qb_49_2=1.8
.ic q_50_2=0
.ic qb_50_2=1.8
.ic q_51_2=0
.ic qb_51_2=1.8
.ic q_52_2=0
.ic qb_52_2=1.8
.ic q_53_2=0
.ic qb_53_2=1.8
.ic q_54_2=0
.ic qb_54_2=1.8
.ic q_55_2=0
.ic qb_55_2=1.8
.ic q_56_2=0
.ic qb_56_2=1.8
.ic q_57_2=0
.ic qb_57_2=1.8
.ic q_58_2=0
.ic qb_58_2=1.8
.ic q_59_2=0
.ic qb_59_2=1.8
.ic q_60_2=0
.ic qb_60_2=1.8
.ic q_61_2=0
.ic qb_61_2=1.8
.ic q_62_2=0
.ic qb_62_2=1.8
.ic q_63_2=0
.ic qb_63_2=1.8
.ic q_64_2=0
.ic qb_64_2=1.8
.ic q_65_2=0
.ic qb_65_2=1.8
.ic q_66_2=0
.ic qb_66_2=1.8
.ic q_67_2=0
.ic qb_67_2=1.8
.ic q_68_2=0
.ic qb_68_2=1.8
.ic q_69_2=0
.ic qb_69_2=1.8
.ic q_70_2=0
.ic qb_70_2=1.8
.ic q_71_2=0
.ic qb_71_2=1.8
.ic q_72_2=0
.ic qb_72_2=1.8
.ic q_73_2=0
.ic qb_73_2=1.8
.ic q_74_2=0
.ic qb_74_2=1.8
.ic q_75_2=0
.ic qb_75_2=1.8
.ic q_76_2=0
.ic qb_76_2=1.8
.ic q_77_2=0
.ic qb_77_2=1.8
.ic q_78_2=0
.ic qb_78_2=1.8
.ic q_79_2=0
.ic qb_79_2=1.8
.ic q_80_2=0
.ic qb_80_2=1.8
.ic q_81_2=0
.ic qb_81_2=1.8
.ic q_82_2=0
.ic qb_82_2=1.8
.ic q_83_2=0
.ic qb_83_2=1.8
.ic q_84_2=0
.ic qb_84_2=1.8
.ic q_85_2=0
.ic qb_85_2=1.8
.ic q_86_2=0
.ic qb_86_2=1.8
.ic q_87_2=0
.ic qb_87_2=1.8
.ic q_88_2=0
.ic qb_88_2=1.8
.ic q_89_2=0
.ic qb_89_2=1.8
.ic q_90_2=0
.ic qb_90_2=1.8
.ic q_91_2=0
.ic qb_91_2=1.8
.ic q_92_2=0
.ic qb_92_2=1.8
.ic q_93_2=0
.ic qb_93_2=1.8
.ic q_94_2=0
.ic qb_94_2=1.8
.ic q_95_2=0
.ic qb_95_2=1.8
.ic q_96_2=0
.ic qb_96_2=1.8
.ic q_97_2=0
.ic qb_97_2=1.8
.ic q_98_2=0
.ic qb_98_2=1.8
.ic q_99_2=0
.ic qb_99_2=1.8
.ic q_0_3=0
.ic qb_0_3=1.8
.ic q_1_3=0
.ic qb_1_3=1.8
.ic q_2_3=0
.ic qb_2_3=1.8
.ic q_3_3=0
.ic qb_3_3=1.8
.ic q_4_3=0
.ic qb_4_3=1.8
.ic q_5_3=0
.ic qb_5_3=1.8
.ic q_6_3=0
.ic qb_6_3=1.8
.ic q_7_3=0
.ic qb_7_3=1.8
.ic q_8_3=0
.ic qb_8_3=1.8
.ic q_9_3=0
.ic qb_9_3=1.8
.ic q_10_3=0
.ic qb_10_3=1.8
.ic q_11_3=0
.ic qb_11_3=1.8
.ic q_12_3=0
.ic qb_12_3=1.8
.ic q_13_3=0
.ic qb_13_3=1.8
.ic q_14_3=0
.ic qb_14_3=1.8
.ic q_15_3=0
.ic qb_15_3=1.8
.ic q_16_3=0
.ic qb_16_3=1.8
.ic q_17_3=0
.ic qb_17_3=1.8
.ic q_18_3=0
.ic qb_18_3=1.8
.ic q_19_3=0
.ic qb_19_3=1.8
.ic q_20_3=0
.ic qb_20_3=1.8
.ic q_21_3=0
.ic qb_21_3=1.8
.ic q_22_3=0
.ic qb_22_3=1.8
.ic q_23_3=0
.ic qb_23_3=1.8
.ic q_24_3=0
.ic qb_24_3=1.8
.ic q_25_3=0
.ic qb_25_3=1.8
.ic q_26_3=0
.ic qb_26_3=1.8
.ic q_27_3=0
.ic qb_27_3=1.8
.ic q_28_3=0
.ic qb_28_3=1.8
.ic q_29_3=0
.ic qb_29_3=1.8
.ic q_30_3=0
.ic qb_30_3=1.8
.ic q_31_3=0
.ic qb_31_3=1.8
.ic q_32_3=0
.ic qb_32_3=1.8
.ic q_33_3=0
.ic qb_33_3=1.8
.ic q_34_3=0
.ic qb_34_3=1.8
.ic q_35_3=0
.ic qb_35_3=1.8
.ic q_36_3=0
.ic qb_36_3=1.8
.ic q_37_3=0
.ic qb_37_3=1.8
.ic q_38_3=0
.ic qb_38_3=1.8
.ic q_39_3=0
.ic qb_39_3=1.8
.ic q_40_3=0
.ic qb_40_3=1.8
.ic q_41_3=0
.ic qb_41_3=1.8
.ic q_42_3=0
.ic qb_42_3=1.8
.ic q_43_3=0
.ic qb_43_3=1.8
.ic q_44_3=0
.ic qb_44_3=1.8
.ic q_45_3=0
.ic qb_45_3=1.8
.ic q_46_3=0
.ic qb_46_3=1.8
.ic q_47_3=0
.ic qb_47_3=1.8
.ic q_48_3=0
.ic qb_48_3=1.8
.ic q_49_3=0
.ic qb_49_3=1.8
.ic q_50_3=0
.ic qb_50_3=1.8
.ic q_51_3=0
.ic qb_51_3=1.8
.ic q_52_3=0
.ic qb_52_3=1.8
.ic q_53_3=0
.ic qb_53_3=1.8
.ic q_54_3=0
.ic qb_54_3=1.8
.ic q_55_3=0
.ic qb_55_3=1.8
.ic q_56_3=0
.ic qb_56_3=1.8
.ic q_57_3=0
.ic qb_57_3=1.8
.ic q_58_3=0
.ic qb_58_3=1.8
.ic q_59_3=0
.ic qb_59_3=1.8
.ic q_60_3=0
.ic qb_60_3=1.8
.ic q_61_3=0
.ic qb_61_3=1.8
.ic q_62_3=0
.ic qb_62_3=1.8
.ic q_63_3=0
.ic qb_63_3=1.8
.ic q_64_3=0
.ic qb_64_3=1.8
.ic q_65_3=0
.ic qb_65_3=1.8
.ic q_66_3=0
.ic qb_66_3=1.8
.ic q_67_3=0
.ic qb_67_3=1.8
.ic q_68_3=0
.ic qb_68_3=1.8
.ic q_69_3=0
.ic qb_69_3=1.8
.ic q_70_3=0
.ic qb_70_3=1.8
.ic q_71_3=0
.ic qb_71_3=1.8
.ic q_72_3=0
.ic qb_72_3=1.8
.ic q_73_3=0
.ic qb_73_3=1.8
.ic q_74_3=0
.ic qb_74_3=1.8
.ic q_75_3=0
.ic qb_75_3=1.8
.ic q_76_3=0
.ic qb_76_3=1.8
.ic q_77_3=0
.ic qb_77_3=1.8
.ic q_78_3=0
.ic qb_78_3=1.8
.ic q_79_3=0
.ic qb_79_3=1.8
.ic q_80_3=0
.ic qb_80_3=1.8
.ic q_81_3=0
.ic qb_81_3=1.8
.ic q_82_3=0
.ic qb_82_3=1.8
.ic q_83_3=0
.ic qb_83_3=1.8
.ic q_84_3=0
.ic qb_84_3=1.8
.ic q_85_3=0
.ic qb_85_3=1.8
.ic q_86_3=0
.ic qb_86_3=1.8
.ic q_87_3=0
.ic qb_87_3=1.8
.ic q_88_3=0
.ic qb_88_3=1.8
.ic q_89_3=0
.ic qb_89_3=1.8
.ic q_90_3=0
.ic qb_90_3=1.8
.ic q_91_3=0
.ic qb_91_3=1.8
.ic q_92_3=0
.ic qb_92_3=1.8
.ic q_93_3=0
.ic qb_93_3=1.8
.ic q_94_3=0
.ic qb_94_3=1.8
.ic q_95_3=0
.ic qb_95_3=1.8
.ic q_96_3=0
.ic qb_96_3=1.8
.ic q_97_3=0
.ic qb_97_3=1.8
.ic q_98_3=0
.ic qb_98_3=1.8
.ic q_99_3=0
.ic qb_99_3=1.8
.ic q_0_4=0
.ic qb_0_4=1.8
.ic q_1_4=0
.ic qb_1_4=1.8
.ic q_2_4=0
.ic qb_2_4=1.8
.ic q_3_4=0
.ic qb_3_4=1.8
.ic q_4_4=0
.ic qb_4_4=1.8
.ic q_5_4=0
.ic qb_5_4=1.8
.ic q_6_4=0
.ic qb_6_4=1.8
.ic q_7_4=0
.ic qb_7_4=1.8
.ic q_8_4=0
.ic qb_8_4=1.8
.ic q_9_4=0
.ic qb_9_4=1.8
.ic q_10_4=0
.ic qb_10_4=1.8
.ic q_11_4=0
.ic qb_11_4=1.8
.ic q_12_4=0
.ic qb_12_4=1.8
.ic q_13_4=0
.ic qb_13_4=1.8
.ic q_14_4=0
.ic qb_14_4=1.8
.ic q_15_4=0
.ic qb_15_4=1.8
.ic q_16_4=0
.ic qb_16_4=1.8
.ic q_17_4=0
.ic qb_17_4=1.8
.ic q_18_4=0
.ic qb_18_4=1.8
.ic q_19_4=0
.ic qb_19_4=1.8
.ic q_20_4=0
.ic qb_20_4=1.8
.ic q_21_4=0
.ic qb_21_4=1.8
.ic q_22_4=0
.ic qb_22_4=1.8
.ic q_23_4=0
.ic qb_23_4=1.8
.ic q_24_4=0
.ic qb_24_4=1.8
.ic q_25_4=0
.ic qb_25_4=1.8
.ic q_26_4=0
.ic qb_26_4=1.8
.ic q_27_4=0
.ic qb_27_4=1.8
.ic q_28_4=0
.ic qb_28_4=1.8
.ic q_29_4=0
.ic qb_29_4=1.8
.ic q_30_4=0
.ic qb_30_4=1.8
.ic q_31_4=0
.ic qb_31_4=1.8
.ic q_32_4=0
.ic qb_32_4=1.8
.ic q_33_4=0
.ic qb_33_4=1.8
.ic q_34_4=0
.ic qb_34_4=1.8
.ic q_35_4=0
.ic qb_35_4=1.8
.ic q_36_4=0
.ic qb_36_4=1.8
.ic q_37_4=0
.ic qb_37_4=1.8
.ic q_38_4=0
.ic qb_38_4=1.8
.ic q_39_4=0
.ic qb_39_4=1.8
.ic q_40_4=0
.ic qb_40_4=1.8
.ic q_41_4=0
.ic qb_41_4=1.8
.ic q_42_4=0
.ic qb_42_4=1.8
.ic q_43_4=0
.ic qb_43_4=1.8
.ic q_44_4=0
.ic qb_44_4=1.8
.ic q_45_4=0
.ic qb_45_4=1.8
.ic q_46_4=0
.ic qb_46_4=1.8
.ic q_47_4=0
.ic qb_47_4=1.8
.ic q_48_4=0
.ic qb_48_4=1.8
.ic q_49_4=0
.ic qb_49_4=1.8
.ic q_50_4=0
.ic qb_50_4=1.8
.ic q_51_4=0
.ic qb_51_4=1.8
.ic q_52_4=0
.ic qb_52_4=1.8
.ic q_53_4=0
.ic qb_53_4=1.8
.ic q_54_4=0
.ic qb_54_4=1.8
.ic q_55_4=0
.ic qb_55_4=1.8
.ic q_56_4=0
.ic qb_56_4=1.8
.ic q_57_4=0
.ic qb_57_4=1.8
.ic q_58_4=0
.ic qb_58_4=1.8
.ic q_59_4=0
.ic qb_59_4=1.8
.ic q_60_4=0
.ic qb_60_4=1.8
.ic q_61_4=0
.ic qb_61_4=1.8
.ic q_62_4=0
.ic qb_62_4=1.8
.ic q_63_4=0
.ic qb_63_4=1.8
.ic q_64_4=0
.ic qb_64_4=1.8
.ic q_65_4=0
.ic qb_65_4=1.8
.ic q_66_4=0
.ic qb_66_4=1.8
.ic q_67_4=0
.ic qb_67_4=1.8
.ic q_68_4=0
.ic qb_68_4=1.8
.ic q_69_4=0
.ic qb_69_4=1.8
.ic q_70_4=0
.ic qb_70_4=1.8
.ic q_71_4=0
.ic qb_71_4=1.8
.ic q_72_4=0
.ic qb_72_4=1.8
.ic q_73_4=0
.ic qb_73_4=1.8
.ic q_74_4=0
.ic qb_74_4=1.8
.ic q_75_4=0
.ic qb_75_4=1.8
.ic q_76_4=0
.ic qb_76_4=1.8
.ic q_77_4=0
.ic qb_77_4=1.8
.ic q_78_4=0
.ic qb_78_4=1.8
.ic q_79_4=0
.ic qb_79_4=1.8
.ic q_80_4=0
.ic qb_80_4=1.8
.ic q_81_4=0
.ic qb_81_4=1.8
.ic q_82_4=0
.ic qb_82_4=1.8
.ic q_83_4=0
.ic qb_83_4=1.8
.ic q_84_4=0
.ic qb_84_4=1.8
.ic q_85_4=0
.ic qb_85_4=1.8
.ic q_86_4=0
.ic qb_86_4=1.8
.ic q_87_4=0
.ic qb_87_4=1.8
.ic q_88_4=0
.ic qb_88_4=1.8
.ic q_89_4=0
.ic qb_89_4=1.8
.ic q_90_4=0
.ic qb_90_4=1.8
.ic q_91_4=0
.ic qb_91_4=1.8
.ic q_92_4=0
.ic qb_92_4=1.8
.ic q_93_4=0
.ic qb_93_4=1.8
.ic q_94_4=0
.ic qb_94_4=1.8
.ic q_95_4=0
.ic qb_95_4=1.8
.ic q_96_4=0
.ic qb_96_4=1.8
.ic q_97_4=0
.ic qb_97_4=1.8
.ic q_98_4=0
.ic qb_98_4=1.8
.ic q_99_4=0
.ic qb_99_4=1.8
.ic q_0_5=0
.ic qb_0_5=1.8
.ic q_1_5=0
.ic qb_1_5=1.8
.ic q_2_5=0
.ic qb_2_5=1.8
.ic q_3_5=0
.ic qb_3_5=1.8
.ic q_4_5=0
.ic qb_4_5=1.8
.ic q_5_5=0
.ic qb_5_5=1.8
.ic q_6_5=0
.ic qb_6_5=1.8
.ic q_7_5=0
.ic qb_7_5=1.8
.ic q_8_5=0
.ic qb_8_5=1.8
.ic q_9_5=0
.ic qb_9_5=1.8
.ic q_10_5=0
.ic qb_10_5=1.8
.ic q_11_5=0
.ic qb_11_5=1.8
.ic q_12_5=0
.ic qb_12_5=1.8
.ic q_13_5=0
.ic qb_13_5=1.8
.ic q_14_5=0
.ic qb_14_5=1.8
.ic q_15_5=0
.ic qb_15_5=1.8
.ic q_16_5=0
.ic qb_16_5=1.8
.ic q_17_5=0
.ic qb_17_5=1.8
.ic q_18_5=0
.ic qb_18_5=1.8
.ic q_19_5=0
.ic qb_19_5=1.8
.ic q_20_5=0
.ic qb_20_5=1.8
.ic q_21_5=0
.ic qb_21_5=1.8
.ic q_22_5=0
.ic qb_22_5=1.8
.ic q_23_5=0
.ic qb_23_5=1.8
.ic q_24_5=0
.ic qb_24_5=1.8
.ic q_25_5=0
.ic qb_25_5=1.8
.ic q_26_5=0
.ic qb_26_5=1.8
.ic q_27_5=0
.ic qb_27_5=1.8
.ic q_28_5=0
.ic qb_28_5=1.8
.ic q_29_5=0
.ic qb_29_5=1.8
.ic q_30_5=0
.ic qb_30_5=1.8
.ic q_31_5=0
.ic qb_31_5=1.8
.ic q_32_5=0
.ic qb_32_5=1.8
.ic q_33_5=0
.ic qb_33_5=1.8
.ic q_34_5=0
.ic qb_34_5=1.8
.ic q_35_5=0
.ic qb_35_5=1.8
.ic q_36_5=0
.ic qb_36_5=1.8
.ic q_37_5=0
.ic qb_37_5=1.8
.ic q_38_5=0
.ic qb_38_5=1.8
.ic q_39_5=0
.ic qb_39_5=1.8
.ic q_40_5=0
.ic qb_40_5=1.8
.ic q_41_5=0
.ic qb_41_5=1.8
.ic q_42_5=0
.ic qb_42_5=1.8
.ic q_43_5=0
.ic qb_43_5=1.8
.ic q_44_5=0
.ic qb_44_5=1.8
.ic q_45_5=0
.ic qb_45_5=1.8
.ic q_46_5=0
.ic qb_46_5=1.8
.ic q_47_5=0
.ic qb_47_5=1.8
.ic q_48_5=0
.ic qb_48_5=1.8
.ic q_49_5=0
.ic qb_49_5=1.8
.ic q_50_5=0
.ic qb_50_5=1.8
.ic q_51_5=0
.ic qb_51_5=1.8
.ic q_52_5=0
.ic qb_52_5=1.8
.ic q_53_5=0
.ic qb_53_5=1.8
.ic q_54_5=0
.ic qb_54_5=1.8
.ic q_55_5=0
.ic qb_55_5=1.8
.ic q_56_5=0
.ic qb_56_5=1.8
.ic q_57_5=0
.ic qb_57_5=1.8
.ic q_58_5=0
.ic qb_58_5=1.8
.ic q_59_5=0
.ic qb_59_5=1.8
.ic q_60_5=0
.ic qb_60_5=1.8
.ic q_61_5=0
.ic qb_61_5=1.8
.ic q_62_5=0
.ic qb_62_5=1.8
.ic q_63_5=0
.ic qb_63_5=1.8
.ic q_64_5=0
.ic qb_64_5=1.8
.ic q_65_5=0
.ic qb_65_5=1.8
.ic q_66_5=0
.ic qb_66_5=1.8
.ic q_67_5=0
.ic qb_67_5=1.8
.ic q_68_5=0
.ic qb_68_5=1.8
.ic q_69_5=0
.ic qb_69_5=1.8
.ic q_70_5=0
.ic qb_70_5=1.8
.ic q_71_5=0
.ic qb_71_5=1.8
.ic q_72_5=0
.ic qb_72_5=1.8
.ic q_73_5=0
.ic qb_73_5=1.8
.ic q_74_5=0
.ic qb_74_5=1.8
.ic q_75_5=0
.ic qb_75_5=1.8
.ic q_76_5=0
.ic qb_76_5=1.8
.ic q_77_5=0
.ic qb_77_5=1.8
.ic q_78_5=0
.ic qb_78_5=1.8
.ic q_79_5=0
.ic qb_79_5=1.8
.ic q_80_5=0
.ic qb_80_5=1.8
.ic q_81_5=0
.ic qb_81_5=1.8
.ic q_82_5=0
.ic qb_82_5=1.8
.ic q_83_5=0
.ic qb_83_5=1.8
.ic q_84_5=0
.ic qb_84_5=1.8
.ic q_85_5=0
.ic qb_85_5=1.8
.ic q_86_5=0
.ic qb_86_5=1.8
.ic q_87_5=0
.ic qb_87_5=1.8
.ic q_88_5=0
.ic qb_88_5=1.8
.ic q_89_5=0
.ic qb_89_5=1.8
.ic q_90_5=0
.ic qb_90_5=1.8
.ic q_91_5=0
.ic qb_91_5=1.8
.ic q_92_5=0
.ic qb_92_5=1.8
.ic q_93_5=0
.ic qb_93_5=1.8
.ic q_94_5=0
.ic qb_94_5=1.8
.ic q_95_5=0
.ic qb_95_5=1.8
.ic q_96_5=0
.ic qb_96_5=1.8
.ic q_97_5=0
.ic qb_97_5=1.8
.ic q_98_5=0
.ic qb_98_5=1.8
.ic q_99_5=0
.ic qb_99_5=1.8
.ic q_0_6=0
.ic qb_0_6=1.8
.ic q_1_6=0
.ic qb_1_6=1.8
.ic q_2_6=0
.ic qb_2_6=1.8
.ic q_3_6=0
.ic qb_3_6=1.8
.ic q_4_6=0
.ic qb_4_6=1.8
.ic q_5_6=0
.ic qb_5_6=1.8
.ic q_6_6=0
.ic qb_6_6=1.8
.ic q_7_6=0
.ic qb_7_6=1.8
.ic q_8_6=0
.ic qb_8_6=1.8
.ic q_9_6=0
.ic qb_9_6=1.8
.ic q_10_6=0
.ic qb_10_6=1.8
.ic q_11_6=0
.ic qb_11_6=1.8
.ic q_12_6=0
.ic qb_12_6=1.8
.ic q_13_6=0
.ic qb_13_6=1.8
.ic q_14_6=0
.ic qb_14_6=1.8
.ic q_15_6=0
.ic qb_15_6=1.8
.ic q_16_6=0
.ic qb_16_6=1.8
.ic q_17_6=0
.ic qb_17_6=1.8
.ic q_18_6=0
.ic qb_18_6=1.8
.ic q_19_6=0
.ic qb_19_6=1.8
.ic q_20_6=0
.ic qb_20_6=1.8
.ic q_21_6=0
.ic qb_21_6=1.8
.ic q_22_6=0
.ic qb_22_6=1.8
.ic q_23_6=0
.ic qb_23_6=1.8
.ic q_24_6=0
.ic qb_24_6=1.8
.ic q_25_6=0
.ic qb_25_6=1.8
.ic q_26_6=0
.ic qb_26_6=1.8
.ic q_27_6=0
.ic qb_27_6=1.8
.ic q_28_6=0
.ic qb_28_6=1.8
.ic q_29_6=0
.ic qb_29_6=1.8
.ic q_30_6=0
.ic qb_30_6=1.8
.ic q_31_6=0
.ic qb_31_6=1.8
.ic q_32_6=0
.ic qb_32_6=1.8
.ic q_33_6=0
.ic qb_33_6=1.8
.ic q_34_6=0
.ic qb_34_6=1.8
.ic q_35_6=0
.ic qb_35_6=1.8
.ic q_36_6=0
.ic qb_36_6=1.8
.ic q_37_6=0
.ic qb_37_6=1.8
.ic q_38_6=0
.ic qb_38_6=1.8
.ic q_39_6=0
.ic qb_39_6=1.8
.ic q_40_6=0
.ic qb_40_6=1.8
.ic q_41_6=0
.ic qb_41_6=1.8
.ic q_42_6=0
.ic qb_42_6=1.8
.ic q_43_6=0
.ic qb_43_6=1.8
.ic q_44_6=0
.ic qb_44_6=1.8
.ic q_45_6=0
.ic qb_45_6=1.8
.ic q_46_6=0
.ic qb_46_6=1.8
.ic q_47_6=0
.ic qb_47_6=1.8
.ic q_48_6=0
.ic qb_48_6=1.8
.ic q_49_6=0
.ic qb_49_6=1.8
.ic q_50_6=0
.ic qb_50_6=1.8
.ic q_51_6=0
.ic qb_51_6=1.8
.ic q_52_6=0
.ic qb_52_6=1.8
.ic q_53_6=0
.ic qb_53_6=1.8
.ic q_54_6=0
.ic qb_54_6=1.8
.ic q_55_6=0
.ic qb_55_6=1.8
.ic q_56_6=0
.ic qb_56_6=1.8
.ic q_57_6=0
.ic qb_57_6=1.8
.ic q_58_6=0
.ic qb_58_6=1.8
.ic q_59_6=0
.ic qb_59_6=1.8
.ic q_60_6=0
.ic qb_60_6=1.8
.ic q_61_6=0
.ic qb_61_6=1.8
.ic q_62_6=0
.ic qb_62_6=1.8
.ic q_63_6=0
.ic qb_63_6=1.8
.ic q_64_6=0
.ic qb_64_6=1.8
.ic q_65_6=0
.ic qb_65_6=1.8
.ic q_66_6=0
.ic qb_66_6=1.8
.ic q_67_6=0
.ic qb_67_6=1.8
.ic q_68_6=0
.ic qb_68_6=1.8
.ic q_69_6=0
.ic qb_69_6=1.8
.ic q_70_6=0
.ic qb_70_6=1.8
.ic q_71_6=0
.ic qb_71_6=1.8
.ic q_72_6=0
.ic qb_72_6=1.8
.ic q_73_6=0
.ic qb_73_6=1.8
.ic q_74_6=0
.ic qb_74_6=1.8
.ic q_75_6=0
.ic qb_75_6=1.8
.ic q_76_6=0
.ic qb_76_6=1.8
.ic q_77_6=0
.ic qb_77_6=1.8
.ic q_78_6=0
.ic qb_78_6=1.8
.ic q_79_6=0
.ic qb_79_6=1.8
.ic q_80_6=0
.ic qb_80_6=1.8
.ic q_81_6=0
.ic qb_81_6=1.8
.ic q_82_6=0
.ic qb_82_6=1.8
.ic q_83_6=0
.ic qb_83_6=1.8
.ic q_84_6=0
.ic qb_84_6=1.8
.ic q_85_6=0
.ic qb_85_6=1.8
.ic q_86_6=0
.ic qb_86_6=1.8
.ic q_87_6=0
.ic qb_87_6=1.8
.ic q_88_6=0
.ic qb_88_6=1.8
.ic q_89_6=0
.ic qb_89_6=1.8
.ic q_90_6=0
.ic qb_90_6=1.8
.ic q_91_6=0
.ic qb_91_6=1.8
.ic q_92_6=0
.ic qb_92_6=1.8
.ic q_93_6=0
.ic qb_93_6=1.8
.ic q_94_6=0
.ic qb_94_6=1.8
.ic q_95_6=0
.ic qb_95_6=1.8
.ic q_96_6=0
.ic qb_96_6=1.8
.ic q_97_6=0
.ic qb_97_6=1.8
.ic q_98_6=0
.ic qb_98_6=1.8
.ic q_99_6=0
.ic qb_99_6=1.8
.ic q_0_7=0
.ic qb_0_7=1.8
.ic q_1_7=0
.ic qb_1_7=1.8
.ic q_2_7=0
.ic qb_2_7=1.8
.ic q_3_7=0
.ic qb_3_7=1.8
.ic q_4_7=0
.ic qb_4_7=1.8
.ic q_5_7=0
.ic qb_5_7=1.8
.ic q_6_7=0
.ic qb_6_7=1.8
.ic q_7_7=0
.ic qb_7_7=1.8
.ic q_8_7=0
.ic qb_8_7=1.8
.ic q_9_7=0
.ic qb_9_7=1.8
.ic q_10_7=0
.ic qb_10_7=1.8
.ic q_11_7=0
.ic qb_11_7=1.8
.ic q_12_7=0
.ic qb_12_7=1.8
.ic q_13_7=0
.ic qb_13_7=1.8
.ic q_14_7=0
.ic qb_14_7=1.8
.ic q_15_7=0
.ic qb_15_7=1.8
.ic q_16_7=0
.ic qb_16_7=1.8
.ic q_17_7=0
.ic qb_17_7=1.8
.ic q_18_7=0
.ic qb_18_7=1.8
.ic q_19_7=0
.ic qb_19_7=1.8
.ic q_20_7=0
.ic qb_20_7=1.8
.ic q_21_7=0
.ic qb_21_7=1.8
.ic q_22_7=0
.ic qb_22_7=1.8
.ic q_23_7=0
.ic qb_23_7=1.8
.ic q_24_7=0
.ic qb_24_7=1.8
.ic q_25_7=0
.ic qb_25_7=1.8
.ic q_26_7=0
.ic qb_26_7=1.8
.ic q_27_7=0
.ic qb_27_7=1.8
.ic q_28_7=0
.ic qb_28_7=1.8
.ic q_29_7=0
.ic qb_29_7=1.8
.ic q_30_7=0
.ic qb_30_7=1.8
.ic q_31_7=0
.ic qb_31_7=1.8
.ic q_32_7=0
.ic qb_32_7=1.8
.ic q_33_7=0
.ic qb_33_7=1.8
.ic q_34_7=0
.ic qb_34_7=1.8
.ic q_35_7=0
.ic qb_35_7=1.8
.ic q_36_7=0
.ic qb_36_7=1.8
.ic q_37_7=0
.ic qb_37_7=1.8
.ic q_38_7=0
.ic qb_38_7=1.8
.ic q_39_7=0
.ic qb_39_7=1.8
.ic q_40_7=0
.ic qb_40_7=1.8
.ic q_41_7=0
.ic qb_41_7=1.8
.ic q_42_7=0
.ic qb_42_7=1.8
.ic q_43_7=0
.ic qb_43_7=1.8
.ic q_44_7=0
.ic qb_44_7=1.8
.ic q_45_7=0
.ic qb_45_7=1.8
.ic q_46_7=0
.ic qb_46_7=1.8
.ic q_47_7=0
.ic qb_47_7=1.8
.ic q_48_7=0
.ic qb_48_7=1.8
.ic q_49_7=0
.ic qb_49_7=1.8
.ic q_50_7=0
.ic qb_50_7=1.8
.ic q_51_7=0
.ic qb_51_7=1.8
.ic q_52_7=0
.ic qb_52_7=1.8
.ic q_53_7=0
.ic qb_53_7=1.8
.ic q_54_7=0
.ic qb_54_7=1.8
.ic q_55_7=0
.ic qb_55_7=1.8
.ic q_56_7=0
.ic qb_56_7=1.8
.ic q_57_7=0
.ic qb_57_7=1.8
.ic q_58_7=0
.ic qb_58_7=1.8
.ic q_59_7=0
.ic qb_59_7=1.8
.ic q_60_7=0
.ic qb_60_7=1.8
.ic q_61_7=0
.ic qb_61_7=1.8
.ic q_62_7=0
.ic qb_62_7=1.8
.ic q_63_7=0
.ic qb_63_7=1.8
.ic q_64_7=0
.ic qb_64_7=1.8
.ic q_65_7=0
.ic qb_65_7=1.8
.ic q_66_7=0
.ic qb_66_7=1.8
.ic q_67_7=0
.ic qb_67_7=1.8
.ic q_68_7=0
.ic qb_68_7=1.8
.ic q_69_7=0
.ic qb_69_7=1.8
.ic q_70_7=0
.ic qb_70_7=1.8
.ic q_71_7=0
.ic qb_71_7=1.8
.ic q_72_7=0
.ic qb_72_7=1.8
.ic q_73_7=0
.ic qb_73_7=1.8
.ic q_74_7=0
.ic qb_74_7=1.8
.ic q_75_7=0
.ic qb_75_7=1.8
.ic q_76_7=0
.ic qb_76_7=1.8
.ic q_77_7=0
.ic qb_77_7=1.8
.ic q_78_7=0
.ic qb_78_7=1.8
.ic q_79_7=0
.ic qb_79_7=1.8
.ic q_80_7=0
.ic qb_80_7=1.8
.ic q_81_7=0
.ic qb_81_7=1.8
.ic q_82_7=0
.ic qb_82_7=1.8
.ic q_83_7=0
.ic qb_83_7=1.8
.ic q_84_7=0
.ic qb_84_7=1.8
.ic q_85_7=0
.ic qb_85_7=1.8
.ic q_86_7=0
.ic qb_86_7=1.8
.ic q_87_7=0
.ic qb_87_7=1.8
.ic q_88_7=0
.ic qb_88_7=1.8
.ic q_89_7=0
.ic qb_89_7=1.8
.ic q_90_7=0
.ic qb_90_7=1.8
.ic q_91_7=0
.ic qb_91_7=1.8
.ic q_92_7=0
.ic qb_92_7=1.8
.ic q_93_7=0
.ic qb_93_7=1.8
.ic q_94_7=0
.ic qb_94_7=1.8
.ic q_95_7=0
.ic qb_95_7=1.8
.ic q_96_7=0
.ic qb_96_7=1.8
.ic q_97_7=0
.ic qb_97_7=1.8
.ic q_98_7=0
.ic qb_98_7=1.8
.ic q_99_7=0
.ic qb_99_7=1.8
.ic q_0_8=0
.ic qb_0_8=1.8
.ic q_1_8=0
.ic qb_1_8=1.8
.ic q_2_8=0
.ic qb_2_8=1.8
.ic q_3_8=0
.ic qb_3_8=1.8
.ic q_4_8=0
.ic qb_4_8=1.8
.ic q_5_8=0
.ic qb_5_8=1.8
.ic q_6_8=0
.ic qb_6_8=1.8
.ic q_7_8=0
.ic qb_7_8=1.8
.ic q_8_8=0
.ic qb_8_8=1.8
.ic q_9_8=0
.ic qb_9_8=1.8
.ic q_10_8=0
.ic qb_10_8=1.8
.ic q_11_8=0
.ic qb_11_8=1.8
.ic q_12_8=0
.ic qb_12_8=1.8
.ic q_13_8=0
.ic qb_13_8=1.8
.ic q_14_8=0
.ic qb_14_8=1.8
.ic q_15_8=0
.ic qb_15_8=1.8
.ic q_16_8=0
.ic qb_16_8=1.8
.ic q_17_8=0
.ic qb_17_8=1.8
.ic q_18_8=0
.ic qb_18_8=1.8
.ic q_19_8=0
.ic qb_19_8=1.8
.ic q_20_8=0
.ic qb_20_8=1.8
.ic q_21_8=0
.ic qb_21_8=1.8
.ic q_22_8=0
.ic qb_22_8=1.8
.ic q_23_8=0
.ic qb_23_8=1.8
.ic q_24_8=0
.ic qb_24_8=1.8
.ic q_25_8=0
.ic qb_25_8=1.8
.ic q_26_8=0
.ic qb_26_8=1.8
.ic q_27_8=0
.ic qb_27_8=1.8
.ic q_28_8=0
.ic qb_28_8=1.8
.ic q_29_8=0
.ic qb_29_8=1.8
.ic q_30_8=0
.ic qb_30_8=1.8
.ic q_31_8=0
.ic qb_31_8=1.8
.ic q_32_8=0
.ic qb_32_8=1.8
.ic q_33_8=0
.ic qb_33_8=1.8
.ic q_34_8=0
.ic qb_34_8=1.8
.ic q_35_8=0
.ic qb_35_8=1.8
.ic q_36_8=0
.ic qb_36_8=1.8
.ic q_37_8=0
.ic qb_37_8=1.8
.ic q_38_8=0
.ic qb_38_8=1.8
.ic q_39_8=0
.ic qb_39_8=1.8
.ic q_40_8=0
.ic qb_40_8=1.8
.ic q_41_8=0
.ic qb_41_8=1.8
.ic q_42_8=0
.ic qb_42_8=1.8
.ic q_43_8=0
.ic qb_43_8=1.8
.ic q_44_8=0
.ic qb_44_8=1.8
.ic q_45_8=0
.ic qb_45_8=1.8
.ic q_46_8=0
.ic qb_46_8=1.8
.ic q_47_8=0
.ic qb_47_8=1.8
.ic q_48_8=0
.ic qb_48_8=1.8
.ic q_49_8=0
.ic qb_49_8=1.8
.ic q_50_8=0
.ic qb_50_8=1.8
.ic q_51_8=0
.ic qb_51_8=1.8
.ic q_52_8=0
.ic qb_52_8=1.8
.ic q_53_8=0
.ic qb_53_8=1.8
.ic q_54_8=0
.ic qb_54_8=1.8
.ic q_55_8=0
.ic qb_55_8=1.8
.ic q_56_8=0
.ic qb_56_8=1.8
.ic q_57_8=0
.ic qb_57_8=1.8
.ic q_58_8=0
.ic qb_58_8=1.8
.ic q_59_8=0
.ic qb_59_8=1.8
.ic q_60_8=0
.ic qb_60_8=1.8
.ic q_61_8=0
.ic qb_61_8=1.8
.ic q_62_8=0
.ic qb_62_8=1.8
.ic q_63_8=0
.ic qb_63_8=1.8
.ic q_64_8=0
.ic qb_64_8=1.8
.ic q_65_8=0
.ic qb_65_8=1.8
.ic q_66_8=0
.ic qb_66_8=1.8
.ic q_67_8=0
.ic qb_67_8=1.8
.ic q_68_8=0
.ic qb_68_8=1.8
.ic q_69_8=0
.ic qb_69_8=1.8
.ic q_70_8=0
.ic qb_70_8=1.8
.ic q_71_8=0
.ic qb_71_8=1.8
.ic q_72_8=0
.ic qb_72_8=1.8
.ic q_73_8=0
.ic qb_73_8=1.8
.ic q_74_8=0
.ic qb_74_8=1.8
.ic q_75_8=0
.ic qb_75_8=1.8
.ic q_76_8=0
.ic qb_76_8=1.8
.ic q_77_8=0
.ic qb_77_8=1.8
.ic q_78_8=0
.ic qb_78_8=1.8
.ic q_79_8=0
.ic qb_79_8=1.8
.ic q_80_8=0
.ic qb_80_8=1.8
.ic q_81_8=0
.ic qb_81_8=1.8
.ic q_82_8=0
.ic qb_82_8=1.8
.ic q_83_8=0
.ic qb_83_8=1.8
.ic q_84_8=0
.ic qb_84_8=1.8
.ic q_85_8=0
.ic qb_85_8=1.8
.ic q_86_8=0
.ic qb_86_8=1.8
.ic q_87_8=0
.ic qb_87_8=1.8
.ic q_88_8=0
.ic qb_88_8=1.8
.ic q_89_8=0
.ic qb_89_8=1.8
.ic q_90_8=0
.ic qb_90_8=1.8
.ic q_91_8=0
.ic qb_91_8=1.8
.ic q_92_8=0
.ic qb_92_8=1.8
.ic q_93_8=0
.ic qb_93_8=1.8
.ic q_94_8=0
.ic qb_94_8=1.8
.ic q_95_8=0
.ic qb_95_8=1.8
.ic q_96_8=0
.ic qb_96_8=1.8
.ic q_97_8=0
.ic qb_97_8=1.8
.ic q_98_8=0
.ic qb_98_8=1.8
.ic q_99_8=0
.ic qb_99_8=1.8
.ic q_0_9=0
.ic qb_0_9=1.8
.ic q_1_9=0
.ic qb_1_9=1.8
.ic q_2_9=0
.ic qb_2_9=1.8
.ic q_3_9=0
.ic qb_3_9=1.8
.ic q_4_9=0
.ic qb_4_9=1.8
.ic q_5_9=0
.ic qb_5_9=1.8
.ic q_6_9=0
.ic qb_6_9=1.8
.ic q_7_9=0
.ic qb_7_9=1.8
.ic q_8_9=0
.ic qb_8_9=1.8
.ic q_9_9=0
.ic qb_9_9=1.8
.ic q_10_9=0
.ic qb_10_9=1.8
.ic q_11_9=0
.ic qb_11_9=1.8
.ic q_12_9=0
.ic qb_12_9=1.8
.ic q_13_9=0
.ic qb_13_9=1.8
.ic q_14_9=0
.ic qb_14_9=1.8
.ic q_15_9=0
.ic qb_15_9=1.8
.ic q_16_9=0
.ic qb_16_9=1.8
.ic q_17_9=0
.ic qb_17_9=1.8
.ic q_18_9=0
.ic qb_18_9=1.8
.ic q_19_9=0
.ic qb_19_9=1.8
.ic q_20_9=0
.ic qb_20_9=1.8
.ic q_21_9=0
.ic qb_21_9=1.8
.ic q_22_9=0
.ic qb_22_9=1.8
.ic q_23_9=0
.ic qb_23_9=1.8
.ic q_24_9=0
.ic qb_24_9=1.8
.ic q_25_9=0
.ic qb_25_9=1.8
.ic q_26_9=0
.ic qb_26_9=1.8
.ic q_27_9=0
.ic qb_27_9=1.8
.ic q_28_9=0
.ic qb_28_9=1.8
.ic q_29_9=0
.ic qb_29_9=1.8
.ic q_30_9=0
.ic qb_30_9=1.8
.ic q_31_9=0
.ic qb_31_9=1.8
.ic q_32_9=0
.ic qb_32_9=1.8
.ic q_33_9=0
.ic qb_33_9=1.8
.ic q_34_9=0
.ic qb_34_9=1.8
.ic q_35_9=0
.ic qb_35_9=1.8
.ic q_36_9=0
.ic qb_36_9=1.8
.ic q_37_9=0
.ic qb_37_9=1.8
.ic q_38_9=0
.ic qb_38_9=1.8
.ic q_39_9=0
.ic qb_39_9=1.8
.ic q_40_9=0
.ic qb_40_9=1.8
.ic q_41_9=0
.ic qb_41_9=1.8
.ic q_42_9=0
.ic qb_42_9=1.8
.ic q_43_9=0
.ic qb_43_9=1.8
.ic q_44_9=0
.ic qb_44_9=1.8
.ic q_45_9=0
.ic qb_45_9=1.8
.ic q_46_9=0
.ic qb_46_9=1.8
.ic q_47_9=0
.ic qb_47_9=1.8
.ic q_48_9=0
.ic qb_48_9=1.8
.ic q_49_9=0
.ic qb_49_9=1.8
.ic q_50_9=0
.ic qb_50_9=1.8
.ic q_51_9=0
.ic qb_51_9=1.8
.ic q_52_9=0
.ic qb_52_9=1.8
.ic q_53_9=0
.ic qb_53_9=1.8
.ic q_54_9=0
.ic qb_54_9=1.8
.ic q_55_9=0
.ic qb_55_9=1.8
.ic q_56_9=0
.ic qb_56_9=1.8
.ic q_57_9=0
.ic qb_57_9=1.8
.ic q_58_9=0
.ic qb_58_9=1.8
.ic q_59_9=0
.ic qb_59_9=1.8
.ic q_60_9=0
.ic qb_60_9=1.8
.ic q_61_9=0
.ic qb_61_9=1.8
.ic q_62_9=0
.ic qb_62_9=1.8
.ic q_63_9=0
.ic qb_63_9=1.8
.ic q_64_9=0
.ic qb_64_9=1.8
.ic q_65_9=0
.ic qb_65_9=1.8
.ic q_66_9=0
.ic qb_66_9=1.8
.ic q_67_9=0
.ic qb_67_9=1.8
.ic q_68_9=0
.ic qb_68_9=1.8
.ic q_69_9=0
.ic qb_69_9=1.8
.ic q_70_9=0
.ic qb_70_9=1.8
.ic q_71_9=0
.ic qb_71_9=1.8
.ic q_72_9=0
.ic qb_72_9=1.8
.ic q_73_9=0
.ic qb_73_9=1.8
.ic q_74_9=0
.ic qb_74_9=1.8
.ic q_75_9=0
.ic qb_75_9=1.8
.ic q_76_9=0
.ic qb_76_9=1.8
.ic q_77_9=0
.ic qb_77_9=1.8
.ic q_78_9=0
.ic qb_78_9=1.8
.ic q_79_9=0
.ic qb_79_9=1.8
.ic q_80_9=0
.ic qb_80_9=1.8
.ic q_81_9=0
.ic qb_81_9=1.8
.ic q_82_9=0
.ic qb_82_9=1.8
.ic q_83_9=0
.ic qb_83_9=1.8
.ic q_84_9=0
.ic qb_84_9=1.8
.ic q_85_9=0
.ic qb_85_9=1.8
.ic q_86_9=0
.ic qb_86_9=1.8
.ic q_87_9=0
.ic qb_87_9=1.8
.ic q_88_9=0
.ic qb_88_9=1.8
.ic q_89_9=0
.ic qb_89_9=1.8
.ic q_90_9=0
.ic qb_90_9=1.8
.ic q_91_9=0
.ic qb_91_9=1.8
.ic q_92_9=0
.ic qb_92_9=1.8
.ic q_93_9=0
.ic qb_93_9=1.8
.ic q_94_9=0
.ic qb_94_9=1.8
.ic q_95_9=0
.ic qb_95_9=1.8
.ic q_96_9=0
.ic qb_96_9=1.8
.ic q_97_9=0
.ic qb_97_9=1.8
.ic q_98_9=0
.ic qb_98_9=1.8
.ic q_99_9=0
.ic qb_99_9=1.8
.ic q_0_10=0
.ic qb_0_10=1.8
.ic q_1_10=0
.ic qb_1_10=1.8
.ic q_2_10=0
.ic qb_2_10=1.8
.ic q_3_10=0
.ic qb_3_10=1.8
.ic q_4_10=0
.ic qb_4_10=1.8
.ic q_5_10=0
.ic qb_5_10=1.8
.ic q_6_10=0
.ic qb_6_10=1.8
.ic q_7_10=0
.ic qb_7_10=1.8
.ic q_8_10=0
.ic qb_8_10=1.8
.ic q_9_10=0
.ic qb_9_10=1.8
.ic q_10_10=0
.ic qb_10_10=1.8
.ic q_11_10=0
.ic qb_11_10=1.8
.ic q_12_10=0
.ic qb_12_10=1.8
.ic q_13_10=0
.ic qb_13_10=1.8
.ic q_14_10=0
.ic qb_14_10=1.8
.ic q_15_10=0
.ic qb_15_10=1.8
.ic q_16_10=0
.ic qb_16_10=1.8
.ic q_17_10=0
.ic qb_17_10=1.8
.ic q_18_10=0
.ic qb_18_10=1.8
.ic q_19_10=0
.ic qb_19_10=1.8
.ic q_20_10=0
.ic qb_20_10=1.8
.ic q_21_10=0
.ic qb_21_10=1.8
.ic q_22_10=0
.ic qb_22_10=1.8
.ic q_23_10=0
.ic qb_23_10=1.8
.ic q_24_10=0
.ic qb_24_10=1.8
.ic q_25_10=0
.ic qb_25_10=1.8
.ic q_26_10=0
.ic qb_26_10=1.8
.ic q_27_10=0
.ic qb_27_10=1.8
.ic q_28_10=0
.ic qb_28_10=1.8
.ic q_29_10=0
.ic qb_29_10=1.8
.ic q_30_10=0
.ic qb_30_10=1.8
.ic q_31_10=0
.ic qb_31_10=1.8
.ic q_32_10=0
.ic qb_32_10=1.8
.ic q_33_10=0
.ic qb_33_10=1.8
.ic q_34_10=0
.ic qb_34_10=1.8
.ic q_35_10=0
.ic qb_35_10=1.8
.ic q_36_10=0
.ic qb_36_10=1.8
.ic q_37_10=0
.ic qb_37_10=1.8
.ic q_38_10=0
.ic qb_38_10=1.8
.ic q_39_10=0
.ic qb_39_10=1.8
.ic q_40_10=0
.ic qb_40_10=1.8
.ic q_41_10=0
.ic qb_41_10=1.8
.ic q_42_10=0
.ic qb_42_10=1.8
.ic q_43_10=0
.ic qb_43_10=1.8
.ic q_44_10=0
.ic qb_44_10=1.8
.ic q_45_10=0
.ic qb_45_10=1.8
.ic q_46_10=0
.ic qb_46_10=1.8
.ic q_47_10=0
.ic qb_47_10=1.8
.ic q_48_10=0
.ic qb_48_10=1.8
.ic q_49_10=0
.ic qb_49_10=1.8
.ic q_50_10=0
.ic qb_50_10=1.8
.ic q_51_10=0
.ic qb_51_10=1.8
.ic q_52_10=0
.ic qb_52_10=1.8
.ic q_53_10=0
.ic qb_53_10=1.8
.ic q_54_10=0
.ic qb_54_10=1.8
.ic q_55_10=0
.ic qb_55_10=1.8
.ic q_56_10=0
.ic qb_56_10=1.8
.ic q_57_10=0
.ic qb_57_10=1.8
.ic q_58_10=0
.ic qb_58_10=1.8
.ic q_59_10=0
.ic qb_59_10=1.8
.ic q_60_10=0
.ic qb_60_10=1.8
.ic q_61_10=0
.ic qb_61_10=1.8
.ic q_62_10=0
.ic qb_62_10=1.8
.ic q_63_10=0
.ic qb_63_10=1.8
.ic q_64_10=0
.ic qb_64_10=1.8
.ic q_65_10=0
.ic qb_65_10=1.8
.ic q_66_10=0
.ic qb_66_10=1.8
.ic q_67_10=0
.ic qb_67_10=1.8
.ic q_68_10=0
.ic qb_68_10=1.8
.ic q_69_10=0
.ic qb_69_10=1.8
.ic q_70_10=0
.ic qb_70_10=1.8
.ic q_71_10=0
.ic qb_71_10=1.8
.ic q_72_10=0
.ic qb_72_10=1.8
.ic q_73_10=0
.ic qb_73_10=1.8
.ic q_74_10=0
.ic qb_74_10=1.8
.ic q_75_10=0
.ic qb_75_10=1.8
.ic q_76_10=0
.ic qb_76_10=1.8
.ic q_77_10=0
.ic qb_77_10=1.8
.ic q_78_10=0
.ic qb_78_10=1.8
.ic q_79_10=0
.ic qb_79_10=1.8
.ic q_80_10=0
.ic qb_80_10=1.8
.ic q_81_10=0
.ic qb_81_10=1.8
.ic q_82_10=0
.ic qb_82_10=1.8
.ic q_83_10=0
.ic qb_83_10=1.8
.ic q_84_10=0
.ic qb_84_10=1.8
.ic q_85_10=0
.ic qb_85_10=1.8
.ic q_86_10=0
.ic qb_86_10=1.8
.ic q_87_10=0
.ic qb_87_10=1.8
.ic q_88_10=0
.ic qb_88_10=1.8
.ic q_89_10=0
.ic qb_89_10=1.8
.ic q_90_10=0
.ic qb_90_10=1.8
.ic q_91_10=0
.ic qb_91_10=1.8
.ic q_92_10=0
.ic qb_92_10=1.8
.ic q_93_10=0
.ic qb_93_10=1.8
.ic q_94_10=0
.ic qb_94_10=1.8
.ic q_95_10=0
.ic qb_95_10=1.8
.ic q_96_10=0
.ic qb_96_10=1.8
.ic q_97_10=0
.ic qb_97_10=1.8
.ic q_98_10=0
.ic qb_98_10=1.8
.ic q_99_10=0
.ic qb_99_10=1.8
.ic q_0_11=0
.ic qb_0_11=1.8
.ic q_1_11=0
.ic qb_1_11=1.8
.ic q_2_11=0
.ic qb_2_11=1.8
.ic q_3_11=0
.ic qb_3_11=1.8
.ic q_4_11=0
.ic qb_4_11=1.8
.ic q_5_11=0
.ic qb_5_11=1.8
.ic q_6_11=0
.ic qb_6_11=1.8
.ic q_7_11=0
.ic qb_7_11=1.8
.ic q_8_11=0
.ic qb_8_11=1.8
.ic q_9_11=0
.ic qb_9_11=1.8
.ic q_10_11=0
.ic qb_10_11=1.8
.ic q_11_11=0
.ic qb_11_11=1.8
.ic q_12_11=0
.ic qb_12_11=1.8
.ic q_13_11=0
.ic qb_13_11=1.8
.ic q_14_11=0
.ic qb_14_11=1.8
.ic q_15_11=0
.ic qb_15_11=1.8
.ic q_16_11=0
.ic qb_16_11=1.8
.ic q_17_11=0
.ic qb_17_11=1.8
.ic q_18_11=0
.ic qb_18_11=1.8
.ic q_19_11=0
.ic qb_19_11=1.8
.ic q_20_11=0
.ic qb_20_11=1.8
.ic q_21_11=0
.ic qb_21_11=1.8
.ic q_22_11=0
.ic qb_22_11=1.8
.ic q_23_11=0
.ic qb_23_11=1.8
.ic q_24_11=0
.ic qb_24_11=1.8
.ic q_25_11=0
.ic qb_25_11=1.8
.ic q_26_11=0
.ic qb_26_11=1.8
.ic q_27_11=0
.ic qb_27_11=1.8
.ic q_28_11=0
.ic qb_28_11=1.8
.ic q_29_11=0
.ic qb_29_11=1.8
.ic q_30_11=0
.ic qb_30_11=1.8
.ic q_31_11=0
.ic qb_31_11=1.8
.ic q_32_11=0
.ic qb_32_11=1.8
.ic q_33_11=0
.ic qb_33_11=1.8
.ic q_34_11=0
.ic qb_34_11=1.8
.ic q_35_11=0
.ic qb_35_11=1.8
.ic q_36_11=0
.ic qb_36_11=1.8
.ic q_37_11=0
.ic qb_37_11=1.8
.ic q_38_11=0
.ic qb_38_11=1.8
.ic q_39_11=0
.ic qb_39_11=1.8
.ic q_40_11=0
.ic qb_40_11=1.8
.ic q_41_11=0
.ic qb_41_11=1.8
.ic q_42_11=0
.ic qb_42_11=1.8
.ic q_43_11=0
.ic qb_43_11=1.8
.ic q_44_11=0
.ic qb_44_11=1.8
.ic q_45_11=0
.ic qb_45_11=1.8
.ic q_46_11=0
.ic qb_46_11=1.8
.ic q_47_11=0
.ic qb_47_11=1.8
.ic q_48_11=0
.ic qb_48_11=1.8
.ic q_49_11=0
.ic qb_49_11=1.8
.ic q_50_11=0
.ic qb_50_11=1.8
.ic q_51_11=0
.ic qb_51_11=1.8
.ic q_52_11=0
.ic qb_52_11=1.8
.ic q_53_11=0
.ic qb_53_11=1.8
.ic q_54_11=0
.ic qb_54_11=1.8
.ic q_55_11=0
.ic qb_55_11=1.8
.ic q_56_11=0
.ic qb_56_11=1.8
.ic q_57_11=0
.ic qb_57_11=1.8
.ic q_58_11=0
.ic qb_58_11=1.8
.ic q_59_11=0
.ic qb_59_11=1.8
.ic q_60_11=0
.ic qb_60_11=1.8
.ic q_61_11=0
.ic qb_61_11=1.8
.ic q_62_11=0
.ic qb_62_11=1.8
.ic q_63_11=0
.ic qb_63_11=1.8
.ic q_64_11=0
.ic qb_64_11=1.8
.ic q_65_11=0
.ic qb_65_11=1.8
.ic q_66_11=0
.ic qb_66_11=1.8
.ic q_67_11=0
.ic qb_67_11=1.8
.ic q_68_11=0
.ic qb_68_11=1.8
.ic q_69_11=0
.ic qb_69_11=1.8
.ic q_70_11=0
.ic qb_70_11=1.8
.ic q_71_11=0
.ic qb_71_11=1.8
.ic q_72_11=0
.ic qb_72_11=1.8
.ic q_73_11=0
.ic qb_73_11=1.8
.ic q_74_11=0
.ic qb_74_11=1.8
.ic q_75_11=0
.ic qb_75_11=1.8
.ic q_76_11=0
.ic qb_76_11=1.8
.ic q_77_11=0
.ic qb_77_11=1.8
.ic q_78_11=0
.ic qb_78_11=1.8
.ic q_79_11=0
.ic qb_79_11=1.8
.ic q_80_11=0
.ic qb_80_11=1.8
.ic q_81_11=0
.ic qb_81_11=1.8
.ic q_82_11=0
.ic qb_82_11=1.8
.ic q_83_11=0
.ic qb_83_11=1.8
.ic q_84_11=0
.ic qb_84_11=1.8
.ic q_85_11=0
.ic qb_85_11=1.8
.ic q_86_11=0
.ic qb_86_11=1.8
.ic q_87_11=0
.ic qb_87_11=1.8
.ic q_88_11=0
.ic qb_88_11=1.8
.ic q_89_11=0
.ic qb_89_11=1.8
.ic q_90_11=0
.ic qb_90_11=1.8
.ic q_91_11=0
.ic qb_91_11=1.8
.ic q_92_11=0
.ic qb_92_11=1.8
.ic q_93_11=0
.ic qb_93_11=1.8
.ic q_94_11=0
.ic qb_94_11=1.8
.ic q_95_11=0
.ic qb_95_11=1.8
.ic q_96_11=0
.ic qb_96_11=1.8
.ic q_97_11=0
.ic qb_97_11=1.8
.ic q_98_11=0
.ic qb_98_11=1.8
.ic q_99_11=0
.ic qb_99_11=1.8
.ic q_0_12=0
.ic qb_0_12=1.8
.ic q_1_12=0
.ic qb_1_12=1.8
.ic q_2_12=0
.ic qb_2_12=1.8
.ic q_3_12=0
.ic qb_3_12=1.8
.ic q_4_12=0
.ic qb_4_12=1.8
.ic q_5_12=0
.ic qb_5_12=1.8
.ic q_6_12=0
.ic qb_6_12=1.8
.ic q_7_12=0
.ic qb_7_12=1.8
.ic q_8_12=0
.ic qb_8_12=1.8
.ic q_9_12=0
.ic qb_9_12=1.8
.ic q_10_12=0
.ic qb_10_12=1.8
.ic q_11_12=0
.ic qb_11_12=1.8
.ic q_12_12=0
.ic qb_12_12=1.8
.ic q_13_12=0
.ic qb_13_12=1.8
.ic q_14_12=0
.ic qb_14_12=1.8
.ic q_15_12=0
.ic qb_15_12=1.8
.ic q_16_12=0
.ic qb_16_12=1.8
.ic q_17_12=0
.ic qb_17_12=1.8
.ic q_18_12=0
.ic qb_18_12=1.8
.ic q_19_12=0
.ic qb_19_12=1.8
.ic q_20_12=0
.ic qb_20_12=1.8
.ic q_21_12=0
.ic qb_21_12=1.8
.ic q_22_12=0
.ic qb_22_12=1.8
.ic q_23_12=0
.ic qb_23_12=1.8
.ic q_24_12=0
.ic qb_24_12=1.8
.ic q_25_12=0
.ic qb_25_12=1.8
.ic q_26_12=0
.ic qb_26_12=1.8
.ic q_27_12=0
.ic qb_27_12=1.8
.ic q_28_12=0
.ic qb_28_12=1.8
.ic q_29_12=0
.ic qb_29_12=1.8
.ic q_30_12=0
.ic qb_30_12=1.8
.ic q_31_12=0
.ic qb_31_12=1.8
.ic q_32_12=0
.ic qb_32_12=1.8
.ic q_33_12=0
.ic qb_33_12=1.8
.ic q_34_12=0
.ic qb_34_12=1.8
.ic q_35_12=0
.ic qb_35_12=1.8
.ic q_36_12=0
.ic qb_36_12=1.8
.ic q_37_12=0
.ic qb_37_12=1.8
.ic q_38_12=0
.ic qb_38_12=1.8
.ic q_39_12=0
.ic qb_39_12=1.8
.ic q_40_12=0
.ic qb_40_12=1.8
.ic q_41_12=0
.ic qb_41_12=1.8
.ic q_42_12=0
.ic qb_42_12=1.8
.ic q_43_12=0
.ic qb_43_12=1.8
.ic q_44_12=0
.ic qb_44_12=1.8
.ic q_45_12=0
.ic qb_45_12=1.8
.ic q_46_12=0
.ic qb_46_12=1.8
.ic q_47_12=0
.ic qb_47_12=1.8
.ic q_48_12=0
.ic qb_48_12=1.8
.ic q_49_12=0
.ic qb_49_12=1.8
.ic q_50_12=0
.ic qb_50_12=1.8
.ic q_51_12=0
.ic qb_51_12=1.8
.ic q_52_12=0
.ic qb_52_12=1.8
.ic q_53_12=0
.ic qb_53_12=1.8
.ic q_54_12=0
.ic qb_54_12=1.8
.ic q_55_12=0
.ic qb_55_12=1.8
.ic q_56_12=0
.ic qb_56_12=1.8
.ic q_57_12=0
.ic qb_57_12=1.8
.ic q_58_12=0
.ic qb_58_12=1.8
.ic q_59_12=0
.ic qb_59_12=1.8
.ic q_60_12=0
.ic qb_60_12=1.8
.ic q_61_12=0
.ic qb_61_12=1.8
.ic q_62_12=0
.ic qb_62_12=1.8
.ic q_63_12=0
.ic qb_63_12=1.8
.ic q_64_12=0
.ic qb_64_12=1.8
.ic q_65_12=0
.ic qb_65_12=1.8
.ic q_66_12=0
.ic qb_66_12=1.8
.ic q_67_12=0
.ic qb_67_12=1.8
.ic q_68_12=0
.ic qb_68_12=1.8
.ic q_69_12=0
.ic qb_69_12=1.8
.ic q_70_12=0
.ic qb_70_12=1.8
.ic q_71_12=0
.ic qb_71_12=1.8
.ic q_72_12=0
.ic qb_72_12=1.8
.ic q_73_12=0
.ic qb_73_12=1.8
.ic q_74_12=0
.ic qb_74_12=1.8
.ic q_75_12=0
.ic qb_75_12=1.8
.ic q_76_12=0
.ic qb_76_12=1.8
.ic q_77_12=0
.ic qb_77_12=1.8
.ic q_78_12=0
.ic qb_78_12=1.8
.ic q_79_12=0
.ic qb_79_12=1.8
.ic q_80_12=0
.ic qb_80_12=1.8
.ic q_81_12=0
.ic qb_81_12=1.8
.ic q_82_12=0
.ic qb_82_12=1.8
.ic q_83_12=0
.ic qb_83_12=1.8
.ic q_84_12=0
.ic qb_84_12=1.8
.ic q_85_12=0
.ic qb_85_12=1.8
.ic q_86_12=0
.ic qb_86_12=1.8
.ic q_87_12=0
.ic qb_87_12=1.8
.ic q_88_12=0
.ic qb_88_12=1.8
.ic q_89_12=0
.ic qb_89_12=1.8
.ic q_90_12=0
.ic qb_90_12=1.8
.ic q_91_12=0
.ic qb_91_12=1.8
.ic q_92_12=0
.ic qb_92_12=1.8
.ic q_93_12=0
.ic qb_93_12=1.8
.ic q_94_12=0
.ic qb_94_12=1.8
.ic q_95_12=0
.ic qb_95_12=1.8
.ic q_96_12=0
.ic qb_96_12=1.8
.ic q_97_12=0
.ic qb_97_12=1.8
.ic q_98_12=0
.ic qb_98_12=1.8
.ic q_99_12=0
.ic qb_99_12=1.8
.ic q_0_13=0
.ic qb_0_13=1.8
.ic q_1_13=0
.ic qb_1_13=1.8
.ic q_2_13=0
.ic qb_2_13=1.8
.ic q_3_13=0
.ic qb_3_13=1.8
.ic q_4_13=0
.ic qb_4_13=1.8
.ic q_5_13=0
.ic qb_5_13=1.8
.ic q_6_13=0
.ic qb_6_13=1.8
.ic q_7_13=0
.ic qb_7_13=1.8
.ic q_8_13=0
.ic qb_8_13=1.8
.ic q_9_13=0
.ic qb_9_13=1.8
.ic q_10_13=0
.ic qb_10_13=1.8
.ic q_11_13=0
.ic qb_11_13=1.8
.ic q_12_13=0
.ic qb_12_13=1.8
.ic q_13_13=0
.ic qb_13_13=1.8
.ic q_14_13=0
.ic qb_14_13=1.8
.ic q_15_13=0
.ic qb_15_13=1.8
.ic q_16_13=0
.ic qb_16_13=1.8
.ic q_17_13=0
.ic qb_17_13=1.8
.ic q_18_13=0
.ic qb_18_13=1.8
.ic q_19_13=0
.ic qb_19_13=1.8
.ic q_20_13=0
.ic qb_20_13=1.8
.ic q_21_13=0
.ic qb_21_13=1.8
.ic q_22_13=0
.ic qb_22_13=1.8
.ic q_23_13=0
.ic qb_23_13=1.8
.ic q_24_13=0
.ic qb_24_13=1.8
.ic q_25_13=0
.ic qb_25_13=1.8
.ic q_26_13=0
.ic qb_26_13=1.8
.ic q_27_13=0
.ic qb_27_13=1.8
.ic q_28_13=0
.ic qb_28_13=1.8
.ic q_29_13=0
.ic qb_29_13=1.8
.ic q_30_13=0
.ic qb_30_13=1.8
.ic q_31_13=0
.ic qb_31_13=1.8
.ic q_32_13=0
.ic qb_32_13=1.8
.ic q_33_13=0
.ic qb_33_13=1.8
.ic q_34_13=0
.ic qb_34_13=1.8
.ic q_35_13=0
.ic qb_35_13=1.8
.ic q_36_13=0
.ic qb_36_13=1.8
.ic q_37_13=0
.ic qb_37_13=1.8
.ic q_38_13=0
.ic qb_38_13=1.8
.ic q_39_13=0
.ic qb_39_13=1.8
.ic q_40_13=0
.ic qb_40_13=1.8
.ic q_41_13=0
.ic qb_41_13=1.8
.ic q_42_13=0
.ic qb_42_13=1.8
.ic q_43_13=0
.ic qb_43_13=1.8
.ic q_44_13=0
.ic qb_44_13=1.8
.ic q_45_13=0
.ic qb_45_13=1.8
.ic q_46_13=0
.ic qb_46_13=1.8
.ic q_47_13=0
.ic qb_47_13=1.8
.ic q_48_13=0
.ic qb_48_13=1.8
.ic q_49_13=0
.ic qb_49_13=1.8
.ic q_50_13=0
.ic qb_50_13=1.8
.ic q_51_13=0
.ic qb_51_13=1.8
.ic q_52_13=0
.ic qb_52_13=1.8
.ic q_53_13=0
.ic qb_53_13=1.8
.ic q_54_13=0
.ic qb_54_13=1.8
.ic q_55_13=0
.ic qb_55_13=1.8
.ic q_56_13=0
.ic qb_56_13=1.8
.ic q_57_13=0
.ic qb_57_13=1.8
.ic q_58_13=0
.ic qb_58_13=1.8
.ic q_59_13=0
.ic qb_59_13=1.8
.ic q_60_13=0
.ic qb_60_13=1.8
.ic q_61_13=0
.ic qb_61_13=1.8
.ic q_62_13=0
.ic qb_62_13=1.8
.ic q_63_13=0
.ic qb_63_13=1.8
.ic q_64_13=0
.ic qb_64_13=1.8
.ic q_65_13=0
.ic qb_65_13=1.8
.ic q_66_13=0
.ic qb_66_13=1.8
.ic q_67_13=0
.ic qb_67_13=1.8
.ic q_68_13=0
.ic qb_68_13=1.8
.ic q_69_13=0
.ic qb_69_13=1.8
.ic q_70_13=0
.ic qb_70_13=1.8
.ic q_71_13=0
.ic qb_71_13=1.8
.ic q_72_13=0
.ic qb_72_13=1.8
.ic q_73_13=0
.ic qb_73_13=1.8
.ic q_74_13=0
.ic qb_74_13=1.8
.ic q_75_13=0
.ic qb_75_13=1.8
.ic q_76_13=0
.ic qb_76_13=1.8
.ic q_77_13=0
.ic qb_77_13=1.8
.ic q_78_13=0
.ic qb_78_13=1.8
.ic q_79_13=0
.ic qb_79_13=1.8
.ic q_80_13=0
.ic qb_80_13=1.8
.ic q_81_13=0
.ic qb_81_13=1.8
.ic q_82_13=0
.ic qb_82_13=1.8
.ic q_83_13=0
.ic qb_83_13=1.8
.ic q_84_13=0
.ic qb_84_13=1.8
.ic q_85_13=0
.ic qb_85_13=1.8
.ic q_86_13=0
.ic qb_86_13=1.8
.ic q_87_13=0
.ic qb_87_13=1.8
.ic q_88_13=0
.ic qb_88_13=1.8
.ic q_89_13=0
.ic qb_89_13=1.8
.ic q_90_13=0
.ic qb_90_13=1.8
.ic q_91_13=0
.ic qb_91_13=1.8
.ic q_92_13=0
.ic qb_92_13=1.8
.ic q_93_13=0
.ic qb_93_13=1.8
.ic q_94_13=0
.ic qb_94_13=1.8
.ic q_95_13=0
.ic qb_95_13=1.8
.ic q_96_13=0
.ic qb_96_13=1.8
.ic q_97_13=0
.ic qb_97_13=1.8
.ic q_98_13=0
.ic qb_98_13=1.8
.ic q_99_13=0
.ic qb_99_13=1.8
.ic q_0_14=0
.ic qb_0_14=1.8
.ic q_1_14=0
.ic qb_1_14=1.8
.ic q_2_14=0
.ic qb_2_14=1.8
.ic q_3_14=0
.ic qb_3_14=1.8
.ic q_4_14=0
.ic qb_4_14=1.8
.ic q_5_14=0
.ic qb_5_14=1.8
.ic q_6_14=0
.ic qb_6_14=1.8
.ic q_7_14=0
.ic qb_7_14=1.8
.ic q_8_14=0
.ic qb_8_14=1.8
.ic q_9_14=0
.ic qb_9_14=1.8
.ic q_10_14=0
.ic qb_10_14=1.8
.ic q_11_14=0
.ic qb_11_14=1.8
.ic q_12_14=0
.ic qb_12_14=1.8
.ic q_13_14=0
.ic qb_13_14=1.8
.ic q_14_14=0
.ic qb_14_14=1.8
.ic q_15_14=0
.ic qb_15_14=1.8
.ic q_16_14=0
.ic qb_16_14=1.8
.ic q_17_14=0
.ic qb_17_14=1.8
.ic q_18_14=0
.ic qb_18_14=1.8
.ic q_19_14=0
.ic qb_19_14=1.8
.ic q_20_14=0
.ic qb_20_14=1.8
.ic q_21_14=0
.ic qb_21_14=1.8
.ic q_22_14=0
.ic qb_22_14=1.8
.ic q_23_14=0
.ic qb_23_14=1.8
.ic q_24_14=0
.ic qb_24_14=1.8
.ic q_25_14=0
.ic qb_25_14=1.8
.ic q_26_14=0
.ic qb_26_14=1.8
.ic q_27_14=0
.ic qb_27_14=1.8
.ic q_28_14=0
.ic qb_28_14=1.8
.ic q_29_14=0
.ic qb_29_14=1.8
.ic q_30_14=0
.ic qb_30_14=1.8
.ic q_31_14=0
.ic qb_31_14=1.8
.ic q_32_14=0
.ic qb_32_14=1.8
.ic q_33_14=0
.ic qb_33_14=1.8
.ic q_34_14=0
.ic qb_34_14=1.8
.ic q_35_14=0
.ic qb_35_14=1.8
.ic q_36_14=0
.ic qb_36_14=1.8
.ic q_37_14=0
.ic qb_37_14=1.8
.ic q_38_14=0
.ic qb_38_14=1.8
.ic q_39_14=0
.ic qb_39_14=1.8
.ic q_40_14=0
.ic qb_40_14=1.8
.ic q_41_14=0
.ic qb_41_14=1.8
.ic q_42_14=0
.ic qb_42_14=1.8
.ic q_43_14=0
.ic qb_43_14=1.8
.ic q_44_14=0
.ic qb_44_14=1.8
.ic q_45_14=0
.ic qb_45_14=1.8
.ic q_46_14=0
.ic qb_46_14=1.8
.ic q_47_14=0
.ic qb_47_14=1.8
.ic q_48_14=0
.ic qb_48_14=1.8
.ic q_49_14=0
.ic qb_49_14=1.8
.ic q_50_14=0
.ic qb_50_14=1.8
.ic q_51_14=0
.ic qb_51_14=1.8
.ic q_52_14=0
.ic qb_52_14=1.8
.ic q_53_14=0
.ic qb_53_14=1.8
.ic q_54_14=0
.ic qb_54_14=1.8
.ic q_55_14=0
.ic qb_55_14=1.8
.ic q_56_14=0
.ic qb_56_14=1.8
.ic q_57_14=0
.ic qb_57_14=1.8
.ic q_58_14=0
.ic qb_58_14=1.8
.ic q_59_14=0
.ic qb_59_14=1.8
.ic q_60_14=0
.ic qb_60_14=1.8
.ic q_61_14=0
.ic qb_61_14=1.8
.ic q_62_14=0
.ic qb_62_14=1.8
.ic q_63_14=0
.ic qb_63_14=1.8
.ic q_64_14=0
.ic qb_64_14=1.8
.ic q_65_14=0
.ic qb_65_14=1.8
.ic q_66_14=0
.ic qb_66_14=1.8
.ic q_67_14=0
.ic qb_67_14=1.8
.ic q_68_14=0
.ic qb_68_14=1.8
.ic q_69_14=0
.ic qb_69_14=1.8
.ic q_70_14=0
.ic qb_70_14=1.8
.ic q_71_14=0
.ic qb_71_14=1.8
.ic q_72_14=0
.ic qb_72_14=1.8
.ic q_73_14=0
.ic qb_73_14=1.8
.ic q_74_14=0
.ic qb_74_14=1.8
.ic q_75_14=0
.ic qb_75_14=1.8
.ic q_76_14=0
.ic qb_76_14=1.8
.ic q_77_14=0
.ic qb_77_14=1.8
.ic q_78_14=0
.ic qb_78_14=1.8
.ic q_79_14=0
.ic qb_79_14=1.8
.ic q_80_14=0
.ic qb_80_14=1.8
.ic q_81_14=0
.ic qb_81_14=1.8
.ic q_82_14=0
.ic qb_82_14=1.8
.ic q_83_14=0
.ic qb_83_14=1.8
.ic q_84_14=0
.ic qb_84_14=1.8
.ic q_85_14=0
.ic qb_85_14=1.8
.ic q_86_14=0
.ic qb_86_14=1.8
.ic q_87_14=0
.ic qb_87_14=1.8
.ic q_88_14=0
.ic qb_88_14=1.8
.ic q_89_14=0
.ic qb_89_14=1.8
.ic q_90_14=0
.ic qb_90_14=1.8
.ic q_91_14=0
.ic qb_91_14=1.8
.ic q_92_14=0
.ic qb_92_14=1.8
.ic q_93_14=0
.ic qb_93_14=1.8
.ic q_94_14=0
.ic qb_94_14=1.8
.ic q_95_14=0
.ic qb_95_14=1.8
.ic q_96_14=0
.ic qb_96_14=1.8
.ic q_97_14=0
.ic qb_97_14=1.8
.ic q_98_14=0
.ic qb_98_14=1.8
.ic q_99_14=0
.ic qb_99_14=1.8
.ic q_0_15=0
.ic qb_0_15=1.8
.ic q_1_15=0
.ic qb_1_15=1.8
.ic q_2_15=0
.ic qb_2_15=1.8
.ic q_3_15=0
.ic qb_3_15=1.8
.ic q_4_15=0
.ic qb_4_15=1.8
.ic q_5_15=0
.ic qb_5_15=1.8
.ic q_6_15=0
.ic qb_6_15=1.8
.ic q_7_15=0
.ic qb_7_15=1.8
.ic q_8_15=0
.ic qb_8_15=1.8
.ic q_9_15=0
.ic qb_9_15=1.8
.ic q_10_15=0
.ic qb_10_15=1.8
.ic q_11_15=0
.ic qb_11_15=1.8
.ic q_12_15=0
.ic qb_12_15=1.8
.ic q_13_15=0
.ic qb_13_15=1.8
.ic q_14_15=0
.ic qb_14_15=1.8
.ic q_15_15=0
.ic qb_15_15=1.8
.ic q_16_15=0
.ic qb_16_15=1.8
.ic q_17_15=0
.ic qb_17_15=1.8
.ic q_18_15=0
.ic qb_18_15=1.8
.ic q_19_15=0
.ic qb_19_15=1.8
.ic q_20_15=0
.ic qb_20_15=1.8
.ic q_21_15=0
.ic qb_21_15=1.8
.ic q_22_15=0
.ic qb_22_15=1.8
.ic q_23_15=0
.ic qb_23_15=1.8
.ic q_24_15=0
.ic qb_24_15=1.8
.ic q_25_15=0
.ic qb_25_15=1.8
.ic q_26_15=0
.ic qb_26_15=1.8
.ic q_27_15=0
.ic qb_27_15=1.8
.ic q_28_15=0
.ic qb_28_15=1.8
.ic q_29_15=0
.ic qb_29_15=1.8
.ic q_30_15=0
.ic qb_30_15=1.8
.ic q_31_15=0
.ic qb_31_15=1.8
.ic q_32_15=0
.ic qb_32_15=1.8
.ic q_33_15=0
.ic qb_33_15=1.8
.ic q_34_15=0
.ic qb_34_15=1.8
.ic q_35_15=0
.ic qb_35_15=1.8
.ic q_36_15=0
.ic qb_36_15=1.8
.ic q_37_15=0
.ic qb_37_15=1.8
.ic q_38_15=0
.ic qb_38_15=1.8
.ic q_39_15=0
.ic qb_39_15=1.8
.ic q_40_15=0
.ic qb_40_15=1.8
.ic q_41_15=0
.ic qb_41_15=1.8
.ic q_42_15=0
.ic qb_42_15=1.8
.ic q_43_15=0
.ic qb_43_15=1.8
.ic q_44_15=0
.ic qb_44_15=1.8
.ic q_45_15=0
.ic qb_45_15=1.8
.ic q_46_15=0
.ic qb_46_15=1.8
.ic q_47_15=0
.ic qb_47_15=1.8
.ic q_48_15=0
.ic qb_48_15=1.8
.ic q_49_15=0
.ic qb_49_15=1.8
.ic q_50_15=0
.ic qb_50_15=1.8
.ic q_51_15=0
.ic qb_51_15=1.8
.ic q_52_15=0
.ic qb_52_15=1.8
.ic q_53_15=0
.ic qb_53_15=1.8
.ic q_54_15=0
.ic qb_54_15=1.8
.ic q_55_15=0
.ic qb_55_15=1.8
.ic q_56_15=0
.ic qb_56_15=1.8
.ic q_57_15=0
.ic qb_57_15=1.8
.ic q_58_15=0
.ic qb_58_15=1.8
.ic q_59_15=0
.ic qb_59_15=1.8
.ic q_60_15=0
.ic qb_60_15=1.8
.ic q_61_15=0
.ic qb_61_15=1.8
.ic q_62_15=0
.ic qb_62_15=1.8
.ic q_63_15=0
.ic qb_63_15=1.8
.ic q_64_15=0
.ic qb_64_15=1.8
.ic q_65_15=0
.ic qb_65_15=1.8
.ic q_66_15=0
.ic qb_66_15=1.8
.ic q_67_15=0
.ic qb_67_15=1.8
.ic q_68_15=0
.ic qb_68_15=1.8
.ic q_69_15=0
.ic qb_69_15=1.8
.ic q_70_15=0
.ic qb_70_15=1.8
.ic q_71_15=0
.ic qb_71_15=1.8
.ic q_72_15=0
.ic qb_72_15=1.8
.ic q_73_15=0
.ic qb_73_15=1.8
.ic q_74_15=0
.ic qb_74_15=1.8
.ic q_75_15=0
.ic qb_75_15=1.8
.ic q_76_15=0
.ic qb_76_15=1.8
.ic q_77_15=0
.ic qb_77_15=1.8
.ic q_78_15=0
.ic qb_78_15=1.8
.ic q_79_15=0
.ic qb_79_15=1.8
.ic q_80_15=0
.ic qb_80_15=1.8
.ic q_81_15=0
.ic qb_81_15=1.8
.ic q_82_15=0
.ic qb_82_15=1.8
.ic q_83_15=0
.ic qb_83_15=1.8
.ic q_84_15=0
.ic qb_84_15=1.8
.ic q_85_15=0
.ic qb_85_15=1.8
.ic q_86_15=0
.ic qb_86_15=1.8
.ic q_87_15=0
.ic qb_87_15=1.8
.ic q_88_15=0
.ic qb_88_15=1.8
.ic q_89_15=0
.ic qb_89_15=1.8
.ic q_90_15=0
.ic qb_90_15=1.8
.ic q_91_15=0
.ic qb_91_15=1.8
.ic q_92_15=0
.ic qb_92_15=1.8
.ic q_93_15=0
.ic qb_93_15=1.8
.ic q_94_15=0
.ic qb_94_15=1.8
.ic q_95_15=0
.ic qb_95_15=1.8
.ic q_96_15=0
.ic qb_96_15=1.8
.ic q_97_15=0
.ic qb_97_15=1.8
.ic q_98_15=0
.ic qb_98_15=1.8
.ic q_99_15=0
.ic qb_99_15=1.8
.ic q_0_16=0
.ic qb_0_16=1.8
.ic q_1_16=0
.ic qb_1_16=1.8
.ic q_2_16=0
.ic qb_2_16=1.8
.ic q_3_16=0
.ic qb_3_16=1.8
.ic q_4_16=0
.ic qb_4_16=1.8
.ic q_5_16=0
.ic qb_5_16=1.8
.ic q_6_16=0
.ic qb_6_16=1.8
.ic q_7_16=0
.ic qb_7_16=1.8
.ic q_8_16=0
.ic qb_8_16=1.8
.ic q_9_16=0
.ic qb_9_16=1.8
.ic q_10_16=0
.ic qb_10_16=1.8
.ic q_11_16=0
.ic qb_11_16=1.8
.ic q_12_16=0
.ic qb_12_16=1.8
.ic q_13_16=0
.ic qb_13_16=1.8
.ic q_14_16=0
.ic qb_14_16=1.8
.ic q_15_16=0
.ic qb_15_16=1.8
.ic q_16_16=0
.ic qb_16_16=1.8
.ic q_17_16=0
.ic qb_17_16=1.8
.ic q_18_16=0
.ic qb_18_16=1.8
.ic q_19_16=0
.ic qb_19_16=1.8
.ic q_20_16=0
.ic qb_20_16=1.8
.ic q_21_16=0
.ic qb_21_16=1.8
.ic q_22_16=0
.ic qb_22_16=1.8
.ic q_23_16=0
.ic qb_23_16=1.8
.ic q_24_16=0
.ic qb_24_16=1.8
.ic q_25_16=0
.ic qb_25_16=1.8
.ic q_26_16=0
.ic qb_26_16=1.8
.ic q_27_16=0
.ic qb_27_16=1.8
.ic q_28_16=0
.ic qb_28_16=1.8
.ic q_29_16=0
.ic qb_29_16=1.8
.ic q_30_16=0
.ic qb_30_16=1.8
.ic q_31_16=0
.ic qb_31_16=1.8
.ic q_32_16=0
.ic qb_32_16=1.8
.ic q_33_16=0
.ic qb_33_16=1.8
.ic q_34_16=0
.ic qb_34_16=1.8
.ic q_35_16=0
.ic qb_35_16=1.8
.ic q_36_16=0
.ic qb_36_16=1.8
.ic q_37_16=0
.ic qb_37_16=1.8
.ic q_38_16=0
.ic qb_38_16=1.8
.ic q_39_16=0
.ic qb_39_16=1.8
.ic q_40_16=0
.ic qb_40_16=1.8
.ic q_41_16=0
.ic qb_41_16=1.8
.ic q_42_16=0
.ic qb_42_16=1.8
.ic q_43_16=0
.ic qb_43_16=1.8
.ic q_44_16=0
.ic qb_44_16=1.8
.ic q_45_16=0
.ic qb_45_16=1.8
.ic q_46_16=0
.ic qb_46_16=1.8
.ic q_47_16=0
.ic qb_47_16=1.8
.ic q_48_16=0
.ic qb_48_16=1.8
.ic q_49_16=0
.ic qb_49_16=1.8
.ic q_50_16=0
.ic qb_50_16=1.8
.ic q_51_16=0
.ic qb_51_16=1.8
.ic q_52_16=0
.ic qb_52_16=1.8
.ic q_53_16=0
.ic qb_53_16=1.8
.ic q_54_16=0
.ic qb_54_16=1.8
.ic q_55_16=0
.ic qb_55_16=1.8
.ic q_56_16=0
.ic qb_56_16=1.8
.ic q_57_16=0
.ic qb_57_16=1.8
.ic q_58_16=0
.ic qb_58_16=1.8
.ic q_59_16=0
.ic qb_59_16=1.8
.ic q_60_16=0
.ic qb_60_16=1.8
.ic q_61_16=0
.ic qb_61_16=1.8
.ic q_62_16=0
.ic qb_62_16=1.8
.ic q_63_16=0
.ic qb_63_16=1.8
.ic q_64_16=0
.ic qb_64_16=1.8
.ic q_65_16=0
.ic qb_65_16=1.8
.ic q_66_16=0
.ic qb_66_16=1.8
.ic q_67_16=0
.ic qb_67_16=1.8
.ic q_68_16=0
.ic qb_68_16=1.8
.ic q_69_16=0
.ic qb_69_16=1.8
.ic q_70_16=0
.ic qb_70_16=1.8
.ic q_71_16=0
.ic qb_71_16=1.8
.ic q_72_16=0
.ic qb_72_16=1.8
.ic q_73_16=0
.ic qb_73_16=1.8
.ic q_74_16=0
.ic qb_74_16=1.8
.ic q_75_16=0
.ic qb_75_16=1.8
.ic q_76_16=0
.ic qb_76_16=1.8
.ic q_77_16=0
.ic qb_77_16=1.8
.ic q_78_16=0
.ic qb_78_16=1.8
.ic q_79_16=0
.ic qb_79_16=1.8
.ic q_80_16=0
.ic qb_80_16=1.8
.ic q_81_16=0
.ic qb_81_16=1.8
.ic q_82_16=0
.ic qb_82_16=1.8
.ic q_83_16=0
.ic qb_83_16=1.8
.ic q_84_16=0
.ic qb_84_16=1.8
.ic q_85_16=0
.ic qb_85_16=1.8
.ic q_86_16=0
.ic qb_86_16=1.8
.ic q_87_16=0
.ic qb_87_16=1.8
.ic q_88_16=0
.ic qb_88_16=1.8
.ic q_89_16=0
.ic qb_89_16=1.8
.ic q_90_16=0
.ic qb_90_16=1.8
.ic q_91_16=0
.ic qb_91_16=1.8
.ic q_92_16=0
.ic qb_92_16=1.8
.ic q_93_16=0
.ic qb_93_16=1.8
.ic q_94_16=0
.ic qb_94_16=1.8
.ic q_95_16=0
.ic qb_95_16=1.8
.ic q_96_16=0
.ic qb_96_16=1.8
.ic q_97_16=0
.ic qb_97_16=1.8
.ic q_98_16=0
.ic qb_98_16=1.8
.ic q_99_16=0
.ic qb_99_16=1.8
.ic q_0_17=0
.ic qb_0_17=1.8
.ic q_1_17=0
.ic qb_1_17=1.8
.ic q_2_17=0
.ic qb_2_17=1.8
.ic q_3_17=0
.ic qb_3_17=1.8
.ic q_4_17=0
.ic qb_4_17=1.8
.ic q_5_17=0
.ic qb_5_17=1.8
.ic q_6_17=0
.ic qb_6_17=1.8
.ic q_7_17=0
.ic qb_7_17=1.8
.ic q_8_17=0
.ic qb_8_17=1.8
.ic q_9_17=0
.ic qb_9_17=1.8
.ic q_10_17=0
.ic qb_10_17=1.8
.ic q_11_17=0
.ic qb_11_17=1.8
.ic q_12_17=0
.ic qb_12_17=1.8
.ic q_13_17=0
.ic qb_13_17=1.8
.ic q_14_17=0
.ic qb_14_17=1.8
.ic q_15_17=0
.ic qb_15_17=1.8
.ic q_16_17=0
.ic qb_16_17=1.8
.ic q_17_17=0
.ic qb_17_17=1.8
.ic q_18_17=0
.ic qb_18_17=1.8
.ic q_19_17=0
.ic qb_19_17=1.8
.ic q_20_17=0
.ic qb_20_17=1.8
.ic q_21_17=0
.ic qb_21_17=1.8
.ic q_22_17=0
.ic qb_22_17=1.8
.ic q_23_17=0
.ic qb_23_17=1.8
.ic q_24_17=0
.ic qb_24_17=1.8
.ic q_25_17=0
.ic qb_25_17=1.8
.ic q_26_17=0
.ic qb_26_17=1.8
.ic q_27_17=0
.ic qb_27_17=1.8
.ic q_28_17=0
.ic qb_28_17=1.8
.ic q_29_17=0
.ic qb_29_17=1.8
.ic q_30_17=0
.ic qb_30_17=1.8
.ic q_31_17=0
.ic qb_31_17=1.8
.ic q_32_17=0
.ic qb_32_17=1.8
.ic q_33_17=0
.ic qb_33_17=1.8
.ic q_34_17=0
.ic qb_34_17=1.8
.ic q_35_17=0
.ic qb_35_17=1.8
.ic q_36_17=0
.ic qb_36_17=1.8
.ic q_37_17=0
.ic qb_37_17=1.8
.ic q_38_17=0
.ic qb_38_17=1.8
.ic q_39_17=0
.ic qb_39_17=1.8
.ic q_40_17=0
.ic qb_40_17=1.8
.ic q_41_17=0
.ic qb_41_17=1.8
.ic q_42_17=0
.ic qb_42_17=1.8
.ic q_43_17=0
.ic qb_43_17=1.8
.ic q_44_17=0
.ic qb_44_17=1.8
.ic q_45_17=0
.ic qb_45_17=1.8
.ic q_46_17=0
.ic qb_46_17=1.8
.ic q_47_17=0
.ic qb_47_17=1.8
.ic q_48_17=0
.ic qb_48_17=1.8
.ic q_49_17=0
.ic qb_49_17=1.8
.ic q_50_17=0
.ic qb_50_17=1.8
.ic q_51_17=0
.ic qb_51_17=1.8
.ic q_52_17=0
.ic qb_52_17=1.8
.ic q_53_17=0
.ic qb_53_17=1.8
.ic q_54_17=0
.ic qb_54_17=1.8
.ic q_55_17=0
.ic qb_55_17=1.8
.ic q_56_17=0
.ic qb_56_17=1.8
.ic q_57_17=0
.ic qb_57_17=1.8
.ic q_58_17=0
.ic qb_58_17=1.8
.ic q_59_17=0
.ic qb_59_17=1.8
.ic q_60_17=0
.ic qb_60_17=1.8
.ic q_61_17=0
.ic qb_61_17=1.8
.ic q_62_17=0
.ic qb_62_17=1.8
.ic q_63_17=0
.ic qb_63_17=1.8
.ic q_64_17=0
.ic qb_64_17=1.8
.ic q_65_17=0
.ic qb_65_17=1.8
.ic q_66_17=0
.ic qb_66_17=1.8
.ic q_67_17=0
.ic qb_67_17=1.8
.ic q_68_17=0
.ic qb_68_17=1.8
.ic q_69_17=0
.ic qb_69_17=1.8
.ic q_70_17=0
.ic qb_70_17=1.8
.ic q_71_17=0
.ic qb_71_17=1.8
.ic q_72_17=0
.ic qb_72_17=1.8
.ic q_73_17=0
.ic qb_73_17=1.8
.ic q_74_17=0
.ic qb_74_17=1.8
.ic q_75_17=0
.ic qb_75_17=1.8
.ic q_76_17=0
.ic qb_76_17=1.8
.ic q_77_17=0
.ic qb_77_17=1.8
.ic q_78_17=0
.ic qb_78_17=1.8
.ic q_79_17=0
.ic qb_79_17=1.8
.ic q_80_17=0
.ic qb_80_17=1.8
.ic q_81_17=0
.ic qb_81_17=1.8
.ic q_82_17=0
.ic qb_82_17=1.8
.ic q_83_17=0
.ic qb_83_17=1.8
.ic q_84_17=0
.ic qb_84_17=1.8
.ic q_85_17=0
.ic qb_85_17=1.8
.ic q_86_17=0
.ic qb_86_17=1.8
.ic q_87_17=0
.ic qb_87_17=1.8
.ic q_88_17=0
.ic qb_88_17=1.8
.ic q_89_17=0
.ic qb_89_17=1.8
.ic q_90_17=0
.ic qb_90_17=1.8
.ic q_91_17=0
.ic qb_91_17=1.8
.ic q_92_17=0
.ic qb_92_17=1.8
.ic q_93_17=0
.ic qb_93_17=1.8
.ic q_94_17=0
.ic qb_94_17=1.8
.ic q_95_17=0
.ic qb_95_17=1.8
.ic q_96_17=0
.ic qb_96_17=1.8
.ic q_97_17=0
.ic qb_97_17=1.8
.ic q_98_17=0
.ic qb_98_17=1.8
.ic q_99_17=0
.ic qb_99_17=1.8
.ic q_0_18=0
.ic qb_0_18=1.8
.ic q_1_18=0
.ic qb_1_18=1.8
.ic q_2_18=0
.ic qb_2_18=1.8
.ic q_3_18=0
.ic qb_3_18=1.8
.ic q_4_18=0
.ic qb_4_18=1.8
.ic q_5_18=0
.ic qb_5_18=1.8
.ic q_6_18=0
.ic qb_6_18=1.8
.ic q_7_18=0
.ic qb_7_18=1.8
.ic q_8_18=0
.ic qb_8_18=1.8
.ic q_9_18=0
.ic qb_9_18=1.8
.ic q_10_18=0
.ic qb_10_18=1.8
.ic q_11_18=0
.ic qb_11_18=1.8
.ic q_12_18=0
.ic qb_12_18=1.8
.ic q_13_18=0
.ic qb_13_18=1.8
.ic q_14_18=0
.ic qb_14_18=1.8
.ic q_15_18=0
.ic qb_15_18=1.8
.ic q_16_18=0
.ic qb_16_18=1.8
.ic q_17_18=0
.ic qb_17_18=1.8
.ic q_18_18=0
.ic qb_18_18=1.8
.ic q_19_18=0
.ic qb_19_18=1.8
.ic q_20_18=0
.ic qb_20_18=1.8
.ic q_21_18=0
.ic qb_21_18=1.8
.ic q_22_18=0
.ic qb_22_18=1.8
.ic q_23_18=0
.ic qb_23_18=1.8
.ic q_24_18=0
.ic qb_24_18=1.8
.ic q_25_18=0
.ic qb_25_18=1.8
.ic q_26_18=0
.ic qb_26_18=1.8
.ic q_27_18=0
.ic qb_27_18=1.8
.ic q_28_18=0
.ic qb_28_18=1.8
.ic q_29_18=0
.ic qb_29_18=1.8
.ic q_30_18=0
.ic qb_30_18=1.8
.ic q_31_18=0
.ic qb_31_18=1.8
.ic q_32_18=0
.ic qb_32_18=1.8
.ic q_33_18=0
.ic qb_33_18=1.8
.ic q_34_18=0
.ic qb_34_18=1.8
.ic q_35_18=0
.ic qb_35_18=1.8
.ic q_36_18=0
.ic qb_36_18=1.8
.ic q_37_18=0
.ic qb_37_18=1.8
.ic q_38_18=0
.ic qb_38_18=1.8
.ic q_39_18=0
.ic qb_39_18=1.8
.ic q_40_18=0
.ic qb_40_18=1.8
.ic q_41_18=0
.ic qb_41_18=1.8
.ic q_42_18=0
.ic qb_42_18=1.8
.ic q_43_18=0
.ic qb_43_18=1.8
.ic q_44_18=0
.ic qb_44_18=1.8
.ic q_45_18=0
.ic qb_45_18=1.8
.ic q_46_18=0
.ic qb_46_18=1.8
.ic q_47_18=0
.ic qb_47_18=1.8
.ic q_48_18=0
.ic qb_48_18=1.8
.ic q_49_18=0
.ic qb_49_18=1.8
.ic q_50_18=0
.ic qb_50_18=1.8
.ic q_51_18=0
.ic qb_51_18=1.8
.ic q_52_18=0
.ic qb_52_18=1.8
.ic q_53_18=0
.ic qb_53_18=1.8
.ic q_54_18=0
.ic qb_54_18=1.8
.ic q_55_18=0
.ic qb_55_18=1.8
.ic q_56_18=0
.ic qb_56_18=1.8
.ic q_57_18=0
.ic qb_57_18=1.8
.ic q_58_18=0
.ic qb_58_18=1.8
.ic q_59_18=0
.ic qb_59_18=1.8
.ic q_60_18=0
.ic qb_60_18=1.8
.ic q_61_18=0
.ic qb_61_18=1.8
.ic q_62_18=0
.ic qb_62_18=1.8
.ic q_63_18=0
.ic qb_63_18=1.8
.ic q_64_18=0
.ic qb_64_18=1.8
.ic q_65_18=0
.ic qb_65_18=1.8
.ic q_66_18=0
.ic qb_66_18=1.8
.ic q_67_18=0
.ic qb_67_18=1.8
.ic q_68_18=0
.ic qb_68_18=1.8
.ic q_69_18=0
.ic qb_69_18=1.8
.ic q_70_18=0
.ic qb_70_18=1.8
.ic q_71_18=0
.ic qb_71_18=1.8
.ic q_72_18=0
.ic qb_72_18=1.8
.ic q_73_18=0
.ic qb_73_18=1.8
.ic q_74_18=0
.ic qb_74_18=1.8
.ic q_75_18=0
.ic qb_75_18=1.8
.ic q_76_18=0
.ic qb_76_18=1.8
.ic q_77_18=0
.ic qb_77_18=1.8
.ic q_78_18=0
.ic qb_78_18=1.8
.ic q_79_18=0
.ic qb_79_18=1.8
.ic q_80_18=0
.ic qb_80_18=1.8
.ic q_81_18=0
.ic qb_81_18=1.8
.ic q_82_18=0
.ic qb_82_18=1.8
.ic q_83_18=0
.ic qb_83_18=1.8
.ic q_84_18=0
.ic qb_84_18=1.8
.ic q_85_18=0
.ic qb_85_18=1.8
.ic q_86_18=0
.ic qb_86_18=1.8
.ic q_87_18=0
.ic qb_87_18=1.8
.ic q_88_18=0
.ic qb_88_18=1.8
.ic q_89_18=0
.ic qb_89_18=1.8
.ic q_90_18=0
.ic qb_90_18=1.8
.ic q_91_18=0
.ic qb_91_18=1.8
.ic q_92_18=0
.ic qb_92_18=1.8
.ic q_93_18=0
.ic qb_93_18=1.8
.ic q_94_18=0
.ic qb_94_18=1.8
.ic q_95_18=0
.ic qb_95_18=1.8
.ic q_96_18=0
.ic qb_96_18=1.8
.ic q_97_18=0
.ic qb_97_18=1.8
.ic q_98_18=0
.ic qb_98_18=1.8
.ic q_99_18=0
.ic qb_99_18=1.8
.ic q_0_19=0
.ic qb_0_19=1.8
.ic q_1_19=0
.ic qb_1_19=1.8
.ic q_2_19=0
.ic qb_2_19=1.8
.ic q_3_19=0
.ic qb_3_19=1.8
.ic q_4_19=0
.ic qb_4_19=1.8
.ic q_5_19=0
.ic qb_5_19=1.8
.ic q_6_19=0
.ic qb_6_19=1.8
.ic q_7_19=0
.ic qb_7_19=1.8
.ic q_8_19=0
.ic qb_8_19=1.8
.ic q_9_19=0
.ic qb_9_19=1.8
.ic q_10_19=0
.ic qb_10_19=1.8
.ic q_11_19=0
.ic qb_11_19=1.8
.ic q_12_19=0
.ic qb_12_19=1.8
.ic q_13_19=0
.ic qb_13_19=1.8
.ic q_14_19=0
.ic qb_14_19=1.8
.ic q_15_19=0
.ic qb_15_19=1.8
.ic q_16_19=0
.ic qb_16_19=1.8
.ic q_17_19=0
.ic qb_17_19=1.8
.ic q_18_19=0
.ic qb_18_19=1.8
.ic q_19_19=0
.ic qb_19_19=1.8
.ic q_20_19=0
.ic qb_20_19=1.8
.ic q_21_19=0
.ic qb_21_19=1.8
.ic q_22_19=0
.ic qb_22_19=1.8
.ic q_23_19=0
.ic qb_23_19=1.8
.ic q_24_19=0
.ic qb_24_19=1.8
.ic q_25_19=0
.ic qb_25_19=1.8
.ic q_26_19=0
.ic qb_26_19=1.8
.ic q_27_19=0
.ic qb_27_19=1.8
.ic q_28_19=0
.ic qb_28_19=1.8
.ic q_29_19=0
.ic qb_29_19=1.8
.ic q_30_19=0
.ic qb_30_19=1.8
.ic q_31_19=0
.ic qb_31_19=1.8
.ic q_32_19=0
.ic qb_32_19=1.8
.ic q_33_19=0
.ic qb_33_19=1.8
.ic q_34_19=0
.ic qb_34_19=1.8
.ic q_35_19=0
.ic qb_35_19=1.8
.ic q_36_19=0
.ic qb_36_19=1.8
.ic q_37_19=0
.ic qb_37_19=1.8
.ic q_38_19=0
.ic qb_38_19=1.8
.ic q_39_19=0
.ic qb_39_19=1.8
.ic q_40_19=0
.ic qb_40_19=1.8
.ic q_41_19=0
.ic qb_41_19=1.8
.ic q_42_19=0
.ic qb_42_19=1.8
.ic q_43_19=0
.ic qb_43_19=1.8
.ic q_44_19=0
.ic qb_44_19=1.8
.ic q_45_19=0
.ic qb_45_19=1.8
.ic q_46_19=0
.ic qb_46_19=1.8
.ic q_47_19=0
.ic qb_47_19=1.8
.ic q_48_19=0
.ic qb_48_19=1.8
.ic q_49_19=0
.ic qb_49_19=1.8
.ic q_50_19=0
.ic qb_50_19=1.8
.ic q_51_19=0
.ic qb_51_19=1.8
.ic q_52_19=0
.ic qb_52_19=1.8
.ic q_53_19=0
.ic qb_53_19=1.8
.ic q_54_19=0
.ic qb_54_19=1.8
.ic q_55_19=0
.ic qb_55_19=1.8
.ic q_56_19=0
.ic qb_56_19=1.8
.ic q_57_19=0
.ic qb_57_19=1.8
.ic q_58_19=0
.ic qb_58_19=1.8
.ic q_59_19=0
.ic qb_59_19=1.8
.ic q_60_19=0
.ic qb_60_19=1.8
.ic q_61_19=0
.ic qb_61_19=1.8
.ic q_62_19=0
.ic qb_62_19=1.8
.ic q_63_19=0
.ic qb_63_19=1.8
.ic q_64_19=0
.ic qb_64_19=1.8
.ic q_65_19=0
.ic qb_65_19=1.8
.ic q_66_19=0
.ic qb_66_19=1.8
.ic q_67_19=0
.ic qb_67_19=1.8
.ic q_68_19=0
.ic qb_68_19=1.8
.ic q_69_19=0
.ic qb_69_19=1.8
.ic q_70_19=0
.ic qb_70_19=1.8
.ic q_71_19=0
.ic qb_71_19=1.8
.ic q_72_19=0
.ic qb_72_19=1.8
.ic q_73_19=0
.ic qb_73_19=1.8
.ic q_74_19=0
.ic qb_74_19=1.8
.ic q_75_19=0
.ic qb_75_19=1.8
.ic q_76_19=0
.ic qb_76_19=1.8
.ic q_77_19=0
.ic qb_77_19=1.8
.ic q_78_19=0
.ic qb_78_19=1.8
.ic q_79_19=0
.ic qb_79_19=1.8
.ic q_80_19=0
.ic qb_80_19=1.8
.ic q_81_19=0
.ic qb_81_19=1.8
.ic q_82_19=0
.ic qb_82_19=1.8
.ic q_83_19=0
.ic qb_83_19=1.8
.ic q_84_19=0
.ic qb_84_19=1.8
.ic q_85_19=0
.ic qb_85_19=1.8
.ic q_86_19=0
.ic qb_86_19=1.8
.ic q_87_19=0
.ic qb_87_19=1.8
.ic q_88_19=0
.ic qb_88_19=1.8
.ic q_89_19=0
.ic qb_89_19=1.8
.ic q_90_19=0
.ic qb_90_19=1.8
.ic q_91_19=0
.ic qb_91_19=1.8
.ic q_92_19=0
.ic qb_92_19=1.8
.ic q_93_19=0
.ic qb_93_19=1.8
.ic q_94_19=0
.ic qb_94_19=1.8
.ic q_95_19=0
.ic qb_95_19=1.8
.ic q_96_19=0
.ic qb_96_19=1.8
.ic q_97_19=0
.ic qb_97_19=1.8
.ic q_98_19=0
.ic qb_98_19=1.8
.ic q_99_19=0
.ic qb_99_19=1.8
.ic q_0_20=0
.ic qb_0_20=1.8
.ic q_1_20=0
.ic qb_1_20=1.8
.ic q_2_20=0
.ic qb_2_20=1.8
.ic q_3_20=0
.ic qb_3_20=1.8
.ic q_4_20=0
.ic qb_4_20=1.8
.ic q_5_20=0
.ic qb_5_20=1.8
.ic q_6_20=0
.ic qb_6_20=1.8
.ic q_7_20=0
.ic qb_7_20=1.8
.ic q_8_20=0
.ic qb_8_20=1.8
.ic q_9_20=0
.ic qb_9_20=1.8
.ic q_10_20=0
.ic qb_10_20=1.8
.ic q_11_20=0
.ic qb_11_20=1.8
.ic q_12_20=0
.ic qb_12_20=1.8
.ic q_13_20=0
.ic qb_13_20=1.8
.ic q_14_20=0
.ic qb_14_20=1.8
.ic q_15_20=0
.ic qb_15_20=1.8
.ic q_16_20=0
.ic qb_16_20=1.8
.ic q_17_20=0
.ic qb_17_20=1.8
.ic q_18_20=0
.ic qb_18_20=1.8
.ic q_19_20=0
.ic qb_19_20=1.8
.ic q_20_20=0
.ic qb_20_20=1.8
.ic q_21_20=0
.ic qb_21_20=1.8
.ic q_22_20=0
.ic qb_22_20=1.8
.ic q_23_20=0
.ic qb_23_20=1.8
.ic q_24_20=0
.ic qb_24_20=1.8
.ic q_25_20=0
.ic qb_25_20=1.8
.ic q_26_20=0
.ic qb_26_20=1.8
.ic q_27_20=0
.ic qb_27_20=1.8
.ic q_28_20=0
.ic qb_28_20=1.8
.ic q_29_20=0
.ic qb_29_20=1.8
.ic q_30_20=0
.ic qb_30_20=1.8
.ic q_31_20=0
.ic qb_31_20=1.8
.ic q_32_20=0
.ic qb_32_20=1.8
.ic q_33_20=0
.ic qb_33_20=1.8
.ic q_34_20=0
.ic qb_34_20=1.8
.ic q_35_20=0
.ic qb_35_20=1.8
.ic q_36_20=0
.ic qb_36_20=1.8
.ic q_37_20=0
.ic qb_37_20=1.8
.ic q_38_20=0
.ic qb_38_20=1.8
.ic q_39_20=0
.ic qb_39_20=1.8
.ic q_40_20=0
.ic qb_40_20=1.8
.ic q_41_20=0
.ic qb_41_20=1.8
.ic q_42_20=0
.ic qb_42_20=1.8
.ic q_43_20=0
.ic qb_43_20=1.8
.ic q_44_20=0
.ic qb_44_20=1.8
.ic q_45_20=0
.ic qb_45_20=1.8
.ic q_46_20=0
.ic qb_46_20=1.8
.ic q_47_20=0
.ic qb_47_20=1.8
.ic q_48_20=0
.ic qb_48_20=1.8
.ic q_49_20=0
.ic qb_49_20=1.8
.ic q_50_20=0
.ic qb_50_20=1.8
.ic q_51_20=0
.ic qb_51_20=1.8
.ic q_52_20=0
.ic qb_52_20=1.8
.ic q_53_20=0
.ic qb_53_20=1.8
.ic q_54_20=0
.ic qb_54_20=1.8
.ic q_55_20=0
.ic qb_55_20=1.8
.ic q_56_20=0
.ic qb_56_20=1.8
.ic q_57_20=0
.ic qb_57_20=1.8
.ic q_58_20=0
.ic qb_58_20=1.8
.ic q_59_20=0
.ic qb_59_20=1.8
.ic q_60_20=0
.ic qb_60_20=1.8
.ic q_61_20=0
.ic qb_61_20=1.8
.ic q_62_20=0
.ic qb_62_20=1.8
.ic q_63_20=0
.ic qb_63_20=1.8
.ic q_64_20=0
.ic qb_64_20=1.8
.ic q_65_20=0
.ic qb_65_20=1.8
.ic q_66_20=0
.ic qb_66_20=1.8
.ic q_67_20=0
.ic qb_67_20=1.8
.ic q_68_20=0
.ic qb_68_20=1.8
.ic q_69_20=0
.ic qb_69_20=1.8
.ic q_70_20=0
.ic qb_70_20=1.8
.ic q_71_20=0
.ic qb_71_20=1.8
.ic q_72_20=0
.ic qb_72_20=1.8
.ic q_73_20=0
.ic qb_73_20=1.8
.ic q_74_20=0
.ic qb_74_20=1.8
.ic q_75_20=0
.ic qb_75_20=1.8
.ic q_76_20=0
.ic qb_76_20=1.8
.ic q_77_20=0
.ic qb_77_20=1.8
.ic q_78_20=0
.ic qb_78_20=1.8
.ic q_79_20=0
.ic qb_79_20=1.8
.ic q_80_20=0
.ic qb_80_20=1.8
.ic q_81_20=0
.ic qb_81_20=1.8
.ic q_82_20=0
.ic qb_82_20=1.8
.ic q_83_20=0
.ic qb_83_20=1.8
.ic q_84_20=0
.ic qb_84_20=1.8
.ic q_85_20=0
.ic qb_85_20=1.8
.ic q_86_20=0
.ic qb_86_20=1.8
.ic q_87_20=0
.ic qb_87_20=1.8
.ic q_88_20=0
.ic qb_88_20=1.8
.ic q_89_20=0
.ic qb_89_20=1.8
.ic q_90_20=0
.ic qb_90_20=1.8
.ic q_91_20=0
.ic qb_91_20=1.8
.ic q_92_20=0
.ic qb_92_20=1.8
.ic q_93_20=0
.ic qb_93_20=1.8
.ic q_94_20=0
.ic qb_94_20=1.8
.ic q_95_20=0
.ic qb_95_20=1.8
.ic q_96_20=0
.ic qb_96_20=1.8
.ic q_97_20=0
.ic qb_97_20=1.8
.ic q_98_20=0
.ic qb_98_20=1.8
.ic q_99_20=0
.ic qb_99_20=1.8
.ic q_0_21=0
.ic qb_0_21=1.8
.ic q_1_21=0
.ic qb_1_21=1.8
.ic q_2_21=0
.ic qb_2_21=1.8
.ic q_3_21=0
.ic qb_3_21=1.8
.ic q_4_21=0
.ic qb_4_21=1.8
.ic q_5_21=0
.ic qb_5_21=1.8
.ic q_6_21=0
.ic qb_6_21=1.8
.ic q_7_21=0
.ic qb_7_21=1.8
.ic q_8_21=0
.ic qb_8_21=1.8
.ic q_9_21=0
.ic qb_9_21=1.8
.ic q_10_21=0
.ic qb_10_21=1.8
.ic q_11_21=0
.ic qb_11_21=1.8
.ic q_12_21=0
.ic qb_12_21=1.8
.ic q_13_21=0
.ic qb_13_21=1.8
.ic q_14_21=0
.ic qb_14_21=1.8
.ic q_15_21=0
.ic qb_15_21=1.8
.ic q_16_21=0
.ic qb_16_21=1.8
.ic q_17_21=0
.ic qb_17_21=1.8
.ic q_18_21=0
.ic qb_18_21=1.8
.ic q_19_21=0
.ic qb_19_21=1.8
.ic q_20_21=0
.ic qb_20_21=1.8
.ic q_21_21=0
.ic qb_21_21=1.8
.ic q_22_21=0
.ic qb_22_21=1.8
.ic q_23_21=0
.ic qb_23_21=1.8
.ic q_24_21=0
.ic qb_24_21=1.8
.ic q_25_21=0
.ic qb_25_21=1.8
.ic q_26_21=0
.ic qb_26_21=1.8
.ic q_27_21=0
.ic qb_27_21=1.8
.ic q_28_21=0
.ic qb_28_21=1.8
.ic q_29_21=0
.ic qb_29_21=1.8
.ic q_30_21=0
.ic qb_30_21=1.8
.ic q_31_21=0
.ic qb_31_21=1.8
.ic q_32_21=0
.ic qb_32_21=1.8
.ic q_33_21=0
.ic qb_33_21=1.8
.ic q_34_21=0
.ic qb_34_21=1.8
.ic q_35_21=0
.ic qb_35_21=1.8
.ic q_36_21=0
.ic qb_36_21=1.8
.ic q_37_21=0
.ic qb_37_21=1.8
.ic q_38_21=0
.ic qb_38_21=1.8
.ic q_39_21=0
.ic qb_39_21=1.8
.ic q_40_21=0
.ic qb_40_21=1.8
.ic q_41_21=0
.ic qb_41_21=1.8
.ic q_42_21=0
.ic qb_42_21=1.8
.ic q_43_21=0
.ic qb_43_21=1.8
.ic q_44_21=0
.ic qb_44_21=1.8
.ic q_45_21=0
.ic qb_45_21=1.8
.ic q_46_21=0
.ic qb_46_21=1.8
.ic q_47_21=0
.ic qb_47_21=1.8
.ic q_48_21=0
.ic qb_48_21=1.8
.ic q_49_21=0
.ic qb_49_21=1.8
.ic q_50_21=0
.ic qb_50_21=1.8
.ic q_51_21=0
.ic qb_51_21=1.8
.ic q_52_21=0
.ic qb_52_21=1.8
.ic q_53_21=0
.ic qb_53_21=1.8
.ic q_54_21=0
.ic qb_54_21=1.8
.ic q_55_21=0
.ic qb_55_21=1.8
.ic q_56_21=0
.ic qb_56_21=1.8
.ic q_57_21=0
.ic qb_57_21=1.8
.ic q_58_21=0
.ic qb_58_21=1.8
.ic q_59_21=0
.ic qb_59_21=1.8
.ic q_60_21=0
.ic qb_60_21=1.8
.ic q_61_21=0
.ic qb_61_21=1.8
.ic q_62_21=0
.ic qb_62_21=1.8
.ic q_63_21=0
.ic qb_63_21=1.8
.ic q_64_21=0
.ic qb_64_21=1.8
.ic q_65_21=0
.ic qb_65_21=1.8
.ic q_66_21=0
.ic qb_66_21=1.8
.ic q_67_21=0
.ic qb_67_21=1.8
.ic q_68_21=0
.ic qb_68_21=1.8
.ic q_69_21=0
.ic qb_69_21=1.8
.ic q_70_21=0
.ic qb_70_21=1.8
.ic q_71_21=0
.ic qb_71_21=1.8
.ic q_72_21=0
.ic qb_72_21=1.8
.ic q_73_21=0
.ic qb_73_21=1.8
.ic q_74_21=0
.ic qb_74_21=1.8
.ic q_75_21=0
.ic qb_75_21=1.8
.ic q_76_21=0
.ic qb_76_21=1.8
.ic q_77_21=0
.ic qb_77_21=1.8
.ic q_78_21=0
.ic qb_78_21=1.8
.ic q_79_21=0
.ic qb_79_21=1.8
.ic q_80_21=0
.ic qb_80_21=1.8
.ic q_81_21=0
.ic qb_81_21=1.8
.ic q_82_21=0
.ic qb_82_21=1.8
.ic q_83_21=0
.ic qb_83_21=1.8
.ic q_84_21=0
.ic qb_84_21=1.8
.ic q_85_21=0
.ic qb_85_21=1.8
.ic q_86_21=0
.ic qb_86_21=1.8
.ic q_87_21=0
.ic qb_87_21=1.8
.ic q_88_21=0
.ic qb_88_21=1.8
.ic q_89_21=0
.ic qb_89_21=1.8
.ic q_90_21=0
.ic qb_90_21=1.8
.ic q_91_21=0
.ic qb_91_21=1.8
.ic q_92_21=0
.ic qb_92_21=1.8
.ic q_93_21=0
.ic qb_93_21=1.8
.ic q_94_21=0
.ic qb_94_21=1.8
.ic q_95_21=0
.ic qb_95_21=1.8
.ic q_96_21=0
.ic qb_96_21=1.8
.ic q_97_21=0
.ic qb_97_21=1.8
.ic q_98_21=0
.ic qb_98_21=1.8
.ic q_99_21=0
.ic qb_99_21=1.8
.ic q_0_22=0
.ic qb_0_22=1.8
.ic q_1_22=0
.ic qb_1_22=1.8
.ic q_2_22=0
.ic qb_2_22=1.8
.ic q_3_22=0
.ic qb_3_22=1.8
.ic q_4_22=0
.ic qb_4_22=1.8
.ic q_5_22=0
.ic qb_5_22=1.8
.ic q_6_22=0
.ic qb_6_22=1.8
.ic q_7_22=0
.ic qb_7_22=1.8
.ic q_8_22=0
.ic qb_8_22=1.8
.ic q_9_22=0
.ic qb_9_22=1.8
.ic q_10_22=0
.ic qb_10_22=1.8
.ic q_11_22=0
.ic qb_11_22=1.8
.ic q_12_22=0
.ic qb_12_22=1.8
.ic q_13_22=0
.ic qb_13_22=1.8
.ic q_14_22=0
.ic qb_14_22=1.8
.ic q_15_22=0
.ic qb_15_22=1.8
.ic q_16_22=0
.ic qb_16_22=1.8
.ic q_17_22=0
.ic qb_17_22=1.8
.ic q_18_22=0
.ic qb_18_22=1.8
.ic q_19_22=0
.ic qb_19_22=1.8
.ic q_20_22=0
.ic qb_20_22=1.8
.ic q_21_22=0
.ic qb_21_22=1.8
.ic q_22_22=0
.ic qb_22_22=1.8
.ic q_23_22=0
.ic qb_23_22=1.8
.ic q_24_22=0
.ic qb_24_22=1.8
.ic q_25_22=0
.ic qb_25_22=1.8
.ic q_26_22=0
.ic qb_26_22=1.8
.ic q_27_22=0
.ic qb_27_22=1.8
.ic q_28_22=0
.ic qb_28_22=1.8
.ic q_29_22=0
.ic qb_29_22=1.8
.ic q_30_22=0
.ic qb_30_22=1.8
.ic q_31_22=0
.ic qb_31_22=1.8
.ic q_32_22=0
.ic qb_32_22=1.8
.ic q_33_22=0
.ic qb_33_22=1.8
.ic q_34_22=0
.ic qb_34_22=1.8
.ic q_35_22=0
.ic qb_35_22=1.8
.ic q_36_22=0
.ic qb_36_22=1.8
.ic q_37_22=0
.ic qb_37_22=1.8
.ic q_38_22=0
.ic qb_38_22=1.8
.ic q_39_22=0
.ic qb_39_22=1.8
.ic q_40_22=0
.ic qb_40_22=1.8
.ic q_41_22=0
.ic qb_41_22=1.8
.ic q_42_22=0
.ic qb_42_22=1.8
.ic q_43_22=0
.ic qb_43_22=1.8
.ic q_44_22=0
.ic qb_44_22=1.8
.ic q_45_22=0
.ic qb_45_22=1.8
.ic q_46_22=0
.ic qb_46_22=1.8
.ic q_47_22=0
.ic qb_47_22=1.8
.ic q_48_22=0
.ic qb_48_22=1.8
.ic q_49_22=0
.ic qb_49_22=1.8
.ic q_50_22=0
.ic qb_50_22=1.8
.ic q_51_22=0
.ic qb_51_22=1.8
.ic q_52_22=0
.ic qb_52_22=1.8
.ic q_53_22=0
.ic qb_53_22=1.8
.ic q_54_22=0
.ic qb_54_22=1.8
.ic q_55_22=0
.ic qb_55_22=1.8
.ic q_56_22=0
.ic qb_56_22=1.8
.ic q_57_22=0
.ic qb_57_22=1.8
.ic q_58_22=0
.ic qb_58_22=1.8
.ic q_59_22=0
.ic qb_59_22=1.8
.ic q_60_22=0
.ic qb_60_22=1.8
.ic q_61_22=0
.ic qb_61_22=1.8
.ic q_62_22=0
.ic qb_62_22=1.8
.ic q_63_22=0
.ic qb_63_22=1.8
.ic q_64_22=0
.ic qb_64_22=1.8
.ic q_65_22=0
.ic qb_65_22=1.8
.ic q_66_22=0
.ic qb_66_22=1.8
.ic q_67_22=0
.ic qb_67_22=1.8
.ic q_68_22=0
.ic qb_68_22=1.8
.ic q_69_22=0
.ic qb_69_22=1.8
.ic q_70_22=0
.ic qb_70_22=1.8
.ic q_71_22=0
.ic qb_71_22=1.8
.ic q_72_22=0
.ic qb_72_22=1.8
.ic q_73_22=0
.ic qb_73_22=1.8
.ic q_74_22=0
.ic qb_74_22=1.8
.ic q_75_22=0
.ic qb_75_22=1.8
.ic q_76_22=0
.ic qb_76_22=1.8
.ic q_77_22=0
.ic qb_77_22=1.8
.ic q_78_22=0
.ic qb_78_22=1.8
.ic q_79_22=0
.ic qb_79_22=1.8
.ic q_80_22=0
.ic qb_80_22=1.8
.ic q_81_22=0
.ic qb_81_22=1.8
.ic q_82_22=0
.ic qb_82_22=1.8
.ic q_83_22=0
.ic qb_83_22=1.8
.ic q_84_22=0
.ic qb_84_22=1.8
.ic q_85_22=0
.ic qb_85_22=1.8
.ic q_86_22=0
.ic qb_86_22=1.8
.ic q_87_22=0
.ic qb_87_22=1.8
.ic q_88_22=0
.ic qb_88_22=1.8
.ic q_89_22=0
.ic qb_89_22=1.8
.ic q_90_22=0
.ic qb_90_22=1.8
.ic q_91_22=0
.ic qb_91_22=1.8
.ic q_92_22=0
.ic qb_92_22=1.8
.ic q_93_22=0
.ic qb_93_22=1.8
.ic q_94_22=0
.ic qb_94_22=1.8
.ic q_95_22=0
.ic qb_95_22=1.8
.ic q_96_22=0
.ic qb_96_22=1.8
.ic q_97_22=0
.ic qb_97_22=1.8
.ic q_98_22=0
.ic qb_98_22=1.8
.ic q_99_22=0
.ic qb_99_22=1.8
.ic q_0_23=0
.ic qb_0_23=1.8
.ic q_1_23=0
.ic qb_1_23=1.8
.ic q_2_23=0
.ic qb_2_23=1.8
.ic q_3_23=0
.ic qb_3_23=1.8
.ic q_4_23=0
.ic qb_4_23=1.8
.ic q_5_23=0
.ic qb_5_23=1.8
.ic q_6_23=0
.ic qb_6_23=1.8
.ic q_7_23=0
.ic qb_7_23=1.8
.ic q_8_23=0
.ic qb_8_23=1.8
.ic q_9_23=0
.ic qb_9_23=1.8
.ic q_10_23=0
.ic qb_10_23=1.8
.ic q_11_23=0
.ic qb_11_23=1.8
.ic q_12_23=0
.ic qb_12_23=1.8
.ic q_13_23=0
.ic qb_13_23=1.8
.ic q_14_23=0
.ic qb_14_23=1.8
.ic q_15_23=0
.ic qb_15_23=1.8
.ic q_16_23=0
.ic qb_16_23=1.8
.ic q_17_23=0
.ic qb_17_23=1.8
.ic q_18_23=0
.ic qb_18_23=1.8
.ic q_19_23=0
.ic qb_19_23=1.8
.ic q_20_23=0
.ic qb_20_23=1.8
.ic q_21_23=0
.ic qb_21_23=1.8
.ic q_22_23=0
.ic qb_22_23=1.8
.ic q_23_23=0
.ic qb_23_23=1.8
.ic q_24_23=0
.ic qb_24_23=1.8
.ic q_25_23=0
.ic qb_25_23=1.8
.ic q_26_23=0
.ic qb_26_23=1.8
.ic q_27_23=0
.ic qb_27_23=1.8
.ic q_28_23=0
.ic qb_28_23=1.8
.ic q_29_23=0
.ic qb_29_23=1.8
.ic q_30_23=0
.ic qb_30_23=1.8
.ic q_31_23=0
.ic qb_31_23=1.8
.ic q_32_23=0
.ic qb_32_23=1.8
.ic q_33_23=0
.ic qb_33_23=1.8
.ic q_34_23=0
.ic qb_34_23=1.8
.ic q_35_23=0
.ic qb_35_23=1.8
.ic q_36_23=0
.ic qb_36_23=1.8
.ic q_37_23=0
.ic qb_37_23=1.8
.ic q_38_23=0
.ic qb_38_23=1.8
.ic q_39_23=0
.ic qb_39_23=1.8
.ic q_40_23=0
.ic qb_40_23=1.8
.ic q_41_23=0
.ic qb_41_23=1.8
.ic q_42_23=0
.ic qb_42_23=1.8
.ic q_43_23=0
.ic qb_43_23=1.8
.ic q_44_23=0
.ic qb_44_23=1.8
.ic q_45_23=0
.ic qb_45_23=1.8
.ic q_46_23=0
.ic qb_46_23=1.8
.ic q_47_23=0
.ic qb_47_23=1.8
.ic q_48_23=0
.ic qb_48_23=1.8
.ic q_49_23=0
.ic qb_49_23=1.8
.ic q_50_23=0
.ic qb_50_23=1.8
.ic q_51_23=0
.ic qb_51_23=1.8
.ic q_52_23=0
.ic qb_52_23=1.8
.ic q_53_23=0
.ic qb_53_23=1.8
.ic q_54_23=0
.ic qb_54_23=1.8
.ic q_55_23=0
.ic qb_55_23=1.8
.ic q_56_23=0
.ic qb_56_23=1.8
.ic q_57_23=0
.ic qb_57_23=1.8
.ic q_58_23=0
.ic qb_58_23=1.8
.ic q_59_23=0
.ic qb_59_23=1.8
.ic q_60_23=0
.ic qb_60_23=1.8
.ic q_61_23=0
.ic qb_61_23=1.8
.ic q_62_23=0
.ic qb_62_23=1.8
.ic q_63_23=0
.ic qb_63_23=1.8
.ic q_64_23=0
.ic qb_64_23=1.8
.ic q_65_23=0
.ic qb_65_23=1.8
.ic q_66_23=0
.ic qb_66_23=1.8
.ic q_67_23=0
.ic qb_67_23=1.8
.ic q_68_23=0
.ic qb_68_23=1.8
.ic q_69_23=0
.ic qb_69_23=1.8
.ic q_70_23=0
.ic qb_70_23=1.8
.ic q_71_23=0
.ic qb_71_23=1.8
.ic q_72_23=0
.ic qb_72_23=1.8
.ic q_73_23=0
.ic qb_73_23=1.8
.ic q_74_23=0
.ic qb_74_23=1.8
.ic q_75_23=0
.ic qb_75_23=1.8
.ic q_76_23=0
.ic qb_76_23=1.8
.ic q_77_23=0
.ic qb_77_23=1.8
.ic q_78_23=0
.ic qb_78_23=1.8
.ic q_79_23=0
.ic qb_79_23=1.8
.ic q_80_23=0
.ic qb_80_23=1.8
.ic q_81_23=0
.ic qb_81_23=1.8
.ic q_82_23=0
.ic qb_82_23=1.8
.ic q_83_23=0
.ic qb_83_23=1.8
.ic q_84_23=0
.ic qb_84_23=1.8
.ic q_85_23=0
.ic qb_85_23=1.8
.ic q_86_23=0
.ic qb_86_23=1.8
.ic q_87_23=0
.ic qb_87_23=1.8
.ic q_88_23=0
.ic qb_88_23=1.8
.ic q_89_23=0
.ic qb_89_23=1.8
.ic q_90_23=0
.ic qb_90_23=1.8
.ic q_91_23=0
.ic qb_91_23=1.8
.ic q_92_23=0
.ic qb_92_23=1.8
.ic q_93_23=0
.ic qb_93_23=1.8
.ic q_94_23=0
.ic qb_94_23=1.8
.ic q_95_23=0
.ic qb_95_23=1.8
.ic q_96_23=0
.ic qb_96_23=1.8
.ic q_97_23=0
.ic qb_97_23=1.8
.ic q_98_23=0
.ic qb_98_23=1.8
.ic q_99_23=0
.ic qb_99_23=1.8
.ic q_0_24=0
.ic qb_0_24=1.8
.ic q_1_24=0
.ic qb_1_24=1.8
.ic q_2_24=0
.ic qb_2_24=1.8
.ic q_3_24=0
.ic qb_3_24=1.8
.ic q_4_24=0
.ic qb_4_24=1.8
.ic q_5_24=0
.ic qb_5_24=1.8
.ic q_6_24=0
.ic qb_6_24=1.8
.ic q_7_24=0
.ic qb_7_24=1.8
.ic q_8_24=0
.ic qb_8_24=1.8
.ic q_9_24=0
.ic qb_9_24=1.8
.ic q_10_24=0
.ic qb_10_24=1.8
.ic q_11_24=0
.ic qb_11_24=1.8
.ic q_12_24=0
.ic qb_12_24=1.8
.ic q_13_24=0
.ic qb_13_24=1.8
.ic q_14_24=0
.ic qb_14_24=1.8
.ic q_15_24=0
.ic qb_15_24=1.8
.ic q_16_24=0
.ic qb_16_24=1.8
.ic q_17_24=0
.ic qb_17_24=1.8
.ic q_18_24=0
.ic qb_18_24=1.8
.ic q_19_24=0
.ic qb_19_24=1.8
.ic q_20_24=0
.ic qb_20_24=1.8
.ic q_21_24=0
.ic qb_21_24=1.8
.ic q_22_24=0
.ic qb_22_24=1.8
.ic q_23_24=0
.ic qb_23_24=1.8
.ic q_24_24=0
.ic qb_24_24=1.8
.ic q_25_24=0
.ic qb_25_24=1.8
.ic q_26_24=0
.ic qb_26_24=1.8
.ic q_27_24=0
.ic qb_27_24=1.8
.ic q_28_24=0
.ic qb_28_24=1.8
.ic q_29_24=0
.ic qb_29_24=1.8
.ic q_30_24=0
.ic qb_30_24=1.8
.ic q_31_24=0
.ic qb_31_24=1.8
.ic q_32_24=0
.ic qb_32_24=1.8
.ic q_33_24=0
.ic qb_33_24=1.8
.ic q_34_24=0
.ic qb_34_24=1.8
.ic q_35_24=0
.ic qb_35_24=1.8
.ic q_36_24=0
.ic qb_36_24=1.8
.ic q_37_24=0
.ic qb_37_24=1.8
.ic q_38_24=0
.ic qb_38_24=1.8
.ic q_39_24=0
.ic qb_39_24=1.8
.ic q_40_24=0
.ic qb_40_24=1.8
.ic q_41_24=0
.ic qb_41_24=1.8
.ic q_42_24=0
.ic qb_42_24=1.8
.ic q_43_24=0
.ic qb_43_24=1.8
.ic q_44_24=0
.ic qb_44_24=1.8
.ic q_45_24=0
.ic qb_45_24=1.8
.ic q_46_24=0
.ic qb_46_24=1.8
.ic q_47_24=0
.ic qb_47_24=1.8
.ic q_48_24=0
.ic qb_48_24=1.8
.ic q_49_24=0
.ic qb_49_24=1.8
.ic q_50_24=0
.ic qb_50_24=1.8
.ic q_51_24=0
.ic qb_51_24=1.8
.ic q_52_24=0
.ic qb_52_24=1.8
.ic q_53_24=0
.ic qb_53_24=1.8
.ic q_54_24=0
.ic qb_54_24=1.8
.ic q_55_24=0
.ic qb_55_24=1.8
.ic q_56_24=0
.ic qb_56_24=1.8
.ic q_57_24=0
.ic qb_57_24=1.8
.ic q_58_24=0
.ic qb_58_24=1.8
.ic q_59_24=0
.ic qb_59_24=1.8
.ic q_60_24=0
.ic qb_60_24=1.8
.ic q_61_24=0
.ic qb_61_24=1.8
.ic q_62_24=0
.ic qb_62_24=1.8
.ic q_63_24=0
.ic qb_63_24=1.8
.ic q_64_24=0
.ic qb_64_24=1.8
.ic q_65_24=0
.ic qb_65_24=1.8
.ic q_66_24=0
.ic qb_66_24=1.8
.ic q_67_24=0
.ic qb_67_24=1.8
.ic q_68_24=0
.ic qb_68_24=1.8
.ic q_69_24=0
.ic qb_69_24=1.8
.ic q_70_24=0
.ic qb_70_24=1.8
.ic q_71_24=0
.ic qb_71_24=1.8
.ic q_72_24=0
.ic qb_72_24=1.8
.ic q_73_24=0
.ic qb_73_24=1.8
.ic q_74_24=0
.ic qb_74_24=1.8
.ic q_75_24=0
.ic qb_75_24=1.8
.ic q_76_24=0
.ic qb_76_24=1.8
.ic q_77_24=0
.ic qb_77_24=1.8
.ic q_78_24=0
.ic qb_78_24=1.8
.ic q_79_24=0
.ic qb_79_24=1.8
.ic q_80_24=0
.ic qb_80_24=1.8
.ic q_81_24=0
.ic qb_81_24=1.8
.ic q_82_24=0
.ic qb_82_24=1.8
.ic q_83_24=0
.ic qb_83_24=1.8
.ic q_84_24=0
.ic qb_84_24=1.8
.ic q_85_24=0
.ic qb_85_24=1.8
.ic q_86_24=0
.ic qb_86_24=1.8
.ic q_87_24=0
.ic qb_87_24=1.8
.ic q_88_24=0
.ic qb_88_24=1.8
.ic q_89_24=0
.ic qb_89_24=1.8
.ic q_90_24=0
.ic qb_90_24=1.8
.ic q_91_24=0
.ic qb_91_24=1.8
.ic q_92_24=0
.ic qb_92_24=1.8
.ic q_93_24=0
.ic qb_93_24=1.8
.ic q_94_24=0
.ic qb_94_24=1.8
.ic q_95_24=0
.ic qb_95_24=1.8
.ic q_96_24=0
.ic qb_96_24=1.8
.ic q_97_24=0
.ic qb_97_24=1.8
.ic q_98_24=0
.ic qb_98_24=1.8
.ic q_99_24=0
.ic qb_99_24=1.8
.ic q_0_25=0
.ic qb_0_25=1.8
.ic q_1_25=0
.ic qb_1_25=1.8
.ic q_2_25=0
.ic qb_2_25=1.8
.ic q_3_25=0
.ic qb_3_25=1.8
.ic q_4_25=0
.ic qb_4_25=1.8
.ic q_5_25=0
.ic qb_5_25=1.8
.ic q_6_25=0
.ic qb_6_25=1.8
.ic q_7_25=0
.ic qb_7_25=1.8
.ic q_8_25=0
.ic qb_8_25=1.8
.ic q_9_25=0
.ic qb_9_25=1.8
.ic q_10_25=0
.ic qb_10_25=1.8
.ic q_11_25=0
.ic qb_11_25=1.8
.ic q_12_25=0
.ic qb_12_25=1.8
.ic q_13_25=0
.ic qb_13_25=1.8
.ic q_14_25=0
.ic qb_14_25=1.8
.ic q_15_25=0
.ic qb_15_25=1.8
.ic q_16_25=0
.ic qb_16_25=1.8
.ic q_17_25=0
.ic qb_17_25=1.8
.ic q_18_25=0
.ic qb_18_25=1.8
.ic q_19_25=0
.ic qb_19_25=1.8
.ic q_20_25=0
.ic qb_20_25=1.8
.ic q_21_25=0
.ic qb_21_25=1.8
.ic q_22_25=0
.ic qb_22_25=1.8
.ic q_23_25=0
.ic qb_23_25=1.8
.ic q_24_25=0
.ic qb_24_25=1.8
.ic q_25_25=0
.ic qb_25_25=1.8
.ic q_26_25=0
.ic qb_26_25=1.8
.ic q_27_25=0
.ic qb_27_25=1.8
.ic q_28_25=0
.ic qb_28_25=1.8
.ic q_29_25=0
.ic qb_29_25=1.8
.ic q_30_25=0
.ic qb_30_25=1.8
.ic q_31_25=0
.ic qb_31_25=1.8
.ic q_32_25=0
.ic qb_32_25=1.8
.ic q_33_25=0
.ic qb_33_25=1.8
.ic q_34_25=0
.ic qb_34_25=1.8
.ic q_35_25=0
.ic qb_35_25=1.8
.ic q_36_25=0
.ic qb_36_25=1.8
.ic q_37_25=0
.ic qb_37_25=1.8
.ic q_38_25=0
.ic qb_38_25=1.8
.ic q_39_25=0
.ic qb_39_25=1.8
.ic q_40_25=0
.ic qb_40_25=1.8
.ic q_41_25=0
.ic qb_41_25=1.8
.ic q_42_25=0
.ic qb_42_25=1.8
.ic q_43_25=0
.ic qb_43_25=1.8
.ic q_44_25=0
.ic qb_44_25=1.8
.ic q_45_25=0
.ic qb_45_25=1.8
.ic q_46_25=0
.ic qb_46_25=1.8
.ic q_47_25=0
.ic qb_47_25=1.8
.ic q_48_25=0
.ic qb_48_25=1.8
.ic q_49_25=0
.ic qb_49_25=1.8
.ic q_50_25=0
.ic qb_50_25=1.8
.ic q_51_25=0
.ic qb_51_25=1.8
.ic q_52_25=0
.ic qb_52_25=1.8
.ic q_53_25=0
.ic qb_53_25=1.8
.ic q_54_25=0
.ic qb_54_25=1.8
.ic q_55_25=0
.ic qb_55_25=1.8
.ic q_56_25=0
.ic qb_56_25=1.8
.ic q_57_25=0
.ic qb_57_25=1.8
.ic q_58_25=0
.ic qb_58_25=1.8
.ic q_59_25=0
.ic qb_59_25=1.8
.ic q_60_25=0
.ic qb_60_25=1.8
.ic q_61_25=0
.ic qb_61_25=1.8
.ic q_62_25=0
.ic qb_62_25=1.8
.ic q_63_25=0
.ic qb_63_25=1.8
.ic q_64_25=0
.ic qb_64_25=1.8
.ic q_65_25=0
.ic qb_65_25=1.8
.ic q_66_25=0
.ic qb_66_25=1.8
.ic q_67_25=0
.ic qb_67_25=1.8
.ic q_68_25=0
.ic qb_68_25=1.8
.ic q_69_25=0
.ic qb_69_25=1.8
.ic q_70_25=0
.ic qb_70_25=1.8
.ic q_71_25=0
.ic qb_71_25=1.8
.ic q_72_25=0
.ic qb_72_25=1.8
.ic q_73_25=0
.ic qb_73_25=1.8
.ic q_74_25=0
.ic qb_74_25=1.8
.ic q_75_25=0
.ic qb_75_25=1.8
.ic q_76_25=0
.ic qb_76_25=1.8
.ic q_77_25=0
.ic qb_77_25=1.8
.ic q_78_25=0
.ic qb_78_25=1.8
.ic q_79_25=0
.ic qb_79_25=1.8
.ic q_80_25=0
.ic qb_80_25=1.8
.ic q_81_25=0
.ic qb_81_25=1.8
.ic q_82_25=0
.ic qb_82_25=1.8
.ic q_83_25=0
.ic qb_83_25=1.8
.ic q_84_25=0
.ic qb_84_25=1.8
.ic q_85_25=0
.ic qb_85_25=1.8
.ic q_86_25=0
.ic qb_86_25=1.8
.ic q_87_25=0
.ic qb_87_25=1.8
.ic q_88_25=0
.ic qb_88_25=1.8
.ic q_89_25=0
.ic qb_89_25=1.8
.ic q_90_25=0
.ic qb_90_25=1.8
.ic q_91_25=0
.ic qb_91_25=1.8
.ic q_92_25=0
.ic qb_92_25=1.8
.ic q_93_25=0
.ic qb_93_25=1.8
.ic q_94_25=0
.ic qb_94_25=1.8
.ic q_95_25=0
.ic qb_95_25=1.8
.ic q_96_25=0
.ic qb_96_25=1.8
.ic q_97_25=0
.ic qb_97_25=1.8
.ic q_98_25=0
.ic qb_98_25=1.8
.ic q_99_25=0
.ic qb_99_25=1.8
.ic q_0_26=0
.ic qb_0_26=1.8
.ic q_1_26=0
.ic qb_1_26=1.8
.ic q_2_26=0
.ic qb_2_26=1.8
.ic q_3_26=0
.ic qb_3_26=1.8
.ic q_4_26=0
.ic qb_4_26=1.8
.ic q_5_26=0
.ic qb_5_26=1.8
.ic q_6_26=0
.ic qb_6_26=1.8
.ic q_7_26=0
.ic qb_7_26=1.8
.ic q_8_26=0
.ic qb_8_26=1.8
.ic q_9_26=0
.ic qb_9_26=1.8
.ic q_10_26=0
.ic qb_10_26=1.8
.ic q_11_26=0
.ic qb_11_26=1.8
.ic q_12_26=0
.ic qb_12_26=1.8
.ic q_13_26=0
.ic qb_13_26=1.8
.ic q_14_26=0
.ic qb_14_26=1.8
.ic q_15_26=0
.ic qb_15_26=1.8
.ic q_16_26=0
.ic qb_16_26=1.8
.ic q_17_26=0
.ic qb_17_26=1.8
.ic q_18_26=0
.ic qb_18_26=1.8
.ic q_19_26=0
.ic qb_19_26=1.8
.ic q_20_26=0
.ic qb_20_26=1.8
.ic q_21_26=0
.ic qb_21_26=1.8
.ic q_22_26=0
.ic qb_22_26=1.8
.ic q_23_26=0
.ic qb_23_26=1.8
.ic q_24_26=0
.ic qb_24_26=1.8
.ic q_25_26=0
.ic qb_25_26=1.8
.ic q_26_26=0
.ic qb_26_26=1.8
.ic q_27_26=0
.ic qb_27_26=1.8
.ic q_28_26=0
.ic qb_28_26=1.8
.ic q_29_26=0
.ic qb_29_26=1.8
.ic q_30_26=0
.ic qb_30_26=1.8
.ic q_31_26=0
.ic qb_31_26=1.8
.ic q_32_26=0
.ic qb_32_26=1.8
.ic q_33_26=0
.ic qb_33_26=1.8
.ic q_34_26=0
.ic qb_34_26=1.8
.ic q_35_26=0
.ic qb_35_26=1.8
.ic q_36_26=0
.ic qb_36_26=1.8
.ic q_37_26=0
.ic qb_37_26=1.8
.ic q_38_26=0
.ic qb_38_26=1.8
.ic q_39_26=0
.ic qb_39_26=1.8
.ic q_40_26=0
.ic qb_40_26=1.8
.ic q_41_26=0
.ic qb_41_26=1.8
.ic q_42_26=0
.ic qb_42_26=1.8
.ic q_43_26=0
.ic qb_43_26=1.8
.ic q_44_26=0
.ic qb_44_26=1.8
.ic q_45_26=0
.ic qb_45_26=1.8
.ic q_46_26=0
.ic qb_46_26=1.8
.ic q_47_26=0
.ic qb_47_26=1.8
.ic q_48_26=0
.ic qb_48_26=1.8
.ic q_49_26=0
.ic qb_49_26=1.8
.ic q_50_26=0
.ic qb_50_26=1.8
.ic q_51_26=0
.ic qb_51_26=1.8
.ic q_52_26=0
.ic qb_52_26=1.8
.ic q_53_26=0
.ic qb_53_26=1.8
.ic q_54_26=0
.ic qb_54_26=1.8
.ic q_55_26=0
.ic qb_55_26=1.8
.ic q_56_26=0
.ic qb_56_26=1.8
.ic q_57_26=0
.ic qb_57_26=1.8
.ic q_58_26=0
.ic qb_58_26=1.8
.ic q_59_26=0
.ic qb_59_26=1.8
.ic q_60_26=0
.ic qb_60_26=1.8
.ic q_61_26=0
.ic qb_61_26=1.8
.ic q_62_26=0
.ic qb_62_26=1.8
.ic q_63_26=0
.ic qb_63_26=1.8
.ic q_64_26=0
.ic qb_64_26=1.8
.ic q_65_26=0
.ic qb_65_26=1.8
.ic q_66_26=0
.ic qb_66_26=1.8
.ic q_67_26=0
.ic qb_67_26=1.8
.ic q_68_26=0
.ic qb_68_26=1.8
.ic q_69_26=0
.ic qb_69_26=1.8
.ic q_70_26=0
.ic qb_70_26=1.8
.ic q_71_26=0
.ic qb_71_26=1.8
.ic q_72_26=0
.ic qb_72_26=1.8
.ic q_73_26=0
.ic qb_73_26=1.8
.ic q_74_26=0
.ic qb_74_26=1.8
.ic q_75_26=0
.ic qb_75_26=1.8
.ic q_76_26=0
.ic qb_76_26=1.8
.ic q_77_26=0
.ic qb_77_26=1.8
.ic q_78_26=0
.ic qb_78_26=1.8
.ic q_79_26=0
.ic qb_79_26=1.8
.ic q_80_26=0
.ic qb_80_26=1.8
.ic q_81_26=0
.ic qb_81_26=1.8
.ic q_82_26=0
.ic qb_82_26=1.8
.ic q_83_26=0
.ic qb_83_26=1.8
.ic q_84_26=0
.ic qb_84_26=1.8
.ic q_85_26=0
.ic qb_85_26=1.8
.ic q_86_26=0
.ic qb_86_26=1.8
.ic q_87_26=0
.ic qb_87_26=1.8
.ic q_88_26=0
.ic qb_88_26=1.8
.ic q_89_26=0
.ic qb_89_26=1.8
.ic q_90_26=0
.ic qb_90_26=1.8
.ic q_91_26=0
.ic qb_91_26=1.8
.ic q_92_26=0
.ic qb_92_26=1.8
.ic q_93_26=0
.ic qb_93_26=1.8
.ic q_94_26=0
.ic qb_94_26=1.8
.ic q_95_26=0
.ic qb_95_26=1.8
.ic q_96_26=0
.ic qb_96_26=1.8
.ic q_97_26=0
.ic qb_97_26=1.8
.ic q_98_26=0
.ic qb_98_26=1.8
.ic q_99_26=0
.ic qb_99_26=1.8
.ic q_0_27=0
.ic qb_0_27=1.8
.ic q_1_27=0
.ic qb_1_27=1.8
.ic q_2_27=0
.ic qb_2_27=1.8
.ic q_3_27=0
.ic qb_3_27=1.8
.ic q_4_27=0
.ic qb_4_27=1.8
.ic q_5_27=0
.ic qb_5_27=1.8
.ic q_6_27=0
.ic qb_6_27=1.8
.ic q_7_27=0
.ic qb_7_27=1.8
.ic q_8_27=0
.ic qb_8_27=1.8
.ic q_9_27=0
.ic qb_9_27=1.8
.ic q_10_27=0
.ic qb_10_27=1.8
.ic q_11_27=0
.ic qb_11_27=1.8
.ic q_12_27=0
.ic qb_12_27=1.8
.ic q_13_27=0
.ic qb_13_27=1.8
.ic q_14_27=0
.ic qb_14_27=1.8
.ic q_15_27=0
.ic qb_15_27=1.8
.ic q_16_27=0
.ic qb_16_27=1.8
.ic q_17_27=0
.ic qb_17_27=1.8
.ic q_18_27=0
.ic qb_18_27=1.8
.ic q_19_27=0
.ic qb_19_27=1.8
.ic q_20_27=0
.ic qb_20_27=1.8
.ic q_21_27=0
.ic qb_21_27=1.8
.ic q_22_27=0
.ic qb_22_27=1.8
.ic q_23_27=0
.ic qb_23_27=1.8
.ic q_24_27=0
.ic qb_24_27=1.8
.ic q_25_27=0
.ic qb_25_27=1.8
.ic q_26_27=0
.ic qb_26_27=1.8
.ic q_27_27=0
.ic qb_27_27=1.8
.ic q_28_27=0
.ic qb_28_27=1.8
.ic q_29_27=0
.ic qb_29_27=1.8
.ic q_30_27=0
.ic qb_30_27=1.8
.ic q_31_27=0
.ic qb_31_27=1.8
.ic q_32_27=0
.ic qb_32_27=1.8
.ic q_33_27=0
.ic qb_33_27=1.8
.ic q_34_27=0
.ic qb_34_27=1.8
.ic q_35_27=0
.ic qb_35_27=1.8
.ic q_36_27=0
.ic qb_36_27=1.8
.ic q_37_27=0
.ic qb_37_27=1.8
.ic q_38_27=0
.ic qb_38_27=1.8
.ic q_39_27=0
.ic qb_39_27=1.8
.ic q_40_27=0
.ic qb_40_27=1.8
.ic q_41_27=0
.ic qb_41_27=1.8
.ic q_42_27=0
.ic qb_42_27=1.8
.ic q_43_27=0
.ic qb_43_27=1.8
.ic q_44_27=0
.ic qb_44_27=1.8
.ic q_45_27=0
.ic qb_45_27=1.8
.ic q_46_27=0
.ic qb_46_27=1.8
.ic q_47_27=0
.ic qb_47_27=1.8
.ic q_48_27=0
.ic qb_48_27=1.8
.ic q_49_27=0
.ic qb_49_27=1.8
.ic q_50_27=0
.ic qb_50_27=1.8
.ic q_51_27=0
.ic qb_51_27=1.8
.ic q_52_27=0
.ic qb_52_27=1.8
.ic q_53_27=0
.ic qb_53_27=1.8
.ic q_54_27=0
.ic qb_54_27=1.8
.ic q_55_27=0
.ic qb_55_27=1.8
.ic q_56_27=0
.ic qb_56_27=1.8
.ic q_57_27=0
.ic qb_57_27=1.8
.ic q_58_27=0
.ic qb_58_27=1.8
.ic q_59_27=0
.ic qb_59_27=1.8
.ic q_60_27=0
.ic qb_60_27=1.8
.ic q_61_27=0
.ic qb_61_27=1.8
.ic q_62_27=0
.ic qb_62_27=1.8
.ic q_63_27=0
.ic qb_63_27=1.8
.ic q_64_27=0
.ic qb_64_27=1.8
.ic q_65_27=0
.ic qb_65_27=1.8
.ic q_66_27=0
.ic qb_66_27=1.8
.ic q_67_27=0
.ic qb_67_27=1.8
.ic q_68_27=0
.ic qb_68_27=1.8
.ic q_69_27=0
.ic qb_69_27=1.8
.ic q_70_27=0
.ic qb_70_27=1.8
.ic q_71_27=0
.ic qb_71_27=1.8
.ic q_72_27=0
.ic qb_72_27=1.8
.ic q_73_27=0
.ic qb_73_27=1.8
.ic q_74_27=0
.ic qb_74_27=1.8
.ic q_75_27=0
.ic qb_75_27=1.8
.ic q_76_27=0
.ic qb_76_27=1.8
.ic q_77_27=0
.ic qb_77_27=1.8
.ic q_78_27=0
.ic qb_78_27=1.8
.ic q_79_27=0
.ic qb_79_27=1.8
.ic q_80_27=0
.ic qb_80_27=1.8
.ic q_81_27=0
.ic qb_81_27=1.8
.ic q_82_27=0
.ic qb_82_27=1.8
.ic q_83_27=0
.ic qb_83_27=1.8
.ic q_84_27=0
.ic qb_84_27=1.8
.ic q_85_27=0
.ic qb_85_27=1.8
.ic q_86_27=0
.ic qb_86_27=1.8
.ic q_87_27=0
.ic qb_87_27=1.8
.ic q_88_27=0
.ic qb_88_27=1.8
.ic q_89_27=0
.ic qb_89_27=1.8
.ic q_90_27=0
.ic qb_90_27=1.8
.ic q_91_27=0
.ic qb_91_27=1.8
.ic q_92_27=0
.ic qb_92_27=1.8
.ic q_93_27=0
.ic qb_93_27=1.8
.ic q_94_27=0
.ic qb_94_27=1.8
.ic q_95_27=0
.ic qb_95_27=1.8
.ic q_96_27=0
.ic qb_96_27=1.8
.ic q_97_27=0
.ic qb_97_27=1.8
.ic q_98_27=0
.ic qb_98_27=1.8
.ic q_99_27=0
.ic qb_99_27=1.8
.ic q_0_28=0
.ic qb_0_28=1.8
.ic q_1_28=0
.ic qb_1_28=1.8
.ic q_2_28=0
.ic qb_2_28=1.8
.ic q_3_28=0
.ic qb_3_28=1.8
.ic q_4_28=0
.ic qb_4_28=1.8
.ic q_5_28=0
.ic qb_5_28=1.8
.ic q_6_28=0
.ic qb_6_28=1.8
.ic q_7_28=0
.ic qb_7_28=1.8
.ic q_8_28=0
.ic qb_8_28=1.8
.ic q_9_28=0
.ic qb_9_28=1.8
.ic q_10_28=0
.ic qb_10_28=1.8
.ic q_11_28=0
.ic qb_11_28=1.8
.ic q_12_28=0
.ic qb_12_28=1.8
.ic q_13_28=0
.ic qb_13_28=1.8
.ic q_14_28=0
.ic qb_14_28=1.8
.ic q_15_28=0
.ic qb_15_28=1.8
.ic q_16_28=0
.ic qb_16_28=1.8
.ic q_17_28=0
.ic qb_17_28=1.8
.ic q_18_28=0
.ic qb_18_28=1.8
.ic q_19_28=0
.ic qb_19_28=1.8
.ic q_20_28=0
.ic qb_20_28=1.8
.ic q_21_28=0
.ic qb_21_28=1.8
.ic q_22_28=0
.ic qb_22_28=1.8
.ic q_23_28=0
.ic qb_23_28=1.8
.ic q_24_28=0
.ic qb_24_28=1.8
.ic q_25_28=0
.ic qb_25_28=1.8
.ic q_26_28=0
.ic qb_26_28=1.8
.ic q_27_28=0
.ic qb_27_28=1.8
.ic q_28_28=0
.ic qb_28_28=1.8
.ic q_29_28=0
.ic qb_29_28=1.8
.ic q_30_28=0
.ic qb_30_28=1.8
.ic q_31_28=0
.ic qb_31_28=1.8
.ic q_32_28=0
.ic qb_32_28=1.8
.ic q_33_28=0
.ic qb_33_28=1.8
.ic q_34_28=0
.ic qb_34_28=1.8
.ic q_35_28=0
.ic qb_35_28=1.8
.ic q_36_28=0
.ic qb_36_28=1.8
.ic q_37_28=0
.ic qb_37_28=1.8
.ic q_38_28=0
.ic qb_38_28=1.8
.ic q_39_28=0
.ic qb_39_28=1.8
.ic q_40_28=0
.ic qb_40_28=1.8
.ic q_41_28=0
.ic qb_41_28=1.8
.ic q_42_28=0
.ic qb_42_28=1.8
.ic q_43_28=0
.ic qb_43_28=1.8
.ic q_44_28=0
.ic qb_44_28=1.8
.ic q_45_28=0
.ic qb_45_28=1.8
.ic q_46_28=0
.ic qb_46_28=1.8
.ic q_47_28=0
.ic qb_47_28=1.8
.ic q_48_28=0
.ic qb_48_28=1.8
.ic q_49_28=0
.ic qb_49_28=1.8
.ic q_50_28=0
.ic qb_50_28=1.8
.ic q_51_28=0
.ic qb_51_28=1.8
.ic q_52_28=0
.ic qb_52_28=1.8
.ic q_53_28=0
.ic qb_53_28=1.8
.ic q_54_28=0
.ic qb_54_28=1.8
.ic q_55_28=0
.ic qb_55_28=1.8
.ic q_56_28=0
.ic qb_56_28=1.8
.ic q_57_28=0
.ic qb_57_28=1.8
.ic q_58_28=0
.ic qb_58_28=1.8
.ic q_59_28=0
.ic qb_59_28=1.8
.ic q_60_28=0
.ic qb_60_28=1.8
.ic q_61_28=0
.ic qb_61_28=1.8
.ic q_62_28=0
.ic qb_62_28=1.8
.ic q_63_28=0
.ic qb_63_28=1.8
.ic q_64_28=0
.ic qb_64_28=1.8
.ic q_65_28=0
.ic qb_65_28=1.8
.ic q_66_28=0
.ic qb_66_28=1.8
.ic q_67_28=0
.ic qb_67_28=1.8
.ic q_68_28=0
.ic qb_68_28=1.8
.ic q_69_28=0
.ic qb_69_28=1.8
.ic q_70_28=0
.ic qb_70_28=1.8
.ic q_71_28=0
.ic qb_71_28=1.8
.ic q_72_28=0
.ic qb_72_28=1.8
.ic q_73_28=0
.ic qb_73_28=1.8
.ic q_74_28=0
.ic qb_74_28=1.8
.ic q_75_28=0
.ic qb_75_28=1.8
.ic q_76_28=0
.ic qb_76_28=1.8
.ic q_77_28=0
.ic qb_77_28=1.8
.ic q_78_28=0
.ic qb_78_28=1.8
.ic q_79_28=0
.ic qb_79_28=1.8
.ic q_80_28=0
.ic qb_80_28=1.8
.ic q_81_28=0
.ic qb_81_28=1.8
.ic q_82_28=0
.ic qb_82_28=1.8
.ic q_83_28=0
.ic qb_83_28=1.8
.ic q_84_28=0
.ic qb_84_28=1.8
.ic q_85_28=0
.ic qb_85_28=1.8
.ic q_86_28=0
.ic qb_86_28=1.8
.ic q_87_28=0
.ic qb_87_28=1.8
.ic q_88_28=0
.ic qb_88_28=1.8
.ic q_89_28=0
.ic qb_89_28=1.8
.ic q_90_28=0
.ic qb_90_28=1.8
.ic q_91_28=0
.ic qb_91_28=1.8
.ic q_92_28=0
.ic qb_92_28=1.8
.ic q_93_28=0
.ic qb_93_28=1.8
.ic q_94_28=0
.ic qb_94_28=1.8
.ic q_95_28=0
.ic qb_95_28=1.8
.ic q_96_28=0
.ic qb_96_28=1.8
.ic q_97_28=0
.ic qb_97_28=1.8
.ic q_98_28=0
.ic qb_98_28=1.8
.ic q_99_28=0
.ic qb_99_28=1.8
.ic q_0_29=0
.ic qb_0_29=1.8
.ic q_1_29=0
.ic qb_1_29=1.8
.ic q_2_29=0
.ic qb_2_29=1.8
.ic q_3_29=0
.ic qb_3_29=1.8
.ic q_4_29=0
.ic qb_4_29=1.8
.ic q_5_29=0
.ic qb_5_29=1.8
.ic q_6_29=0
.ic qb_6_29=1.8
.ic q_7_29=0
.ic qb_7_29=1.8
.ic q_8_29=0
.ic qb_8_29=1.8
.ic q_9_29=0
.ic qb_9_29=1.8
.ic q_10_29=0
.ic qb_10_29=1.8
.ic q_11_29=0
.ic qb_11_29=1.8
.ic q_12_29=0
.ic qb_12_29=1.8
.ic q_13_29=0
.ic qb_13_29=1.8
.ic q_14_29=0
.ic qb_14_29=1.8
.ic q_15_29=0
.ic qb_15_29=1.8
.ic q_16_29=0
.ic qb_16_29=1.8
.ic q_17_29=0
.ic qb_17_29=1.8
.ic q_18_29=0
.ic qb_18_29=1.8
.ic q_19_29=0
.ic qb_19_29=1.8
.ic q_20_29=0
.ic qb_20_29=1.8
.ic q_21_29=0
.ic qb_21_29=1.8
.ic q_22_29=0
.ic qb_22_29=1.8
.ic q_23_29=0
.ic qb_23_29=1.8
.ic q_24_29=0
.ic qb_24_29=1.8
.ic q_25_29=0
.ic qb_25_29=1.8
.ic q_26_29=0
.ic qb_26_29=1.8
.ic q_27_29=0
.ic qb_27_29=1.8
.ic q_28_29=0
.ic qb_28_29=1.8
.ic q_29_29=0
.ic qb_29_29=1.8
.ic q_30_29=0
.ic qb_30_29=1.8
.ic q_31_29=0
.ic qb_31_29=1.8
.ic q_32_29=0
.ic qb_32_29=1.8
.ic q_33_29=0
.ic qb_33_29=1.8
.ic q_34_29=0
.ic qb_34_29=1.8
.ic q_35_29=0
.ic qb_35_29=1.8
.ic q_36_29=0
.ic qb_36_29=1.8
.ic q_37_29=0
.ic qb_37_29=1.8
.ic q_38_29=0
.ic qb_38_29=1.8
.ic q_39_29=0
.ic qb_39_29=1.8
.ic q_40_29=0
.ic qb_40_29=1.8
.ic q_41_29=0
.ic qb_41_29=1.8
.ic q_42_29=0
.ic qb_42_29=1.8
.ic q_43_29=0
.ic qb_43_29=1.8
.ic q_44_29=0
.ic qb_44_29=1.8
.ic q_45_29=0
.ic qb_45_29=1.8
.ic q_46_29=0
.ic qb_46_29=1.8
.ic q_47_29=0
.ic qb_47_29=1.8
.ic q_48_29=0
.ic qb_48_29=1.8
.ic q_49_29=0
.ic qb_49_29=1.8
.ic q_50_29=0
.ic qb_50_29=1.8
.ic q_51_29=0
.ic qb_51_29=1.8
.ic q_52_29=0
.ic qb_52_29=1.8
.ic q_53_29=0
.ic qb_53_29=1.8
.ic q_54_29=0
.ic qb_54_29=1.8
.ic q_55_29=0
.ic qb_55_29=1.8
.ic q_56_29=0
.ic qb_56_29=1.8
.ic q_57_29=0
.ic qb_57_29=1.8
.ic q_58_29=0
.ic qb_58_29=1.8
.ic q_59_29=0
.ic qb_59_29=1.8
.ic q_60_29=0
.ic qb_60_29=1.8
.ic q_61_29=0
.ic qb_61_29=1.8
.ic q_62_29=0
.ic qb_62_29=1.8
.ic q_63_29=0
.ic qb_63_29=1.8
.ic q_64_29=0
.ic qb_64_29=1.8
.ic q_65_29=0
.ic qb_65_29=1.8
.ic q_66_29=0
.ic qb_66_29=1.8
.ic q_67_29=0
.ic qb_67_29=1.8
.ic q_68_29=0
.ic qb_68_29=1.8
.ic q_69_29=0
.ic qb_69_29=1.8
.ic q_70_29=0
.ic qb_70_29=1.8
.ic q_71_29=0
.ic qb_71_29=1.8
.ic q_72_29=0
.ic qb_72_29=1.8
.ic q_73_29=0
.ic qb_73_29=1.8
.ic q_74_29=0
.ic qb_74_29=1.8
.ic q_75_29=0
.ic qb_75_29=1.8
.ic q_76_29=0
.ic qb_76_29=1.8
.ic q_77_29=0
.ic qb_77_29=1.8
.ic q_78_29=0
.ic qb_78_29=1.8
.ic q_79_29=0
.ic qb_79_29=1.8
.ic q_80_29=0
.ic qb_80_29=1.8
.ic q_81_29=0
.ic qb_81_29=1.8
.ic q_82_29=0
.ic qb_82_29=1.8
.ic q_83_29=0
.ic qb_83_29=1.8
.ic q_84_29=0
.ic qb_84_29=1.8
.ic q_85_29=0
.ic qb_85_29=1.8
.ic q_86_29=0
.ic qb_86_29=1.8
.ic q_87_29=0
.ic qb_87_29=1.8
.ic q_88_29=0
.ic qb_88_29=1.8
.ic q_89_29=0
.ic qb_89_29=1.8
.ic q_90_29=0
.ic qb_90_29=1.8
.ic q_91_29=0
.ic qb_91_29=1.8
.ic q_92_29=0
.ic qb_92_29=1.8
.ic q_93_29=0
.ic qb_93_29=1.8
.ic q_94_29=0
.ic qb_94_29=1.8
.ic q_95_29=0
.ic qb_95_29=1.8
.ic q_96_29=0
.ic qb_96_29=1.8
.ic q_97_29=0
.ic qb_97_29=1.8
.ic q_98_29=0
.ic qb_98_29=1.8
.ic q_99_29=0
.ic qb_99_29=1.8
.ic q_0_30=0
.ic qb_0_30=1.8
.ic q_1_30=0
.ic qb_1_30=1.8
.ic q_2_30=0
.ic qb_2_30=1.8
.ic q_3_30=0
.ic qb_3_30=1.8
.ic q_4_30=0
.ic qb_4_30=1.8
.ic q_5_30=0
.ic qb_5_30=1.8
.ic q_6_30=0
.ic qb_6_30=1.8
.ic q_7_30=0
.ic qb_7_30=1.8
.ic q_8_30=0
.ic qb_8_30=1.8
.ic q_9_30=0
.ic qb_9_30=1.8
.ic q_10_30=0
.ic qb_10_30=1.8
.ic q_11_30=0
.ic qb_11_30=1.8
.ic q_12_30=0
.ic qb_12_30=1.8
.ic q_13_30=0
.ic qb_13_30=1.8
.ic q_14_30=0
.ic qb_14_30=1.8
.ic q_15_30=0
.ic qb_15_30=1.8
.ic q_16_30=0
.ic qb_16_30=1.8
.ic q_17_30=0
.ic qb_17_30=1.8
.ic q_18_30=0
.ic qb_18_30=1.8
.ic q_19_30=0
.ic qb_19_30=1.8
.ic q_20_30=0
.ic qb_20_30=1.8
.ic q_21_30=0
.ic qb_21_30=1.8
.ic q_22_30=0
.ic qb_22_30=1.8
.ic q_23_30=0
.ic qb_23_30=1.8
.ic q_24_30=0
.ic qb_24_30=1.8
.ic q_25_30=0
.ic qb_25_30=1.8
.ic q_26_30=0
.ic qb_26_30=1.8
.ic q_27_30=0
.ic qb_27_30=1.8
.ic q_28_30=0
.ic qb_28_30=1.8
.ic q_29_30=0
.ic qb_29_30=1.8
.ic q_30_30=0
.ic qb_30_30=1.8
.ic q_31_30=0
.ic qb_31_30=1.8
.ic q_32_30=0
.ic qb_32_30=1.8
.ic q_33_30=0
.ic qb_33_30=1.8
.ic q_34_30=0
.ic qb_34_30=1.8
.ic q_35_30=0
.ic qb_35_30=1.8
.ic q_36_30=0
.ic qb_36_30=1.8
.ic q_37_30=0
.ic qb_37_30=1.8
.ic q_38_30=0
.ic qb_38_30=1.8
.ic q_39_30=0
.ic qb_39_30=1.8
.ic q_40_30=0
.ic qb_40_30=1.8
.ic q_41_30=0
.ic qb_41_30=1.8
.ic q_42_30=0
.ic qb_42_30=1.8
.ic q_43_30=0
.ic qb_43_30=1.8
.ic q_44_30=0
.ic qb_44_30=1.8
.ic q_45_30=0
.ic qb_45_30=1.8
.ic q_46_30=0
.ic qb_46_30=1.8
.ic q_47_30=0
.ic qb_47_30=1.8
.ic q_48_30=0
.ic qb_48_30=1.8
.ic q_49_30=0
.ic qb_49_30=1.8
.ic q_50_30=0
.ic qb_50_30=1.8
.ic q_51_30=0
.ic qb_51_30=1.8
.ic q_52_30=0
.ic qb_52_30=1.8
.ic q_53_30=0
.ic qb_53_30=1.8
.ic q_54_30=0
.ic qb_54_30=1.8
.ic q_55_30=0
.ic qb_55_30=1.8
.ic q_56_30=0
.ic qb_56_30=1.8
.ic q_57_30=0
.ic qb_57_30=1.8
.ic q_58_30=0
.ic qb_58_30=1.8
.ic q_59_30=0
.ic qb_59_30=1.8
.ic q_60_30=0
.ic qb_60_30=1.8
.ic q_61_30=0
.ic qb_61_30=1.8
.ic q_62_30=0
.ic qb_62_30=1.8
.ic q_63_30=0
.ic qb_63_30=1.8
.ic q_64_30=0
.ic qb_64_30=1.8
.ic q_65_30=0
.ic qb_65_30=1.8
.ic q_66_30=0
.ic qb_66_30=1.8
.ic q_67_30=0
.ic qb_67_30=1.8
.ic q_68_30=0
.ic qb_68_30=1.8
.ic q_69_30=0
.ic qb_69_30=1.8
.ic q_70_30=0
.ic qb_70_30=1.8
.ic q_71_30=0
.ic qb_71_30=1.8
.ic q_72_30=0
.ic qb_72_30=1.8
.ic q_73_30=0
.ic qb_73_30=1.8
.ic q_74_30=0
.ic qb_74_30=1.8
.ic q_75_30=0
.ic qb_75_30=1.8
.ic q_76_30=0
.ic qb_76_30=1.8
.ic q_77_30=0
.ic qb_77_30=1.8
.ic q_78_30=0
.ic qb_78_30=1.8
.ic q_79_30=0
.ic qb_79_30=1.8
.ic q_80_30=0
.ic qb_80_30=1.8
.ic q_81_30=0
.ic qb_81_30=1.8
.ic q_82_30=0
.ic qb_82_30=1.8
.ic q_83_30=0
.ic qb_83_30=1.8
.ic q_84_30=0
.ic qb_84_30=1.8
.ic q_85_30=0
.ic qb_85_30=1.8
.ic q_86_30=0
.ic qb_86_30=1.8
.ic q_87_30=0
.ic qb_87_30=1.8
.ic q_88_30=0
.ic qb_88_30=1.8
.ic q_89_30=0
.ic qb_89_30=1.8
.ic q_90_30=0
.ic qb_90_30=1.8
.ic q_91_30=0
.ic qb_91_30=1.8
.ic q_92_30=0
.ic qb_92_30=1.8
.ic q_93_30=0
.ic qb_93_30=1.8
.ic q_94_30=0
.ic qb_94_30=1.8
.ic q_95_30=0
.ic qb_95_30=1.8
.ic q_96_30=0
.ic qb_96_30=1.8
.ic q_97_30=0
.ic qb_97_30=1.8
.ic q_98_30=0
.ic qb_98_30=1.8
.ic q_99_30=0
.ic qb_99_30=1.8
.ic q_0_31=0
.ic qb_0_31=1.8
.ic q_1_31=0
.ic qb_1_31=1.8
.ic q_2_31=0
.ic qb_2_31=1.8
.ic q_3_31=0
.ic qb_3_31=1.8
.ic q_4_31=0
.ic qb_4_31=1.8
.ic q_5_31=0
.ic qb_5_31=1.8
.ic q_6_31=0
.ic qb_6_31=1.8
.ic q_7_31=0
.ic qb_7_31=1.8
.ic q_8_31=0
.ic qb_8_31=1.8
.ic q_9_31=0
.ic qb_9_31=1.8
.ic q_10_31=0
.ic qb_10_31=1.8
.ic q_11_31=0
.ic qb_11_31=1.8
.ic q_12_31=0
.ic qb_12_31=1.8
.ic q_13_31=0
.ic qb_13_31=1.8
.ic q_14_31=0
.ic qb_14_31=1.8
.ic q_15_31=0
.ic qb_15_31=1.8
.ic q_16_31=0
.ic qb_16_31=1.8
.ic q_17_31=0
.ic qb_17_31=1.8
.ic q_18_31=0
.ic qb_18_31=1.8
.ic q_19_31=0
.ic qb_19_31=1.8
.ic q_20_31=0
.ic qb_20_31=1.8
.ic q_21_31=0
.ic qb_21_31=1.8
.ic q_22_31=0
.ic qb_22_31=1.8
.ic q_23_31=0
.ic qb_23_31=1.8
.ic q_24_31=0
.ic qb_24_31=1.8
.ic q_25_31=0
.ic qb_25_31=1.8
.ic q_26_31=0
.ic qb_26_31=1.8
.ic q_27_31=0
.ic qb_27_31=1.8
.ic q_28_31=0
.ic qb_28_31=1.8
.ic q_29_31=0
.ic qb_29_31=1.8
.ic q_30_31=0
.ic qb_30_31=1.8
.ic q_31_31=0
.ic qb_31_31=1.8
.ic q_32_31=0
.ic qb_32_31=1.8
.ic q_33_31=0
.ic qb_33_31=1.8
.ic q_34_31=0
.ic qb_34_31=1.8
.ic q_35_31=0
.ic qb_35_31=1.8
.ic q_36_31=0
.ic qb_36_31=1.8
.ic q_37_31=0
.ic qb_37_31=1.8
.ic q_38_31=0
.ic qb_38_31=1.8
.ic q_39_31=0
.ic qb_39_31=1.8
.ic q_40_31=0
.ic qb_40_31=1.8
.ic q_41_31=0
.ic qb_41_31=1.8
.ic q_42_31=0
.ic qb_42_31=1.8
.ic q_43_31=0
.ic qb_43_31=1.8
.ic q_44_31=0
.ic qb_44_31=1.8
.ic q_45_31=0
.ic qb_45_31=1.8
.ic q_46_31=0
.ic qb_46_31=1.8
.ic q_47_31=0
.ic qb_47_31=1.8
.ic q_48_31=0
.ic qb_48_31=1.8
.ic q_49_31=0
.ic qb_49_31=1.8
.ic q_50_31=0
.ic qb_50_31=1.8
.ic q_51_31=0
.ic qb_51_31=1.8
.ic q_52_31=0
.ic qb_52_31=1.8
.ic q_53_31=0
.ic qb_53_31=1.8
.ic q_54_31=0
.ic qb_54_31=1.8
.ic q_55_31=0
.ic qb_55_31=1.8
.ic q_56_31=0
.ic qb_56_31=1.8
.ic q_57_31=0
.ic qb_57_31=1.8
.ic q_58_31=0
.ic qb_58_31=1.8
.ic q_59_31=0
.ic qb_59_31=1.8
.ic q_60_31=0
.ic qb_60_31=1.8
.ic q_61_31=0
.ic qb_61_31=1.8
.ic q_62_31=0
.ic qb_62_31=1.8
.ic q_63_31=0
.ic qb_63_31=1.8
.ic q_64_31=0
.ic qb_64_31=1.8
.ic q_65_31=0
.ic qb_65_31=1.8
.ic q_66_31=0
.ic qb_66_31=1.8
.ic q_67_31=0
.ic qb_67_31=1.8
.ic q_68_31=0
.ic qb_68_31=1.8
.ic q_69_31=0
.ic qb_69_31=1.8
.ic q_70_31=0
.ic qb_70_31=1.8
.ic q_71_31=0
.ic qb_71_31=1.8
.ic q_72_31=0
.ic qb_72_31=1.8
.ic q_73_31=0
.ic qb_73_31=1.8
.ic q_74_31=0
.ic qb_74_31=1.8
.ic q_75_31=0
.ic qb_75_31=1.8
.ic q_76_31=0
.ic qb_76_31=1.8
.ic q_77_31=0
.ic qb_77_31=1.8
.ic q_78_31=0
.ic qb_78_31=1.8
.ic q_79_31=0
.ic qb_79_31=1.8
.ic q_80_31=0
.ic qb_80_31=1.8
.ic q_81_31=0
.ic qb_81_31=1.8
.ic q_82_31=0
.ic qb_82_31=1.8
.ic q_83_31=0
.ic qb_83_31=1.8
.ic q_84_31=0
.ic qb_84_31=1.8
.ic q_85_31=0
.ic qb_85_31=1.8
.ic q_86_31=0
.ic qb_86_31=1.8
.ic q_87_31=0
.ic qb_87_31=1.8
.ic q_88_31=0
.ic qb_88_31=1.8
.ic q_89_31=0
.ic qb_89_31=1.8
.ic q_90_31=0
.ic qb_90_31=1.8
.ic q_91_31=0
.ic qb_91_31=1.8
.ic q_92_31=0
.ic qb_92_31=1.8
.ic q_93_31=0
.ic qb_93_31=1.8
.ic q_94_31=0
.ic qb_94_31=1.8
.ic q_95_31=0
.ic qb_95_31=1.8
.ic q_96_31=0
.ic qb_96_31=1.8
.ic q_97_31=0
.ic qb_97_31=1.8
.ic q_98_31=0
.ic qb_98_31=1.8
.ic q_99_31=0
.ic qb_99_31=1.8
.ic q_0_32=0
.ic qb_0_32=1.8
.ic q_1_32=0
.ic qb_1_32=1.8
.ic q_2_32=0
.ic qb_2_32=1.8
.ic q_3_32=0
.ic qb_3_32=1.8
.ic q_4_32=0
.ic qb_4_32=1.8
.ic q_5_32=0
.ic qb_5_32=1.8
.ic q_6_32=0
.ic qb_6_32=1.8
.ic q_7_32=0
.ic qb_7_32=1.8
.ic q_8_32=0
.ic qb_8_32=1.8
.ic q_9_32=0
.ic qb_9_32=1.8
.ic q_10_32=0
.ic qb_10_32=1.8
.ic q_11_32=0
.ic qb_11_32=1.8
.ic q_12_32=0
.ic qb_12_32=1.8
.ic q_13_32=0
.ic qb_13_32=1.8
.ic q_14_32=0
.ic qb_14_32=1.8
.ic q_15_32=0
.ic qb_15_32=1.8
.ic q_16_32=0
.ic qb_16_32=1.8
.ic q_17_32=0
.ic qb_17_32=1.8
.ic q_18_32=0
.ic qb_18_32=1.8
.ic q_19_32=0
.ic qb_19_32=1.8
.ic q_20_32=0
.ic qb_20_32=1.8
.ic q_21_32=0
.ic qb_21_32=1.8
.ic q_22_32=0
.ic qb_22_32=1.8
.ic q_23_32=0
.ic qb_23_32=1.8
.ic q_24_32=0
.ic qb_24_32=1.8
.ic q_25_32=0
.ic qb_25_32=1.8
.ic q_26_32=0
.ic qb_26_32=1.8
.ic q_27_32=0
.ic qb_27_32=1.8
.ic q_28_32=0
.ic qb_28_32=1.8
.ic q_29_32=0
.ic qb_29_32=1.8
.ic q_30_32=0
.ic qb_30_32=1.8
.ic q_31_32=0
.ic qb_31_32=1.8
.ic q_32_32=0
.ic qb_32_32=1.8
.ic q_33_32=0
.ic qb_33_32=1.8
.ic q_34_32=0
.ic qb_34_32=1.8
.ic q_35_32=0
.ic qb_35_32=1.8
.ic q_36_32=0
.ic qb_36_32=1.8
.ic q_37_32=0
.ic qb_37_32=1.8
.ic q_38_32=0
.ic qb_38_32=1.8
.ic q_39_32=0
.ic qb_39_32=1.8
.ic q_40_32=0
.ic qb_40_32=1.8
.ic q_41_32=0
.ic qb_41_32=1.8
.ic q_42_32=0
.ic qb_42_32=1.8
.ic q_43_32=0
.ic qb_43_32=1.8
.ic q_44_32=0
.ic qb_44_32=1.8
.ic q_45_32=0
.ic qb_45_32=1.8
.ic q_46_32=0
.ic qb_46_32=1.8
.ic q_47_32=0
.ic qb_47_32=1.8
.ic q_48_32=0
.ic qb_48_32=1.8
.ic q_49_32=0
.ic qb_49_32=1.8
.ic q_50_32=0
.ic qb_50_32=1.8
.ic q_51_32=0
.ic qb_51_32=1.8
.ic q_52_32=0
.ic qb_52_32=1.8
.ic q_53_32=0
.ic qb_53_32=1.8
.ic q_54_32=0
.ic qb_54_32=1.8
.ic q_55_32=0
.ic qb_55_32=1.8
.ic q_56_32=0
.ic qb_56_32=1.8
.ic q_57_32=0
.ic qb_57_32=1.8
.ic q_58_32=0
.ic qb_58_32=1.8
.ic q_59_32=0
.ic qb_59_32=1.8
.ic q_60_32=0
.ic qb_60_32=1.8
.ic q_61_32=0
.ic qb_61_32=1.8
.ic q_62_32=0
.ic qb_62_32=1.8
.ic q_63_32=0
.ic qb_63_32=1.8
.ic q_64_32=0
.ic qb_64_32=1.8
.ic q_65_32=0
.ic qb_65_32=1.8
.ic q_66_32=0
.ic qb_66_32=1.8
.ic q_67_32=0
.ic qb_67_32=1.8
.ic q_68_32=0
.ic qb_68_32=1.8
.ic q_69_32=0
.ic qb_69_32=1.8
.ic q_70_32=0
.ic qb_70_32=1.8
.ic q_71_32=0
.ic qb_71_32=1.8
.ic q_72_32=0
.ic qb_72_32=1.8
.ic q_73_32=0
.ic qb_73_32=1.8
.ic q_74_32=0
.ic qb_74_32=1.8
.ic q_75_32=0
.ic qb_75_32=1.8
.ic q_76_32=0
.ic qb_76_32=1.8
.ic q_77_32=0
.ic qb_77_32=1.8
.ic q_78_32=0
.ic qb_78_32=1.8
.ic q_79_32=0
.ic qb_79_32=1.8
.ic q_80_32=0
.ic qb_80_32=1.8
.ic q_81_32=0
.ic qb_81_32=1.8
.ic q_82_32=0
.ic qb_82_32=1.8
.ic q_83_32=0
.ic qb_83_32=1.8
.ic q_84_32=0
.ic qb_84_32=1.8
.ic q_85_32=0
.ic qb_85_32=1.8
.ic q_86_32=0
.ic qb_86_32=1.8
.ic q_87_32=0
.ic qb_87_32=1.8
.ic q_88_32=0
.ic qb_88_32=1.8
.ic q_89_32=0
.ic qb_89_32=1.8
.ic q_90_32=0
.ic qb_90_32=1.8
.ic q_91_32=0
.ic qb_91_32=1.8
.ic q_92_32=0
.ic qb_92_32=1.8
.ic q_93_32=0
.ic qb_93_32=1.8
.ic q_94_32=0
.ic qb_94_32=1.8
.ic q_95_32=0
.ic qb_95_32=1.8
.ic q_96_32=0
.ic qb_96_32=1.8
.ic q_97_32=0
.ic qb_97_32=1.8
.ic q_98_32=0
.ic qb_98_32=1.8
.ic q_99_32=0
.ic qb_99_32=1.8
.ic q_0_33=0
.ic qb_0_33=1.8
.ic q_1_33=0
.ic qb_1_33=1.8
.ic q_2_33=0
.ic qb_2_33=1.8
.ic q_3_33=0
.ic qb_3_33=1.8
.ic q_4_33=0
.ic qb_4_33=1.8
.ic q_5_33=0
.ic qb_5_33=1.8
.ic q_6_33=0
.ic qb_6_33=1.8
.ic q_7_33=0
.ic qb_7_33=1.8
.ic q_8_33=0
.ic qb_8_33=1.8
.ic q_9_33=0
.ic qb_9_33=1.8
.ic q_10_33=0
.ic qb_10_33=1.8
.ic q_11_33=0
.ic qb_11_33=1.8
.ic q_12_33=0
.ic qb_12_33=1.8
.ic q_13_33=0
.ic qb_13_33=1.8
.ic q_14_33=0
.ic qb_14_33=1.8
.ic q_15_33=0
.ic qb_15_33=1.8
.ic q_16_33=0
.ic qb_16_33=1.8
.ic q_17_33=0
.ic qb_17_33=1.8
.ic q_18_33=0
.ic qb_18_33=1.8
.ic q_19_33=0
.ic qb_19_33=1.8
.ic q_20_33=0
.ic qb_20_33=1.8
.ic q_21_33=0
.ic qb_21_33=1.8
.ic q_22_33=0
.ic qb_22_33=1.8
.ic q_23_33=0
.ic qb_23_33=1.8
.ic q_24_33=0
.ic qb_24_33=1.8
.ic q_25_33=0
.ic qb_25_33=1.8
.ic q_26_33=0
.ic qb_26_33=1.8
.ic q_27_33=0
.ic qb_27_33=1.8
.ic q_28_33=0
.ic qb_28_33=1.8
.ic q_29_33=0
.ic qb_29_33=1.8
.ic q_30_33=0
.ic qb_30_33=1.8
.ic q_31_33=0
.ic qb_31_33=1.8
.ic q_32_33=0
.ic qb_32_33=1.8
.ic q_33_33=0
.ic qb_33_33=1.8
.ic q_34_33=0
.ic qb_34_33=1.8
.ic q_35_33=0
.ic qb_35_33=1.8
.ic q_36_33=0
.ic qb_36_33=1.8
.ic q_37_33=0
.ic qb_37_33=1.8
.ic q_38_33=0
.ic qb_38_33=1.8
.ic q_39_33=0
.ic qb_39_33=1.8
.ic q_40_33=0
.ic qb_40_33=1.8
.ic q_41_33=0
.ic qb_41_33=1.8
.ic q_42_33=0
.ic qb_42_33=1.8
.ic q_43_33=0
.ic qb_43_33=1.8
.ic q_44_33=0
.ic qb_44_33=1.8
.ic q_45_33=0
.ic qb_45_33=1.8
.ic q_46_33=0
.ic qb_46_33=1.8
.ic q_47_33=0
.ic qb_47_33=1.8
.ic q_48_33=0
.ic qb_48_33=1.8
.ic q_49_33=0
.ic qb_49_33=1.8
.ic q_50_33=0
.ic qb_50_33=1.8
.ic q_51_33=0
.ic qb_51_33=1.8
.ic q_52_33=0
.ic qb_52_33=1.8
.ic q_53_33=0
.ic qb_53_33=1.8
.ic q_54_33=0
.ic qb_54_33=1.8
.ic q_55_33=0
.ic qb_55_33=1.8
.ic q_56_33=0
.ic qb_56_33=1.8
.ic q_57_33=0
.ic qb_57_33=1.8
.ic q_58_33=0
.ic qb_58_33=1.8
.ic q_59_33=0
.ic qb_59_33=1.8
.ic q_60_33=0
.ic qb_60_33=1.8
.ic q_61_33=0
.ic qb_61_33=1.8
.ic q_62_33=0
.ic qb_62_33=1.8
.ic q_63_33=0
.ic qb_63_33=1.8
.ic q_64_33=0
.ic qb_64_33=1.8
.ic q_65_33=0
.ic qb_65_33=1.8
.ic q_66_33=0
.ic qb_66_33=1.8
.ic q_67_33=0
.ic qb_67_33=1.8
.ic q_68_33=0
.ic qb_68_33=1.8
.ic q_69_33=0
.ic qb_69_33=1.8
.ic q_70_33=0
.ic qb_70_33=1.8
.ic q_71_33=0
.ic qb_71_33=1.8
.ic q_72_33=0
.ic qb_72_33=1.8
.ic q_73_33=0
.ic qb_73_33=1.8
.ic q_74_33=0
.ic qb_74_33=1.8
.ic q_75_33=0
.ic qb_75_33=1.8
.ic q_76_33=0
.ic qb_76_33=1.8
.ic q_77_33=0
.ic qb_77_33=1.8
.ic q_78_33=0
.ic qb_78_33=1.8
.ic q_79_33=0
.ic qb_79_33=1.8
.ic q_80_33=0
.ic qb_80_33=1.8
.ic q_81_33=0
.ic qb_81_33=1.8
.ic q_82_33=0
.ic qb_82_33=1.8
.ic q_83_33=0
.ic qb_83_33=1.8
.ic q_84_33=0
.ic qb_84_33=1.8
.ic q_85_33=0
.ic qb_85_33=1.8
.ic q_86_33=0
.ic qb_86_33=1.8
.ic q_87_33=0
.ic qb_87_33=1.8
.ic q_88_33=0
.ic qb_88_33=1.8
.ic q_89_33=0
.ic qb_89_33=1.8
.ic q_90_33=0
.ic qb_90_33=1.8
.ic q_91_33=0
.ic qb_91_33=1.8
.ic q_92_33=0
.ic qb_92_33=1.8
.ic q_93_33=0
.ic qb_93_33=1.8
.ic q_94_33=0
.ic qb_94_33=1.8
.ic q_95_33=0
.ic qb_95_33=1.8
.ic q_96_33=0
.ic qb_96_33=1.8
.ic q_97_33=0
.ic qb_97_33=1.8
.ic q_98_33=0
.ic qb_98_33=1.8
.ic q_99_33=0
.ic qb_99_33=1.8
.ic q_0_34=0
.ic qb_0_34=1.8
.ic q_1_34=0
.ic qb_1_34=1.8
.ic q_2_34=0
.ic qb_2_34=1.8
.ic q_3_34=0
.ic qb_3_34=1.8
.ic q_4_34=0
.ic qb_4_34=1.8
.ic q_5_34=0
.ic qb_5_34=1.8
.ic q_6_34=0
.ic qb_6_34=1.8
.ic q_7_34=0
.ic qb_7_34=1.8
.ic q_8_34=0
.ic qb_8_34=1.8
.ic q_9_34=0
.ic qb_9_34=1.8
.ic q_10_34=0
.ic qb_10_34=1.8
.ic q_11_34=0
.ic qb_11_34=1.8
.ic q_12_34=0
.ic qb_12_34=1.8
.ic q_13_34=0
.ic qb_13_34=1.8
.ic q_14_34=0
.ic qb_14_34=1.8
.ic q_15_34=0
.ic qb_15_34=1.8
.ic q_16_34=0
.ic qb_16_34=1.8
.ic q_17_34=0
.ic qb_17_34=1.8
.ic q_18_34=0
.ic qb_18_34=1.8
.ic q_19_34=0
.ic qb_19_34=1.8
.ic q_20_34=0
.ic qb_20_34=1.8
.ic q_21_34=0
.ic qb_21_34=1.8
.ic q_22_34=0
.ic qb_22_34=1.8
.ic q_23_34=0
.ic qb_23_34=1.8
.ic q_24_34=0
.ic qb_24_34=1.8
.ic q_25_34=0
.ic qb_25_34=1.8
.ic q_26_34=0
.ic qb_26_34=1.8
.ic q_27_34=0
.ic qb_27_34=1.8
.ic q_28_34=0
.ic qb_28_34=1.8
.ic q_29_34=0
.ic qb_29_34=1.8
.ic q_30_34=0
.ic qb_30_34=1.8
.ic q_31_34=0
.ic qb_31_34=1.8
.ic q_32_34=0
.ic qb_32_34=1.8
.ic q_33_34=0
.ic qb_33_34=1.8
.ic q_34_34=0
.ic qb_34_34=1.8
.ic q_35_34=0
.ic qb_35_34=1.8
.ic q_36_34=0
.ic qb_36_34=1.8
.ic q_37_34=0
.ic qb_37_34=1.8
.ic q_38_34=0
.ic qb_38_34=1.8
.ic q_39_34=0
.ic qb_39_34=1.8
.ic q_40_34=0
.ic qb_40_34=1.8
.ic q_41_34=0
.ic qb_41_34=1.8
.ic q_42_34=0
.ic qb_42_34=1.8
.ic q_43_34=0
.ic qb_43_34=1.8
.ic q_44_34=0
.ic qb_44_34=1.8
.ic q_45_34=0
.ic qb_45_34=1.8
.ic q_46_34=0
.ic qb_46_34=1.8
.ic q_47_34=0
.ic qb_47_34=1.8
.ic q_48_34=0
.ic qb_48_34=1.8
.ic q_49_34=0
.ic qb_49_34=1.8
.ic q_50_34=0
.ic qb_50_34=1.8
.ic q_51_34=0
.ic qb_51_34=1.8
.ic q_52_34=0
.ic qb_52_34=1.8
.ic q_53_34=0
.ic qb_53_34=1.8
.ic q_54_34=0
.ic qb_54_34=1.8
.ic q_55_34=0
.ic qb_55_34=1.8
.ic q_56_34=0
.ic qb_56_34=1.8
.ic q_57_34=0
.ic qb_57_34=1.8
.ic q_58_34=0
.ic qb_58_34=1.8
.ic q_59_34=0
.ic qb_59_34=1.8
.ic q_60_34=0
.ic qb_60_34=1.8
.ic q_61_34=0
.ic qb_61_34=1.8
.ic q_62_34=0
.ic qb_62_34=1.8
.ic q_63_34=0
.ic qb_63_34=1.8
.ic q_64_34=0
.ic qb_64_34=1.8
.ic q_65_34=0
.ic qb_65_34=1.8
.ic q_66_34=0
.ic qb_66_34=1.8
.ic q_67_34=0
.ic qb_67_34=1.8
.ic q_68_34=0
.ic qb_68_34=1.8
.ic q_69_34=0
.ic qb_69_34=1.8
.ic q_70_34=0
.ic qb_70_34=1.8
.ic q_71_34=0
.ic qb_71_34=1.8
.ic q_72_34=0
.ic qb_72_34=1.8
.ic q_73_34=0
.ic qb_73_34=1.8
.ic q_74_34=0
.ic qb_74_34=1.8
.ic q_75_34=0
.ic qb_75_34=1.8
.ic q_76_34=0
.ic qb_76_34=1.8
.ic q_77_34=0
.ic qb_77_34=1.8
.ic q_78_34=0
.ic qb_78_34=1.8
.ic q_79_34=0
.ic qb_79_34=1.8
.ic q_80_34=0
.ic qb_80_34=1.8
.ic q_81_34=0
.ic qb_81_34=1.8
.ic q_82_34=0
.ic qb_82_34=1.8
.ic q_83_34=0
.ic qb_83_34=1.8
.ic q_84_34=0
.ic qb_84_34=1.8
.ic q_85_34=0
.ic qb_85_34=1.8
.ic q_86_34=0
.ic qb_86_34=1.8
.ic q_87_34=0
.ic qb_87_34=1.8
.ic q_88_34=0
.ic qb_88_34=1.8
.ic q_89_34=0
.ic qb_89_34=1.8
.ic q_90_34=0
.ic qb_90_34=1.8
.ic q_91_34=0
.ic qb_91_34=1.8
.ic q_92_34=0
.ic qb_92_34=1.8
.ic q_93_34=0
.ic qb_93_34=1.8
.ic q_94_34=0
.ic qb_94_34=1.8
.ic q_95_34=0
.ic qb_95_34=1.8
.ic q_96_34=0
.ic qb_96_34=1.8
.ic q_97_34=0
.ic qb_97_34=1.8
.ic q_98_34=0
.ic qb_98_34=1.8
.ic q_99_34=0
.ic qb_99_34=1.8
.ic q_0_35=0
.ic qb_0_35=1.8
.ic q_1_35=0
.ic qb_1_35=1.8
.ic q_2_35=0
.ic qb_2_35=1.8
.ic q_3_35=0
.ic qb_3_35=1.8
.ic q_4_35=0
.ic qb_4_35=1.8
.ic q_5_35=0
.ic qb_5_35=1.8
.ic q_6_35=0
.ic qb_6_35=1.8
.ic q_7_35=0
.ic qb_7_35=1.8
.ic q_8_35=0
.ic qb_8_35=1.8
.ic q_9_35=0
.ic qb_9_35=1.8
.ic q_10_35=0
.ic qb_10_35=1.8
.ic q_11_35=0
.ic qb_11_35=1.8
.ic q_12_35=0
.ic qb_12_35=1.8
.ic q_13_35=0
.ic qb_13_35=1.8
.ic q_14_35=0
.ic qb_14_35=1.8
.ic q_15_35=0
.ic qb_15_35=1.8
.ic q_16_35=0
.ic qb_16_35=1.8
.ic q_17_35=0
.ic qb_17_35=1.8
.ic q_18_35=0
.ic qb_18_35=1.8
.ic q_19_35=0
.ic qb_19_35=1.8
.ic q_20_35=0
.ic qb_20_35=1.8
.ic q_21_35=0
.ic qb_21_35=1.8
.ic q_22_35=0
.ic qb_22_35=1.8
.ic q_23_35=0
.ic qb_23_35=1.8
.ic q_24_35=0
.ic qb_24_35=1.8
.ic q_25_35=0
.ic qb_25_35=1.8
.ic q_26_35=0
.ic qb_26_35=1.8
.ic q_27_35=0
.ic qb_27_35=1.8
.ic q_28_35=0
.ic qb_28_35=1.8
.ic q_29_35=0
.ic qb_29_35=1.8
.ic q_30_35=0
.ic qb_30_35=1.8
.ic q_31_35=0
.ic qb_31_35=1.8
.ic q_32_35=0
.ic qb_32_35=1.8
.ic q_33_35=0
.ic qb_33_35=1.8
.ic q_34_35=0
.ic qb_34_35=1.8
.ic q_35_35=0
.ic qb_35_35=1.8
.ic q_36_35=0
.ic qb_36_35=1.8
.ic q_37_35=0
.ic qb_37_35=1.8
.ic q_38_35=0
.ic qb_38_35=1.8
.ic q_39_35=0
.ic qb_39_35=1.8
.ic q_40_35=0
.ic qb_40_35=1.8
.ic q_41_35=0
.ic qb_41_35=1.8
.ic q_42_35=0
.ic qb_42_35=1.8
.ic q_43_35=0
.ic qb_43_35=1.8
.ic q_44_35=0
.ic qb_44_35=1.8
.ic q_45_35=0
.ic qb_45_35=1.8
.ic q_46_35=0
.ic qb_46_35=1.8
.ic q_47_35=0
.ic qb_47_35=1.8
.ic q_48_35=0
.ic qb_48_35=1.8
.ic q_49_35=0
.ic qb_49_35=1.8
.ic q_50_35=0
.ic qb_50_35=1.8
.ic q_51_35=0
.ic qb_51_35=1.8
.ic q_52_35=0
.ic qb_52_35=1.8
.ic q_53_35=0
.ic qb_53_35=1.8
.ic q_54_35=0
.ic qb_54_35=1.8
.ic q_55_35=0
.ic qb_55_35=1.8
.ic q_56_35=0
.ic qb_56_35=1.8
.ic q_57_35=0
.ic qb_57_35=1.8
.ic q_58_35=0
.ic qb_58_35=1.8
.ic q_59_35=0
.ic qb_59_35=1.8
.ic q_60_35=0
.ic qb_60_35=1.8
.ic q_61_35=0
.ic qb_61_35=1.8
.ic q_62_35=0
.ic qb_62_35=1.8
.ic q_63_35=0
.ic qb_63_35=1.8
.ic q_64_35=0
.ic qb_64_35=1.8
.ic q_65_35=0
.ic qb_65_35=1.8
.ic q_66_35=0
.ic qb_66_35=1.8
.ic q_67_35=0
.ic qb_67_35=1.8
.ic q_68_35=0
.ic qb_68_35=1.8
.ic q_69_35=0
.ic qb_69_35=1.8
.ic q_70_35=0
.ic qb_70_35=1.8
.ic q_71_35=0
.ic qb_71_35=1.8
.ic q_72_35=0
.ic qb_72_35=1.8
.ic q_73_35=0
.ic qb_73_35=1.8
.ic q_74_35=0
.ic qb_74_35=1.8
.ic q_75_35=0
.ic qb_75_35=1.8
.ic q_76_35=0
.ic qb_76_35=1.8
.ic q_77_35=0
.ic qb_77_35=1.8
.ic q_78_35=0
.ic qb_78_35=1.8
.ic q_79_35=0
.ic qb_79_35=1.8
.ic q_80_35=0
.ic qb_80_35=1.8
.ic q_81_35=0
.ic qb_81_35=1.8
.ic q_82_35=0
.ic qb_82_35=1.8
.ic q_83_35=0
.ic qb_83_35=1.8
.ic q_84_35=0
.ic qb_84_35=1.8
.ic q_85_35=0
.ic qb_85_35=1.8
.ic q_86_35=0
.ic qb_86_35=1.8
.ic q_87_35=0
.ic qb_87_35=1.8
.ic q_88_35=0
.ic qb_88_35=1.8
.ic q_89_35=0
.ic qb_89_35=1.8
.ic q_90_35=0
.ic qb_90_35=1.8
.ic q_91_35=0
.ic qb_91_35=1.8
.ic q_92_35=0
.ic qb_92_35=1.8
.ic q_93_35=0
.ic qb_93_35=1.8
.ic q_94_35=0
.ic qb_94_35=1.8
.ic q_95_35=0
.ic qb_95_35=1.8
.ic q_96_35=0
.ic qb_96_35=1.8
.ic q_97_35=0
.ic qb_97_35=1.8
.ic q_98_35=0
.ic qb_98_35=1.8
.ic q_99_35=0
.ic qb_99_35=1.8
.ic q_0_36=0
.ic qb_0_36=1.8
.ic q_1_36=0
.ic qb_1_36=1.8
.ic q_2_36=0
.ic qb_2_36=1.8
.ic q_3_36=0
.ic qb_3_36=1.8
.ic q_4_36=0
.ic qb_4_36=1.8
.ic q_5_36=0
.ic qb_5_36=1.8
.ic q_6_36=0
.ic qb_6_36=1.8
.ic q_7_36=0
.ic qb_7_36=1.8
.ic q_8_36=0
.ic qb_8_36=1.8
.ic q_9_36=0
.ic qb_9_36=1.8
.ic q_10_36=0
.ic qb_10_36=1.8
.ic q_11_36=0
.ic qb_11_36=1.8
.ic q_12_36=0
.ic qb_12_36=1.8
.ic q_13_36=0
.ic qb_13_36=1.8
.ic q_14_36=0
.ic qb_14_36=1.8
.ic q_15_36=0
.ic qb_15_36=1.8
.ic q_16_36=0
.ic qb_16_36=1.8
.ic q_17_36=0
.ic qb_17_36=1.8
.ic q_18_36=0
.ic qb_18_36=1.8
.ic q_19_36=0
.ic qb_19_36=1.8
.ic q_20_36=0
.ic qb_20_36=1.8
.ic q_21_36=0
.ic qb_21_36=1.8
.ic q_22_36=0
.ic qb_22_36=1.8
.ic q_23_36=0
.ic qb_23_36=1.8
.ic q_24_36=0
.ic qb_24_36=1.8
.ic q_25_36=0
.ic qb_25_36=1.8
.ic q_26_36=0
.ic qb_26_36=1.8
.ic q_27_36=0
.ic qb_27_36=1.8
.ic q_28_36=0
.ic qb_28_36=1.8
.ic q_29_36=0
.ic qb_29_36=1.8
.ic q_30_36=0
.ic qb_30_36=1.8
.ic q_31_36=0
.ic qb_31_36=1.8
.ic q_32_36=0
.ic qb_32_36=1.8
.ic q_33_36=0
.ic qb_33_36=1.8
.ic q_34_36=0
.ic qb_34_36=1.8
.ic q_35_36=0
.ic qb_35_36=1.8
.ic q_36_36=0
.ic qb_36_36=1.8
.ic q_37_36=0
.ic qb_37_36=1.8
.ic q_38_36=0
.ic qb_38_36=1.8
.ic q_39_36=0
.ic qb_39_36=1.8
.ic q_40_36=0
.ic qb_40_36=1.8
.ic q_41_36=0
.ic qb_41_36=1.8
.ic q_42_36=0
.ic qb_42_36=1.8
.ic q_43_36=0
.ic qb_43_36=1.8
.ic q_44_36=0
.ic qb_44_36=1.8
.ic q_45_36=0
.ic qb_45_36=1.8
.ic q_46_36=0
.ic qb_46_36=1.8
.ic q_47_36=0
.ic qb_47_36=1.8
.ic q_48_36=0
.ic qb_48_36=1.8
.ic q_49_36=0
.ic qb_49_36=1.8
.ic q_50_36=0
.ic qb_50_36=1.8
.ic q_51_36=0
.ic qb_51_36=1.8
.ic q_52_36=0
.ic qb_52_36=1.8
.ic q_53_36=0
.ic qb_53_36=1.8
.ic q_54_36=0
.ic qb_54_36=1.8
.ic q_55_36=0
.ic qb_55_36=1.8
.ic q_56_36=0
.ic qb_56_36=1.8
.ic q_57_36=0
.ic qb_57_36=1.8
.ic q_58_36=0
.ic qb_58_36=1.8
.ic q_59_36=0
.ic qb_59_36=1.8
.ic q_60_36=0
.ic qb_60_36=1.8
.ic q_61_36=0
.ic qb_61_36=1.8
.ic q_62_36=0
.ic qb_62_36=1.8
.ic q_63_36=0
.ic qb_63_36=1.8
.ic q_64_36=0
.ic qb_64_36=1.8
.ic q_65_36=0
.ic qb_65_36=1.8
.ic q_66_36=0
.ic qb_66_36=1.8
.ic q_67_36=0
.ic qb_67_36=1.8
.ic q_68_36=0
.ic qb_68_36=1.8
.ic q_69_36=0
.ic qb_69_36=1.8
.ic q_70_36=0
.ic qb_70_36=1.8
.ic q_71_36=0
.ic qb_71_36=1.8
.ic q_72_36=0
.ic qb_72_36=1.8
.ic q_73_36=0
.ic qb_73_36=1.8
.ic q_74_36=0
.ic qb_74_36=1.8
.ic q_75_36=0
.ic qb_75_36=1.8
.ic q_76_36=0
.ic qb_76_36=1.8
.ic q_77_36=0
.ic qb_77_36=1.8
.ic q_78_36=0
.ic qb_78_36=1.8
.ic q_79_36=0
.ic qb_79_36=1.8
.ic q_80_36=0
.ic qb_80_36=1.8
.ic q_81_36=0
.ic qb_81_36=1.8
.ic q_82_36=0
.ic qb_82_36=1.8
.ic q_83_36=0
.ic qb_83_36=1.8
.ic q_84_36=0
.ic qb_84_36=1.8
.ic q_85_36=0
.ic qb_85_36=1.8
.ic q_86_36=0
.ic qb_86_36=1.8
.ic q_87_36=0
.ic qb_87_36=1.8
.ic q_88_36=0
.ic qb_88_36=1.8
.ic q_89_36=0
.ic qb_89_36=1.8
.ic q_90_36=0
.ic qb_90_36=1.8
.ic q_91_36=0
.ic qb_91_36=1.8
.ic q_92_36=0
.ic qb_92_36=1.8
.ic q_93_36=0
.ic qb_93_36=1.8
.ic q_94_36=0
.ic qb_94_36=1.8
.ic q_95_36=0
.ic qb_95_36=1.8
.ic q_96_36=0
.ic qb_96_36=1.8
.ic q_97_36=0
.ic qb_97_36=1.8
.ic q_98_36=0
.ic qb_98_36=1.8
.ic q_99_36=0
.ic qb_99_36=1.8
.ic q_0_37=0
.ic qb_0_37=1.8
.ic q_1_37=0
.ic qb_1_37=1.8
.ic q_2_37=0
.ic qb_2_37=1.8
.ic q_3_37=0
.ic qb_3_37=1.8
.ic q_4_37=0
.ic qb_4_37=1.8
.ic q_5_37=0
.ic qb_5_37=1.8
.ic q_6_37=0
.ic qb_6_37=1.8
.ic q_7_37=0
.ic qb_7_37=1.8
.ic q_8_37=0
.ic qb_8_37=1.8
.ic q_9_37=0
.ic qb_9_37=1.8
.ic q_10_37=0
.ic qb_10_37=1.8
.ic q_11_37=0
.ic qb_11_37=1.8
.ic q_12_37=0
.ic qb_12_37=1.8
.ic q_13_37=0
.ic qb_13_37=1.8
.ic q_14_37=0
.ic qb_14_37=1.8
.ic q_15_37=0
.ic qb_15_37=1.8
.ic q_16_37=0
.ic qb_16_37=1.8
.ic q_17_37=0
.ic qb_17_37=1.8
.ic q_18_37=0
.ic qb_18_37=1.8
.ic q_19_37=0
.ic qb_19_37=1.8
.ic q_20_37=0
.ic qb_20_37=1.8
.ic q_21_37=0
.ic qb_21_37=1.8
.ic q_22_37=0
.ic qb_22_37=1.8
.ic q_23_37=0
.ic qb_23_37=1.8
.ic q_24_37=0
.ic qb_24_37=1.8
.ic q_25_37=0
.ic qb_25_37=1.8
.ic q_26_37=0
.ic qb_26_37=1.8
.ic q_27_37=0
.ic qb_27_37=1.8
.ic q_28_37=0
.ic qb_28_37=1.8
.ic q_29_37=0
.ic qb_29_37=1.8
.ic q_30_37=0
.ic qb_30_37=1.8
.ic q_31_37=0
.ic qb_31_37=1.8
.ic q_32_37=0
.ic qb_32_37=1.8
.ic q_33_37=0
.ic qb_33_37=1.8
.ic q_34_37=0
.ic qb_34_37=1.8
.ic q_35_37=0
.ic qb_35_37=1.8
.ic q_36_37=0
.ic qb_36_37=1.8
.ic q_37_37=0
.ic qb_37_37=1.8
.ic q_38_37=0
.ic qb_38_37=1.8
.ic q_39_37=0
.ic qb_39_37=1.8
.ic q_40_37=0
.ic qb_40_37=1.8
.ic q_41_37=0
.ic qb_41_37=1.8
.ic q_42_37=0
.ic qb_42_37=1.8
.ic q_43_37=0
.ic qb_43_37=1.8
.ic q_44_37=0
.ic qb_44_37=1.8
.ic q_45_37=0
.ic qb_45_37=1.8
.ic q_46_37=0
.ic qb_46_37=1.8
.ic q_47_37=0
.ic qb_47_37=1.8
.ic q_48_37=0
.ic qb_48_37=1.8
.ic q_49_37=0
.ic qb_49_37=1.8
.ic q_50_37=0
.ic qb_50_37=1.8
.ic q_51_37=0
.ic qb_51_37=1.8
.ic q_52_37=0
.ic qb_52_37=1.8
.ic q_53_37=0
.ic qb_53_37=1.8
.ic q_54_37=0
.ic qb_54_37=1.8
.ic q_55_37=0
.ic qb_55_37=1.8
.ic q_56_37=0
.ic qb_56_37=1.8
.ic q_57_37=0
.ic qb_57_37=1.8
.ic q_58_37=0
.ic qb_58_37=1.8
.ic q_59_37=0
.ic qb_59_37=1.8
.ic q_60_37=0
.ic qb_60_37=1.8
.ic q_61_37=0
.ic qb_61_37=1.8
.ic q_62_37=0
.ic qb_62_37=1.8
.ic q_63_37=0
.ic qb_63_37=1.8
.ic q_64_37=0
.ic qb_64_37=1.8
.ic q_65_37=0
.ic qb_65_37=1.8
.ic q_66_37=0
.ic qb_66_37=1.8
.ic q_67_37=0
.ic qb_67_37=1.8
.ic q_68_37=0
.ic qb_68_37=1.8
.ic q_69_37=0
.ic qb_69_37=1.8
.ic q_70_37=0
.ic qb_70_37=1.8
.ic q_71_37=0
.ic qb_71_37=1.8
.ic q_72_37=0
.ic qb_72_37=1.8
.ic q_73_37=0
.ic qb_73_37=1.8
.ic q_74_37=0
.ic qb_74_37=1.8
.ic q_75_37=0
.ic qb_75_37=1.8
.ic q_76_37=0
.ic qb_76_37=1.8
.ic q_77_37=0
.ic qb_77_37=1.8
.ic q_78_37=0
.ic qb_78_37=1.8
.ic q_79_37=0
.ic qb_79_37=1.8
.ic q_80_37=0
.ic qb_80_37=1.8
.ic q_81_37=0
.ic qb_81_37=1.8
.ic q_82_37=0
.ic qb_82_37=1.8
.ic q_83_37=0
.ic qb_83_37=1.8
.ic q_84_37=0
.ic qb_84_37=1.8
.ic q_85_37=0
.ic qb_85_37=1.8
.ic q_86_37=0
.ic qb_86_37=1.8
.ic q_87_37=0
.ic qb_87_37=1.8
.ic q_88_37=0
.ic qb_88_37=1.8
.ic q_89_37=0
.ic qb_89_37=1.8
.ic q_90_37=0
.ic qb_90_37=1.8
.ic q_91_37=0
.ic qb_91_37=1.8
.ic q_92_37=0
.ic qb_92_37=1.8
.ic q_93_37=0
.ic qb_93_37=1.8
.ic q_94_37=0
.ic qb_94_37=1.8
.ic q_95_37=0
.ic qb_95_37=1.8
.ic q_96_37=0
.ic qb_96_37=1.8
.ic q_97_37=0
.ic qb_97_37=1.8
.ic q_98_37=0
.ic qb_98_37=1.8
.ic q_99_37=0
.ic qb_99_37=1.8
.ic q_0_38=0
.ic qb_0_38=1.8
.ic q_1_38=0
.ic qb_1_38=1.8
.ic q_2_38=0
.ic qb_2_38=1.8
.ic q_3_38=0
.ic qb_3_38=1.8
.ic q_4_38=0
.ic qb_4_38=1.8
.ic q_5_38=0
.ic qb_5_38=1.8
.ic q_6_38=0
.ic qb_6_38=1.8
.ic q_7_38=0
.ic qb_7_38=1.8
.ic q_8_38=0
.ic qb_8_38=1.8
.ic q_9_38=0
.ic qb_9_38=1.8
.ic q_10_38=0
.ic qb_10_38=1.8
.ic q_11_38=0
.ic qb_11_38=1.8
.ic q_12_38=0
.ic qb_12_38=1.8
.ic q_13_38=0
.ic qb_13_38=1.8
.ic q_14_38=0
.ic qb_14_38=1.8
.ic q_15_38=0
.ic qb_15_38=1.8
.ic q_16_38=0
.ic qb_16_38=1.8
.ic q_17_38=0
.ic qb_17_38=1.8
.ic q_18_38=0
.ic qb_18_38=1.8
.ic q_19_38=0
.ic qb_19_38=1.8
.ic q_20_38=0
.ic qb_20_38=1.8
.ic q_21_38=0
.ic qb_21_38=1.8
.ic q_22_38=0
.ic qb_22_38=1.8
.ic q_23_38=0
.ic qb_23_38=1.8
.ic q_24_38=0
.ic qb_24_38=1.8
.ic q_25_38=0
.ic qb_25_38=1.8
.ic q_26_38=0
.ic qb_26_38=1.8
.ic q_27_38=0
.ic qb_27_38=1.8
.ic q_28_38=0
.ic qb_28_38=1.8
.ic q_29_38=0
.ic qb_29_38=1.8
.ic q_30_38=0
.ic qb_30_38=1.8
.ic q_31_38=0
.ic qb_31_38=1.8
.ic q_32_38=0
.ic qb_32_38=1.8
.ic q_33_38=0
.ic qb_33_38=1.8
.ic q_34_38=0
.ic qb_34_38=1.8
.ic q_35_38=0
.ic qb_35_38=1.8
.ic q_36_38=0
.ic qb_36_38=1.8
.ic q_37_38=0
.ic qb_37_38=1.8
.ic q_38_38=0
.ic qb_38_38=1.8
.ic q_39_38=0
.ic qb_39_38=1.8
.ic q_40_38=0
.ic qb_40_38=1.8
.ic q_41_38=0
.ic qb_41_38=1.8
.ic q_42_38=0
.ic qb_42_38=1.8
.ic q_43_38=0
.ic qb_43_38=1.8
.ic q_44_38=0
.ic qb_44_38=1.8
.ic q_45_38=0
.ic qb_45_38=1.8
.ic q_46_38=0
.ic qb_46_38=1.8
.ic q_47_38=0
.ic qb_47_38=1.8
.ic q_48_38=0
.ic qb_48_38=1.8
.ic q_49_38=0
.ic qb_49_38=1.8
.ic q_50_38=0
.ic qb_50_38=1.8
.ic q_51_38=0
.ic qb_51_38=1.8
.ic q_52_38=0
.ic qb_52_38=1.8
.ic q_53_38=0
.ic qb_53_38=1.8
.ic q_54_38=0
.ic qb_54_38=1.8
.ic q_55_38=0
.ic qb_55_38=1.8
.ic q_56_38=0
.ic qb_56_38=1.8
.ic q_57_38=0
.ic qb_57_38=1.8
.ic q_58_38=0
.ic qb_58_38=1.8
.ic q_59_38=0
.ic qb_59_38=1.8
.ic q_60_38=0
.ic qb_60_38=1.8
.ic q_61_38=0
.ic qb_61_38=1.8
.ic q_62_38=0
.ic qb_62_38=1.8
.ic q_63_38=0
.ic qb_63_38=1.8
.ic q_64_38=0
.ic qb_64_38=1.8
.ic q_65_38=0
.ic qb_65_38=1.8
.ic q_66_38=0
.ic qb_66_38=1.8
.ic q_67_38=0
.ic qb_67_38=1.8
.ic q_68_38=0
.ic qb_68_38=1.8
.ic q_69_38=0
.ic qb_69_38=1.8
.ic q_70_38=0
.ic qb_70_38=1.8
.ic q_71_38=0
.ic qb_71_38=1.8
.ic q_72_38=0
.ic qb_72_38=1.8
.ic q_73_38=0
.ic qb_73_38=1.8
.ic q_74_38=0
.ic qb_74_38=1.8
.ic q_75_38=0
.ic qb_75_38=1.8
.ic q_76_38=0
.ic qb_76_38=1.8
.ic q_77_38=0
.ic qb_77_38=1.8
.ic q_78_38=0
.ic qb_78_38=1.8
.ic q_79_38=0
.ic qb_79_38=1.8
.ic q_80_38=0
.ic qb_80_38=1.8
.ic q_81_38=0
.ic qb_81_38=1.8
.ic q_82_38=0
.ic qb_82_38=1.8
.ic q_83_38=0
.ic qb_83_38=1.8
.ic q_84_38=0
.ic qb_84_38=1.8
.ic q_85_38=0
.ic qb_85_38=1.8
.ic q_86_38=0
.ic qb_86_38=1.8
.ic q_87_38=0
.ic qb_87_38=1.8
.ic q_88_38=0
.ic qb_88_38=1.8
.ic q_89_38=0
.ic qb_89_38=1.8
.ic q_90_38=0
.ic qb_90_38=1.8
.ic q_91_38=0
.ic qb_91_38=1.8
.ic q_92_38=0
.ic qb_92_38=1.8
.ic q_93_38=0
.ic qb_93_38=1.8
.ic q_94_38=0
.ic qb_94_38=1.8
.ic q_95_38=0
.ic qb_95_38=1.8
.ic q_96_38=0
.ic qb_96_38=1.8
.ic q_97_38=0
.ic qb_97_38=1.8
.ic q_98_38=0
.ic qb_98_38=1.8
.ic q_99_38=0
.ic qb_99_38=1.8
.ic q_0_39=0
.ic qb_0_39=1.8
.ic q_1_39=0
.ic qb_1_39=1.8
.ic q_2_39=0
.ic qb_2_39=1.8
.ic q_3_39=0
.ic qb_3_39=1.8
.ic q_4_39=0
.ic qb_4_39=1.8
.ic q_5_39=0
.ic qb_5_39=1.8
.ic q_6_39=0
.ic qb_6_39=1.8
.ic q_7_39=0
.ic qb_7_39=1.8
.ic q_8_39=0
.ic qb_8_39=1.8
.ic q_9_39=0
.ic qb_9_39=1.8
.ic q_10_39=0
.ic qb_10_39=1.8
.ic q_11_39=0
.ic qb_11_39=1.8
.ic q_12_39=0
.ic qb_12_39=1.8
.ic q_13_39=0
.ic qb_13_39=1.8
.ic q_14_39=0
.ic qb_14_39=1.8
.ic q_15_39=0
.ic qb_15_39=1.8
.ic q_16_39=0
.ic qb_16_39=1.8
.ic q_17_39=0
.ic qb_17_39=1.8
.ic q_18_39=0
.ic qb_18_39=1.8
.ic q_19_39=0
.ic qb_19_39=1.8
.ic q_20_39=0
.ic qb_20_39=1.8
.ic q_21_39=0
.ic qb_21_39=1.8
.ic q_22_39=0
.ic qb_22_39=1.8
.ic q_23_39=0
.ic qb_23_39=1.8
.ic q_24_39=0
.ic qb_24_39=1.8
.ic q_25_39=0
.ic qb_25_39=1.8
.ic q_26_39=0
.ic qb_26_39=1.8
.ic q_27_39=0
.ic qb_27_39=1.8
.ic q_28_39=0
.ic qb_28_39=1.8
.ic q_29_39=0
.ic qb_29_39=1.8
.ic q_30_39=0
.ic qb_30_39=1.8
.ic q_31_39=0
.ic qb_31_39=1.8
.ic q_32_39=0
.ic qb_32_39=1.8
.ic q_33_39=0
.ic qb_33_39=1.8
.ic q_34_39=0
.ic qb_34_39=1.8
.ic q_35_39=0
.ic qb_35_39=1.8
.ic q_36_39=0
.ic qb_36_39=1.8
.ic q_37_39=0
.ic qb_37_39=1.8
.ic q_38_39=0
.ic qb_38_39=1.8
.ic q_39_39=0
.ic qb_39_39=1.8
.ic q_40_39=0
.ic qb_40_39=1.8
.ic q_41_39=0
.ic qb_41_39=1.8
.ic q_42_39=0
.ic qb_42_39=1.8
.ic q_43_39=0
.ic qb_43_39=1.8
.ic q_44_39=0
.ic qb_44_39=1.8
.ic q_45_39=0
.ic qb_45_39=1.8
.ic q_46_39=0
.ic qb_46_39=1.8
.ic q_47_39=0
.ic qb_47_39=1.8
.ic q_48_39=0
.ic qb_48_39=1.8
.ic q_49_39=0
.ic qb_49_39=1.8
.ic q_50_39=0
.ic qb_50_39=1.8
.ic q_51_39=0
.ic qb_51_39=1.8
.ic q_52_39=0
.ic qb_52_39=1.8
.ic q_53_39=0
.ic qb_53_39=1.8
.ic q_54_39=0
.ic qb_54_39=1.8
.ic q_55_39=0
.ic qb_55_39=1.8
.ic q_56_39=0
.ic qb_56_39=1.8
.ic q_57_39=0
.ic qb_57_39=1.8
.ic q_58_39=0
.ic qb_58_39=1.8
.ic q_59_39=0
.ic qb_59_39=1.8
.ic q_60_39=0
.ic qb_60_39=1.8
.ic q_61_39=0
.ic qb_61_39=1.8
.ic q_62_39=0
.ic qb_62_39=1.8
.ic q_63_39=0
.ic qb_63_39=1.8
.ic q_64_39=0
.ic qb_64_39=1.8
.ic q_65_39=0
.ic qb_65_39=1.8
.ic q_66_39=0
.ic qb_66_39=1.8
.ic q_67_39=0
.ic qb_67_39=1.8
.ic q_68_39=0
.ic qb_68_39=1.8
.ic q_69_39=0
.ic qb_69_39=1.8
.ic q_70_39=0
.ic qb_70_39=1.8
.ic q_71_39=0
.ic qb_71_39=1.8
.ic q_72_39=0
.ic qb_72_39=1.8
.ic q_73_39=0
.ic qb_73_39=1.8
.ic q_74_39=0
.ic qb_74_39=1.8
.ic q_75_39=0
.ic qb_75_39=1.8
.ic q_76_39=0
.ic qb_76_39=1.8
.ic q_77_39=0
.ic qb_77_39=1.8
.ic q_78_39=0
.ic qb_78_39=1.8
.ic q_79_39=0
.ic qb_79_39=1.8
.ic q_80_39=0
.ic qb_80_39=1.8
.ic q_81_39=0
.ic qb_81_39=1.8
.ic q_82_39=0
.ic qb_82_39=1.8
.ic q_83_39=0
.ic qb_83_39=1.8
.ic q_84_39=0
.ic qb_84_39=1.8
.ic q_85_39=0
.ic qb_85_39=1.8
.ic q_86_39=0
.ic qb_86_39=1.8
.ic q_87_39=0
.ic qb_87_39=1.8
.ic q_88_39=0
.ic qb_88_39=1.8
.ic q_89_39=0
.ic qb_89_39=1.8
.ic q_90_39=0
.ic qb_90_39=1.8
.ic q_91_39=0
.ic qb_91_39=1.8
.ic q_92_39=0
.ic qb_92_39=1.8
.ic q_93_39=0
.ic qb_93_39=1.8
.ic q_94_39=0
.ic qb_94_39=1.8
.ic q_95_39=0
.ic qb_95_39=1.8
.ic q_96_39=0
.ic qb_96_39=1.8
.ic q_97_39=0
.ic qb_97_39=1.8
.ic q_98_39=0
.ic qb_98_39=1.8
.ic q_99_39=0
.ic qb_99_39=1.8
.ic q_0_40=0
.ic qb_0_40=1.8
.ic q_1_40=0
.ic qb_1_40=1.8
.ic q_2_40=0
.ic qb_2_40=1.8
.ic q_3_40=0
.ic qb_3_40=1.8
.ic q_4_40=0
.ic qb_4_40=1.8
.ic q_5_40=0
.ic qb_5_40=1.8
.ic q_6_40=0
.ic qb_6_40=1.8
.ic q_7_40=0
.ic qb_7_40=1.8
.ic q_8_40=0
.ic qb_8_40=1.8
.ic q_9_40=0
.ic qb_9_40=1.8
.ic q_10_40=0
.ic qb_10_40=1.8
.ic q_11_40=0
.ic qb_11_40=1.8
.ic q_12_40=0
.ic qb_12_40=1.8
.ic q_13_40=0
.ic qb_13_40=1.8
.ic q_14_40=0
.ic qb_14_40=1.8
.ic q_15_40=0
.ic qb_15_40=1.8
.ic q_16_40=0
.ic qb_16_40=1.8
.ic q_17_40=0
.ic qb_17_40=1.8
.ic q_18_40=0
.ic qb_18_40=1.8
.ic q_19_40=0
.ic qb_19_40=1.8
.ic q_20_40=0
.ic qb_20_40=1.8
.ic q_21_40=0
.ic qb_21_40=1.8
.ic q_22_40=0
.ic qb_22_40=1.8
.ic q_23_40=0
.ic qb_23_40=1.8
.ic q_24_40=0
.ic qb_24_40=1.8
.ic q_25_40=0
.ic qb_25_40=1.8
.ic q_26_40=0
.ic qb_26_40=1.8
.ic q_27_40=0
.ic qb_27_40=1.8
.ic q_28_40=0
.ic qb_28_40=1.8
.ic q_29_40=0
.ic qb_29_40=1.8
.ic q_30_40=0
.ic qb_30_40=1.8
.ic q_31_40=0
.ic qb_31_40=1.8
.ic q_32_40=0
.ic qb_32_40=1.8
.ic q_33_40=0
.ic qb_33_40=1.8
.ic q_34_40=0
.ic qb_34_40=1.8
.ic q_35_40=0
.ic qb_35_40=1.8
.ic q_36_40=0
.ic qb_36_40=1.8
.ic q_37_40=0
.ic qb_37_40=1.8
.ic q_38_40=0
.ic qb_38_40=1.8
.ic q_39_40=0
.ic qb_39_40=1.8
.ic q_40_40=0
.ic qb_40_40=1.8
.ic q_41_40=0
.ic qb_41_40=1.8
.ic q_42_40=0
.ic qb_42_40=1.8
.ic q_43_40=0
.ic qb_43_40=1.8
.ic q_44_40=0
.ic qb_44_40=1.8
.ic q_45_40=0
.ic qb_45_40=1.8
.ic q_46_40=0
.ic qb_46_40=1.8
.ic q_47_40=0
.ic qb_47_40=1.8
.ic q_48_40=0
.ic qb_48_40=1.8
.ic q_49_40=0
.ic qb_49_40=1.8
.ic q_50_40=0
.ic qb_50_40=1.8
.ic q_51_40=0
.ic qb_51_40=1.8
.ic q_52_40=0
.ic qb_52_40=1.8
.ic q_53_40=0
.ic qb_53_40=1.8
.ic q_54_40=0
.ic qb_54_40=1.8
.ic q_55_40=0
.ic qb_55_40=1.8
.ic q_56_40=0
.ic qb_56_40=1.8
.ic q_57_40=0
.ic qb_57_40=1.8
.ic q_58_40=0
.ic qb_58_40=1.8
.ic q_59_40=0
.ic qb_59_40=1.8
.ic q_60_40=0
.ic qb_60_40=1.8
.ic q_61_40=0
.ic qb_61_40=1.8
.ic q_62_40=0
.ic qb_62_40=1.8
.ic q_63_40=0
.ic qb_63_40=1.8
.ic q_64_40=0
.ic qb_64_40=1.8
.ic q_65_40=0
.ic qb_65_40=1.8
.ic q_66_40=0
.ic qb_66_40=1.8
.ic q_67_40=0
.ic qb_67_40=1.8
.ic q_68_40=0
.ic qb_68_40=1.8
.ic q_69_40=0
.ic qb_69_40=1.8
.ic q_70_40=0
.ic qb_70_40=1.8
.ic q_71_40=0
.ic qb_71_40=1.8
.ic q_72_40=0
.ic qb_72_40=1.8
.ic q_73_40=0
.ic qb_73_40=1.8
.ic q_74_40=0
.ic qb_74_40=1.8
.ic q_75_40=0
.ic qb_75_40=1.8
.ic q_76_40=0
.ic qb_76_40=1.8
.ic q_77_40=0
.ic qb_77_40=1.8
.ic q_78_40=0
.ic qb_78_40=1.8
.ic q_79_40=0
.ic qb_79_40=1.8
.ic q_80_40=0
.ic qb_80_40=1.8
.ic q_81_40=0
.ic qb_81_40=1.8
.ic q_82_40=0
.ic qb_82_40=1.8
.ic q_83_40=0
.ic qb_83_40=1.8
.ic q_84_40=0
.ic qb_84_40=1.8
.ic q_85_40=0
.ic qb_85_40=1.8
.ic q_86_40=0
.ic qb_86_40=1.8
.ic q_87_40=0
.ic qb_87_40=1.8
.ic q_88_40=0
.ic qb_88_40=1.8
.ic q_89_40=0
.ic qb_89_40=1.8
.ic q_90_40=0
.ic qb_90_40=1.8
.ic q_91_40=0
.ic qb_91_40=1.8
.ic q_92_40=0
.ic qb_92_40=1.8
.ic q_93_40=0
.ic qb_93_40=1.8
.ic q_94_40=0
.ic qb_94_40=1.8
.ic q_95_40=0
.ic qb_95_40=1.8
.ic q_96_40=0
.ic qb_96_40=1.8
.ic q_97_40=0
.ic qb_97_40=1.8
.ic q_98_40=0
.ic qb_98_40=1.8
.ic q_99_40=0
.ic qb_99_40=1.8
.ic q_0_41=0
.ic qb_0_41=1.8
.ic q_1_41=0
.ic qb_1_41=1.8
.ic q_2_41=0
.ic qb_2_41=1.8
.ic q_3_41=0
.ic qb_3_41=1.8
.ic q_4_41=0
.ic qb_4_41=1.8
.ic q_5_41=0
.ic qb_5_41=1.8
.ic q_6_41=0
.ic qb_6_41=1.8
.ic q_7_41=0
.ic qb_7_41=1.8
.ic q_8_41=0
.ic qb_8_41=1.8
.ic q_9_41=0
.ic qb_9_41=1.8
.ic q_10_41=0
.ic qb_10_41=1.8
.ic q_11_41=0
.ic qb_11_41=1.8
.ic q_12_41=0
.ic qb_12_41=1.8
.ic q_13_41=0
.ic qb_13_41=1.8
.ic q_14_41=0
.ic qb_14_41=1.8
.ic q_15_41=0
.ic qb_15_41=1.8
.ic q_16_41=0
.ic qb_16_41=1.8
.ic q_17_41=0
.ic qb_17_41=1.8
.ic q_18_41=0
.ic qb_18_41=1.8
.ic q_19_41=0
.ic qb_19_41=1.8
.ic q_20_41=0
.ic qb_20_41=1.8
.ic q_21_41=0
.ic qb_21_41=1.8
.ic q_22_41=0
.ic qb_22_41=1.8
.ic q_23_41=0
.ic qb_23_41=1.8
.ic q_24_41=0
.ic qb_24_41=1.8
.ic q_25_41=0
.ic qb_25_41=1.8
.ic q_26_41=0
.ic qb_26_41=1.8
.ic q_27_41=0
.ic qb_27_41=1.8
.ic q_28_41=0
.ic qb_28_41=1.8
.ic q_29_41=0
.ic qb_29_41=1.8
.ic q_30_41=0
.ic qb_30_41=1.8
.ic q_31_41=0
.ic qb_31_41=1.8
.ic q_32_41=0
.ic qb_32_41=1.8
.ic q_33_41=0
.ic qb_33_41=1.8
.ic q_34_41=0
.ic qb_34_41=1.8
.ic q_35_41=0
.ic qb_35_41=1.8
.ic q_36_41=0
.ic qb_36_41=1.8
.ic q_37_41=0
.ic qb_37_41=1.8
.ic q_38_41=0
.ic qb_38_41=1.8
.ic q_39_41=0
.ic qb_39_41=1.8
.ic q_40_41=0
.ic qb_40_41=1.8
.ic q_41_41=0
.ic qb_41_41=1.8
.ic q_42_41=0
.ic qb_42_41=1.8
.ic q_43_41=0
.ic qb_43_41=1.8
.ic q_44_41=0
.ic qb_44_41=1.8
.ic q_45_41=0
.ic qb_45_41=1.8
.ic q_46_41=0
.ic qb_46_41=1.8
.ic q_47_41=0
.ic qb_47_41=1.8
.ic q_48_41=0
.ic qb_48_41=1.8
.ic q_49_41=0
.ic qb_49_41=1.8
.ic q_50_41=0
.ic qb_50_41=1.8
.ic q_51_41=0
.ic qb_51_41=1.8
.ic q_52_41=0
.ic qb_52_41=1.8
.ic q_53_41=0
.ic qb_53_41=1.8
.ic q_54_41=0
.ic qb_54_41=1.8
.ic q_55_41=0
.ic qb_55_41=1.8
.ic q_56_41=0
.ic qb_56_41=1.8
.ic q_57_41=0
.ic qb_57_41=1.8
.ic q_58_41=0
.ic qb_58_41=1.8
.ic q_59_41=0
.ic qb_59_41=1.8
.ic q_60_41=0
.ic qb_60_41=1.8
.ic q_61_41=0
.ic qb_61_41=1.8
.ic q_62_41=0
.ic qb_62_41=1.8
.ic q_63_41=0
.ic qb_63_41=1.8
.ic q_64_41=0
.ic qb_64_41=1.8
.ic q_65_41=0
.ic qb_65_41=1.8
.ic q_66_41=0
.ic qb_66_41=1.8
.ic q_67_41=0
.ic qb_67_41=1.8
.ic q_68_41=0
.ic qb_68_41=1.8
.ic q_69_41=0
.ic qb_69_41=1.8
.ic q_70_41=0
.ic qb_70_41=1.8
.ic q_71_41=0
.ic qb_71_41=1.8
.ic q_72_41=0
.ic qb_72_41=1.8
.ic q_73_41=0
.ic qb_73_41=1.8
.ic q_74_41=0
.ic qb_74_41=1.8
.ic q_75_41=0
.ic qb_75_41=1.8
.ic q_76_41=0
.ic qb_76_41=1.8
.ic q_77_41=0
.ic qb_77_41=1.8
.ic q_78_41=0
.ic qb_78_41=1.8
.ic q_79_41=0
.ic qb_79_41=1.8
.ic q_80_41=0
.ic qb_80_41=1.8
.ic q_81_41=0
.ic qb_81_41=1.8
.ic q_82_41=0
.ic qb_82_41=1.8
.ic q_83_41=0
.ic qb_83_41=1.8
.ic q_84_41=0
.ic qb_84_41=1.8
.ic q_85_41=0
.ic qb_85_41=1.8
.ic q_86_41=0
.ic qb_86_41=1.8
.ic q_87_41=0
.ic qb_87_41=1.8
.ic q_88_41=0
.ic qb_88_41=1.8
.ic q_89_41=0
.ic qb_89_41=1.8
.ic q_90_41=0
.ic qb_90_41=1.8
.ic q_91_41=0
.ic qb_91_41=1.8
.ic q_92_41=0
.ic qb_92_41=1.8
.ic q_93_41=0
.ic qb_93_41=1.8
.ic q_94_41=0
.ic qb_94_41=1.8
.ic q_95_41=0
.ic qb_95_41=1.8
.ic q_96_41=0
.ic qb_96_41=1.8
.ic q_97_41=0
.ic qb_97_41=1.8
.ic q_98_41=0
.ic qb_98_41=1.8
.ic q_99_41=0
.ic qb_99_41=1.8
.ic q_0_42=0
.ic qb_0_42=1.8
.ic q_1_42=0
.ic qb_1_42=1.8
.ic q_2_42=0
.ic qb_2_42=1.8
.ic q_3_42=0
.ic qb_3_42=1.8
.ic q_4_42=0
.ic qb_4_42=1.8
.ic q_5_42=0
.ic qb_5_42=1.8
.ic q_6_42=0
.ic qb_6_42=1.8
.ic q_7_42=0
.ic qb_7_42=1.8
.ic q_8_42=0
.ic qb_8_42=1.8
.ic q_9_42=0
.ic qb_9_42=1.8
.ic q_10_42=0
.ic qb_10_42=1.8
.ic q_11_42=0
.ic qb_11_42=1.8
.ic q_12_42=0
.ic qb_12_42=1.8
.ic q_13_42=0
.ic qb_13_42=1.8
.ic q_14_42=0
.ic qb_14_42=1.8
.ic q_15_42=0
.ic qb_15_42=1.8
.ic q_16_42=0
.ic qb_16_42=1.8
.ic q_17_42=0
.ic qb_17_42=1.8
.ic q_18_42=0
.ic qb_18_42=1.8
.ic q_19_42=0
.ic qb_19_42=1.8
.ic q_20_42=0
.ic qb_20_42=1.8
.ic q_21_42=0
.ic qb_21_42=1.8
.ic q_22_42=0
.ic qb_22_42=1.8
.ic q_23_42=0
.ic qb_23_42=1.8
.ic q_24_42=0
.ic qb_24_42=1.8
.ic q_25_42=0
.ic qb_25_42=1.8
.ic q_26_42=0
.ic qb_26_42=1.8
.ic q_27_42=0
.ic qb_27_42=1.8
.ic q_28_42=0
.ic qb_28_42=1.8
.ic q_29_42=0
.ic qb_29_42=1.8
.ic q_30_42=0
.ic qb_30_42=1.8
.ic q_31_42=0
.ic qb_31_42=1.8
.ic q_32_42=0
.ic qb_32_42=1.8
.ic q_33_42=0
.ic qb_33_42=1.8
.ic q_34_42=0
.ic qb_34_42=1.8
.ic q_35_42=0
.ic qb_35_42=1.8
.ic q_36_42=0
.ic qb_36_42=1.8
.ic q_37_42=0
.ic qb_37_42=1.8
.ic q_38_42=0
.ic qb_38_42=1.8
.ic q_39_42=0
.ic qb_39_42=1.8
.ic q_40_42=0
.ic qb_40_42=1.8
.ic q_41_42=0
.ic qb_41_42=1.8
.ic q_42_42=0
.ic qb_42_42=1.8
.ic q_43_42=0
.ic qb_43_42=1.8
.ic q_44_42=0
.ic qb_44_42=1.8
.ic q_45_42=0
.ic qb_45_42=1.8
.ic q_46_42=0
.ic qb_46_42=1.8
.ic q_47_42=0
.ic qb_47_42=1.8
.ic q_48_42=0
.ic qb_48_42=1.8
.ic q_49_42=0
.ic qb_49_42=1.8
.ic q_50_42=0
.ic qb_50_42=1.8
.ic q_51_42=0
.ic qb_51_42=1.8
.ic q_52_42=0
.ic qb_52_42=1.8
.ic q_53_42=0
.ic qb_53_42=1.8
.ic q_54_42=0
.ic qb_54_42=1.8
.ic q_55_42=0
.ic qb_55_42=1.8
.ic q_56_42=0
.ic qb_56_42=1.8
.ic q_57_42=0
.ic qb_57_42=1.8
.ic q_58_42=0
.ic qb_58_42=1.8
.ic q_59_42=0
.ic qb_59_42=1.8
.ic q_60_42=0
.ic qb_60_42=1.8
.ic q_61_42=0
.ic qb_61_42=1.8
.ic q_62_42=0
.ic qb_62_42=1.8
.ic q_63_42=0
.ic qb_63_42=1.8
.ic q_64_42=0
.ic qb_64_42=1.8
.ic q_65_42=0
.ic qb_65_42=1.8
.ic q_66_42=0
.ic qb_66_42=1.8
.ic q_67_42=0
.ic qb_67_42=1.8
.ic q_68_42=0
.ic qb_68_42=1.8
.ic q_69_42=0
.ic qb_69_42=1.8
.ic q_70_42=0
.ic qb_70_42=1.8
.ic q_71_42=0
.ic qb_71_42=1.8
.ic q_72_42=0
.ic qb_72_42=1.8
.ic q_73_42=0
.ic qb_73_42=1.8
.ic q_74_42=0
.ic qb_74_42=1.8
.ic q_75_42=0
.ic qb_75_42=1.8
.ic q_76_42=0
.ic qb_76_42=1.8
.ic q_77_42=0
.ic qb_77_42=1.8
.ic q_78_42=0
.ic qb_78_42=1.8
.ic q_79_42=0
.ic qb_79_42=1.8
.ic q_80_42=0
.ic qb_80_42=1.8
.ic q_81_42=0
.ic qb_81_42=1.8
.ic q_82_42=0
.ic qb_82_42=1.8
.ic q_83_42=0
.ic qb_83_42=1.8
.ic q_84_42=0
.ic qb_84_42=1.8
.ic q_85_42=0
.ic qb_85_42=1.8
.ic q_86_42=0
.ic qb_86_42=1.8
.ic q_87_42=0
.ic qb_87_42=1.8
.ic q_88_42=0
.ic qb_88_42=1.8
.ic q_89_42=0
.ic qb_89_42=1.8
.ic q_90_42=0
.ic qb_90_42=1.8
.ic q_91_42=0
.ic qb_91_42=1.8
.ic q_92_42=0
.ic qb_92_42=1.8
.ic q_93_42=0
.ic qb_93_42=1.8
.ic q_94_42=0
.ic qb_94_42=1.8
.ic q_95_42=0
.ic qb_95_42=1.8
.ic q_96_42=0
.ic qb_96_42=1.8
.ic q_97_42=0
.ic qb_97_42=1.8
.ic q_98_42=0
.ic qb_98_42=1.8
.ic q_99_42=0
.ic qb_99_42=1.8
.ic q_0_43=0
.ic qb_0_43=1.8
.ic q_1_43=0
.ic qb_1_43=1.8
.ic q_2_43=0
.ic qb_2_43=1.8
.ic q_3_43=0
.ic qb_3_43=1.8
.ic q_4_43=0
.ic qb_4_43=1.8
.ic q_5_43=0
.ic qb_5_43=1.8
.ic q_6_43=0
.ic qb_6_43=1.8
.ic q_7_43=0
.ic qb_7_43=1.8
.ic q_8_43=0
.ic qb_8_43=1.8
.ic q_9_43=0
.ic qb_9_43=1.8
.ic q_10_43=0
.ic qb_10_43=1.8
.ic q_11_43=0
.ic qb_11_43=1.8
.ic q_12_43=0
.ic qb_12_43=1.8
.ic q_13_43=0
.ic qb_13_43=1.8
.ic q_14_43=0
.ic qb_14_43=1.8
.ic q_15_43=0
.ic qb_15_43=1.8
.ic q_16_43=0
.ic qb_16_43=1.8
.ic q_17_43=0
.ic qb_17_43=1.8
.ic q_18_43=0
.ic qb_18_43=1.8
.ic q_19_43=0
.ic qb_19_43=1.8
.ic q_20_43=0
.ic qb_20_43=1.8
.ic q_21_43=0
.ic qb_21_43=1.8
.ic q_22_43=0
.ic qb_22_43=1.8
.ic q_23_43=0
.ic qb_23_43=1.8
.ic q_24_43=0
.ic qb_24_43=1.8
.ic q_25_43=0
.ic qb_25_43=1.8
.ic q_26_43=0
.ic qb_26_43=1.8
.ic q_27_43=0
.ic qb_27_43=1.8
.ic q_28_43=0
.ic qb_28_43=1.8
.ic q_29_43=0
.ic qb_29_43=1.8
.ic q_30_43=0
.ic qb_30_43=1.8
.ic q_31_43=0
.ic qb_31_43=1.8
.ic q_32_43=0
.ic qb_32_43=1.8
.ic q_33_43=0
.ic qb_33_43=1.8
.ic q_34_43=0
.ic qb_34_43=1.8
.ic q_35_43=0
.ic qb_35_43=1.8
.ic q_36_43=0
.ic qb_36_43=1.8
.ic q_37_43=0
.ic qb_37_43=1.8
.ic q_38_43=0
.ic qb_38_43=1.8
.ic q_39_43=0
.ic qb_39_43=1.8
.ic q_40_43=0
.ic qb_40_43=1.8
.ic q_41_43=0
.ic qb_41_43=1.8
.ic q_42_43=0
.ic qb_42_43=1.8
.ic q_43_43=0
.ic qb_43_43=1.8
.ic q_44_43=0
.ic qb_44_43=1.8
.ic q_45_43=0
.ic qb_45_43=1.8
.ic q_46_43=0
.ic qb_46_43=1.8
.ic q_47_43=0
.ic qb_47_43=1.8
.ic q_48_43=0
.ic qb_48_43=1.8
.ic q_49_43=0
.ic qb_49_43=1.8
.ic q_50_43=0
.ic qb_50_43=1.8
.ic q_51_43=0
.ic qb_51_43=1.8
.ic q_52_43=0
.ic qb_52_43=1.8
.ic q_53_43=0
.ic qb_53_43=1.8
.ic q_54_43=0
.ic qb_54_43=1.8
.ic q_55_43=0
.ic qb_55_43=1.8
.ic q_56_43=0
.ic qb_56_43=1.8
.ic q_57_43=0
.ic qb_57_43=1.8
.ic q_58_43=0
.ic qb_58_43=1.8
.ic q_59_43=0
.ic qb_59_43=1.8
.ic q_60_43=0
.ic qb_60_43=1.8
.ic q_61_43=0
.ic qb_61_43=1.8
.ic q_62_43=0
.ic qb_62_43=1.8
.ic q_63_43=0
.ic qb_63_43=1.8
.ic q_64_43=0
.ic qb_64_43=1.8
.ic q_65_43=0
.ic qb_65_43=1.8
.ic q_66_43=0
.ic qb_66_43=1.8
.ic q_67_43=0
.ic qb_67_43=1.8
.ic q_68_43=0
.ic qb_68_43=1.8
.ic q_69_43=0
.ic qb_69_43=1.8
.ic q_70_43=0
.ic qb_70_43=1.8
.ic q_71_43=0
.ic qb_71_43=1.8
.ic q_72_43=0
.ic qb_72_43=1.8
.ic q_73_43=0
.ic qb_73_43=1.8
.ic q_74_43=0
.ic qb_74_43=1.8
.ic q_75_43=0
.ic qb_75_43=1.8
.ic q_76_43=0
.ic qb_76_43=1.8
.ic q_77_43=0
.ic qb_77_43=1.8
.ic q_78_43=0
.ic qb_78_43=1.8
.ic q_79_43=0
.ic qb_79_43=1.8
.ic q_80_43=0
.ic qb_80_43=1.8
.ic q_81_43=0
.ic qb_81_43=1.8
.ic q_82_43=0
.ic qb_82_43=1.8
.ic q_83_43=0
.ic qb_83_43=1.8
.ic q_84_43=0
.ic qb_84_43=1.8
.ic q_85_43=0
.ic qb_85_43=1.8
.ic q_86_43=0
.ic qb_86_43=1.8
.ic q_87_43=0
.ic qb_87_43=1.8
.ic q_88_43=0
.ic qb_88_43=1.8
.ic q_89_43=0
.ic qb_89_43=1.8
.ic q_90_43=0
.ic qb_90_43=1.8
.ic q_91_43=0
.ic qb_91_43=1.8
.ic q_92_43=0
.ic qb_92_43=1.8
.ic q_93_43=0
.ic qb_93_43=1.8
.ic q_94_43=0
.ic qb_94_43=1.8
.ic q_95_43=0
.ic qb_95_43=1.8
.ic q_96_43=0
.ic qb_96_43=1.8
.ic q_97_43=0
.ic qb_97_43=1.8
.ic q_98_43=0
.ic qb_98_43=1.8
.ic q_99_43=0
.ic qb_99_43=1.8
.ic q_0_44=0
.ic qb_0_44=1.8
.ic q_1_44=0
.ic qb_1_44=1.8
.ic q_2_44=0
.ic qb_2_44=1.8
.ic q_3_44=0
.ic qb_3_44=1.8
.ic q_4_44=0
.ic qb_4_44=1.8
.ic q_5_44=0
.ic qb_5_44=1.8
.ic q_6_44=0
.ic qb_6_44=1.8
.ic q_7_44=0
.ic qb_7_44=1.8
.ic q_8_44=0
.ic qb_8_44=1.8
.ic q_9_44=0
.ic qb_9_44=1.8
.ic q_10_44=0
.ic qb_10_44=1.8
.ic q_11_44=0
.ic qb_11_44=1.8
.ic q_12_44=0
.ic qb_12_44=1.8
.ic q_13_44=0
.ic qb_13_44=1.8
.ic q_14_44=0
.ic qb_14_44=1.8
.ic q_15_44=0
.ic qb_15_44=1.8
.ic q_16_44=0
.ic qb_16_44=1.8
.ic q_17_44=0
.ic qb_17_44=1.8
.ic q_18_44=0
.ic qb_18_44=1.8
.ic q_19_44=0
.ic qb_19_44=1.8
.ic q_20_44=0
.ic qb_20_44=1.8
.ic q_21_44=0
.ic qb_21_44=1.8
.ic q_22_44=0
.ic qb_22_44=1.8
.ic q_23_44=0
.ic qb_23_44=1.8
.ic q_24_44=0
.ic qb_24_44=1.8
.ic q_25_44=0
.ic qb_25_44=1.8
.ic q_26_44=0
.ic qb_26_44=1.8
.ic q_27_44=0
.ic qb_27_44=1.8
.ic q_28_44=0
.ic qb_28_44=1.8
.ic q_29_44=0
.ic qb_29_44=1.8
.ic q_30_44=0
.ic qb_30_44=1.8
.ic q_31_44=0
.ic qb_31_44=1.8
.ic q_32_44=0
.ic qb_32_44=1.8
.ic q_33_44=0
.ic qb_33_44=1.8
.ic q_34_44=0
.ic qb_34_44=1.8
.ic q_35_44=0
.ic qb_35_44=1.8
.ic q_36_44=0
.ic qb_36_44=1.8
.ic q_37_44=0
.ic qb_37_44=1.8
.ic q_38_44=0
.ic qb_38_44=1.8
.ic q_39_44=0
.ic qb_39_44=1.8
.ic q_40_44=0
.ic qb_40_44=1.8
.ic q_41_44=0
.ic qb_41_44=1.8
.ic q_42_44=0
.ic qb_42_44=1.8
.ic q_43_44=0
.ic qb_43_44=1.8
.ic q_44_44=0
.ic qb_44_44=1.8
.ic q_45_44=0
.ic qb_45_44=1.8
.ic q_46_44=0
.ic qb_46_44=1.8
.ic q_47_44=0
.ic qb_47_44=1.8
.ic q_48_44=0
.ic qb_48_44=1.8
.ic q_49_44=0
.ic qb_49_44=1.8
.ic q_50_44=0
.ic qb_50_44=1.8
.ic q_51_44=0
.ic qb_51_44=1.8
.ic q_52_44=0
.ic qb_52_44=1.8
.ic q_53_44=0
.ic qb_53_44=1.8
.ic q_54_44=0
.ic qb_54_44=1.8
.ic q_55_44=0
.ic qb_55_44=1.8
.ic q_56_44=0
.ic qb_56_44=1.8
.ic q_57_44=0
.ic qb_57_44=1.8
.ic q_58_44=0
.ic qb_58_44=1.8
.ic q_59_44=0
.ic qb_59_44=1.8
.ic q_60_44=0
.ic qb_60_44=1.8
.ic q_61_44=0
.ic qb_61_44=1.8
.ic q_62_44=0
.ic qb_62_44=1.8
.ic q_63_44=0
.ic qb_63_44=1.8
.ic q_64_44=0
.ic qb_64_44=1.8
.ic q_65_44=0
.ic qb_65_44=1.8
.ic q_66_44=0
.ic qb_66_44=1.8
.ic q_67_44=0
.ic qb_67_44=1.8
.ic q_68_44=0
.ic qb_68_44=1.8
.ic q_69_44=0
.ic qb_69_44=1.8
.ic q_70_44=0
.ic qb_70_44=1.8
.ic q_71_44=0
.ic qb_71_44=1.8
.ic q_72_44=0
.ic qb_72_44=1.8
.ic q_73_44=0
.ic qb_73_44=1.8
.ic q_74_44=0
.ic qb_74_44=1.8
.ic q_75_44=0
.ic qb_75_44=1.8
.ic q_76_44=0
.ic qb_76_44=1.8
.ic q_77_44=0
.ic qb_77_44=1.8
.ic q_78_44=0
.ic qb_78_44=1.8
.ic q_79_44=0
.ic qb_79_44=1.8
.ic q_80_44=0
.ic qb_80_44=1.8
.ic q_81_44=0
.ic qb_81_44=1.8
.ic q_82_44=0
.ic qb_82_44=1.8
.ic q_83_44=0
.ic qb_83_44=1.8
.ic q_84_44=0
.ic qb_84_44=1.8
.ic q_85_44=0
.ic qb_85_44=1.8
.ic q_86_44=0
.ic qb_86_44=1.8
.ic q_87_44=0
.ic qb_87_44=1.8
.ic q_88_44=0
.ic qb_88_44=1.8
.ic q_89_44=0
.ic qb_89_44=1.8
.ic q_90_44=0
.ic qb_90_44=1.8
.ic q_91_44=0
.ic qb_91_44=1.8
.ic q_92_44=0
.ic qb_92_44=1.8
.ic q_93_44=0
.ic qb_93_44=1.8
.ic q_94_44=0
.ic qb_94_44=1.8
.ic q_95_44=0
.ic qb_95_44=1.8
.ic q_96_44=0
.ic qb_96_44=1.8
.ic q_97_44=0
.ic qb_97_44=1.8
.ic q_98_44=0
.ic qb_98_44=1.8
.ic q_99_44=0
.ic qb_99_44=1.8
.ic q_0_45=0
.ic qb_0_45=1.8
.ic q_1_45=0
.ic qb_1_45=1.8
.ic q_2_45=0
.ic qb_2_45=1.8
.ic q_3_45=0
.ic qb_3_45=1.8
.ic q_4_45=0
.ic qb_4_45=1.8
.ic q_5_45=0
.ic qb_5_45=1.8
.ic q_6_45=0
.ic qb_6_45=1.8
.ic q_7_45=0
.ic qb_7_45=1.8
.ic q_8_45=0
.ic qb_8_45=1.8
.ic q_9_45=0
.ic qb_9_45=1.8
.ic q_10_45=0
.ic qb_10_45=1.8
.ic q_11_45=0
.ic qb_11_45=1.8
.ic q_12_45=0
.ic qb_12_45=1.8
.ic q_13_45=0
.ic qb_13_45=1.8
.ic q_14_45=0
.ic qb_14_45=1.8
.ic q_15_45=0
.ic qb_15_45=1.8
.ic q_16_45=0
.ic qb_16_45=1.8
.ic q_17_45=0
.ic qb_17_45=1.8
.ic q_18_45=0
.ic qb_18_45=1.8
.ic q_19_45=0
.ic qb_19_45=1.8
.ic q_20_45=0
.ic qb_20_45=1.8
.ic q_21_45=0
.ic qb_21_45=1.8
.ic q_22_45=0
.ic qb_22_45=1.8
.ic q_23_45=0
.ic qb_23_45=1.8
.ic q_24_45=0
.ic qb_24_45=1.8
.ic q_25_45=0
.ic qb_25_45=1.8
.ic q_26_45=0
.ic qb_26_45=1.8
.ic q_27_45=0
.ic qb_27_45=1.8
.ic q_28_45=0
.ic qb_28_45=1.8
.ic q_29_45=0
.ic qb_29_45=1.8
.ic q_30_45=0
.ic qb_30_45=1.8
.ic q_31_45=0
.ic qb_31_45=1.8
.ic q_32_45=0
.ic qb_32_45=1.8
.ic q_33_45=0
.ic qb_33_45=1.8
.ic q_34_45=0
.ic qb_34_45=1.8
.ic q_35_45=0
.ic qb_35_45=1.8
.ic q_36_45=0
.ic qb_36_45=1.8
.ic q_37_45=0
.ic qb_37_45=1.8
.ic q_38_45=0
.ic qb_38_45=1.8
.ic q_39_45=0
.ic qb_39_45=1.8
.ic q_40_45=0
.ic qb_40_45=1.8
.ic q_41_45=0
.ic qb_41_45=1.8
.ic q_42_45=0
.ic qb_42_45=1.8
.ic q_43_45=0
.ic qb_43_45=1.8
.ic q_44_45=0
.ic qb_44_45=1.8
.ic q_45_45=0
.ic qb_45_45=1.8
.ic q_46_45=0
.ic qb_46_45=1.8
.ic q_47_45=0
.ic qb_47_45=1.8
.ic q_48_45=0
.ic qb_48_45=1.8
.ic q_49_45=0
.ic qb_49_45=1.8
.ic q_50_45=0
.ic qb_50_45=1.8
.ic q_51_45=0
.ic qb_51_45=1.8
.ic q_52_45=0
.ic qb_52_45=1.8
.ic q_53_45=0
.ic qb_53_45=1.8
.ic q_54_45=0
.ic qb_54_45=1.8
.ic q_55_45=0
.ic qb_55_45=1.8
.ic q_56_45=0
.ic qb_56_45=1.8
.ic q_57_45=0
.ic qb_57_45=1.8
.ic q_58_45=0
.ic qb_58_45=1.8
.ic q_59_45=0
.ic qb_59_45=1.8
.ic q_60_45=0
.ic qb_60_45=1.8
.ic q_61_45=0
.ic qb_61_45=1.8
.ic q_62_45=0
.ic qb_62_45=1.8
.ic q_63_45=0
.ic qb_63_45=1.8
.ic q_64_45=0
.ic qb_64_45=1.8
.ic q_65_45=0
.ic qb_65_45=1.8
.ic q_66_45=0
.ic qb_66_45=1.8
.ic q_67_45=0
.ic qb_67_45=1.8
.ic q_68_45=0
.ic qb_68_45=1.8
.ic q_69_45=0
.ic qb_69_45=1.8
.ic q_70_45=0
.ic qb_70_45=1.8
.ic q_71_45=0
.ic qb_71_45=1.8
.ic q_72_45=0
.ic qb_72_45=1.8
.ic q_73_45=0
.ic qb_73_45=1.8
.ic q_74_45=0
.ic qb_74_45=1.8
.ic q_75_45=0
.ic qb_75_45=1.8
.ic q_76_45=0
.ic qb_76_45=1.8
.ic q_77_45=0
.ic qb_77_45=1.8
.ic q_78_45=0
.ic qb_78_45=1.8
.ic q_79_45=0
.ic qb_79_45=1.8
.ic q_80_45=0
.ic qb_80_45=1.8
.ic q_81_45=0
.ic qb_81_45=1.8
.ic q_82_45=0
.ic qb_82_45=1.8
.ic q_83_45=0
.ic qb_83_45=1.8
.ic q_84_45=0
.ic qb_84_45=1.8
.ic q_85_45=0
.ic qb_85_45=1.8
.ic q_86_45=0
.ic qb_86_45=1.8
.ic q_87_45=0
.ic qb_87_45=1.8
.ic q_88_45=0
.ic qb_88_45=1.8
.ic q_89_45=0
.ic qb_89_45=1.8
.ic q_90_45=0
.ic qb_90_45=1.8
.ic q_91_45=0
.ic qb_91_45=1.8
.ic q_92_45=0
.ic qb_92_45=1.8
.ic q_93_45=0
.ic qb_93_45=1.8
.ic q_94_45=0
.ic qb_94_45=1.8
.ic q_95_45=0
.ic qb_95_45=1.8
.ic q_96_45=0
.ic qb_96_45=1.8
.ic q_97_45=0
.ic qb_97_45=1.8
.ic q_98_45=0
.ic qb_98_45=1.8
.ic q_99_45=0
.ic qb_99_45=1.8
.ic q_0_46=0
.ic qb_0_46=1.8
.ic q_1_46=0
.ic qb_1_46=1.8
.ic q_2_46=0
.ic qb_2_46=1.8
.ic q_3_46=0
.ic qb_3_46=1.8
.ic q_4_46=0
.ic qb_4_46=1.8
.ic q_5_46=0
.ic qb_5_46=1.8
.ic q_6_46=0
.ic qb_6_46=1.8
.ic q_7_46=0
.ic qb_7_46=1.8
.ic q_8_46=0
.ic qb_8_46=1.8
.ic q_9_46=0
.ic qb_9_46=1.8
.ic q_10_46=0
.ic qb_10_46=1.8
.ic q_11_46=0
.ic qb_11_46=1.8
.ic q_12_46=0
.ic qb_12_46=1.8
.ic q_13_46=0
.ic qb_13_46=1.8
.ic q_14_46=0
.ic qb_14_46=1.8
.ic q_15_46=0
.ic qb_15_46=1.8
.ic q_16_46=0
.ic qb_16_46=1.8
.ic q_17_46=0
.ic qb_17_46=1.8
.ic q_18_46=0
.ic qb_18_46=1.8
.ic q_19_46=0
.ic qb_19_46=1.8
.ic q_20_46=0
.ic qb_20_46=1.8
.ic q_21_46=0
.ic qb_21_46=1.8
.ic q_22_46=0
.ic qb_22_46=1.8
.ic q_23_46=0
.ic qb_23_46=1.8
.ic q_24_46=0
.ic qb_24_46=1.8
.ic q_25_46=0
.ic qb_25_46=1.8
.ic q_26_46=0
.ic qb_26_46=1.8
.ic q_27_46=0
.ic qb_27_46=1.8
.ic q_28_46=0
.ic qb_28_46=1.8
.ic q_29_46=0
.ic qb_29_46=1.8
.ic q_30_46=0
.ic qb_30_46=1.8
.ic q_31_46=0
.ic qb_31_46=1.8
.ic q_32_46=0
.ic qb_32_46=1.8
.ic q_33_46=0
.ic qb_33_46=1.8
.ic q_34_46=0
.ic qb_34_46=1.8
.ic q_35_46=0
.ic qb_35_46=1.8
.ic q_36_46=0
.ic qb_36_46=1.8
.ic q_37_46=0
.ic qb_37_46=1.8
.ic q_38_46=0
.ic qb_38_46=1.8
.ic q_39_46=0
.ic qb_39_46=1.8
.ic q_40_46=0
.ic qb_40_46=1.8
.ic q_41_46=0
.ic qb_41_46=1.8
.ic q_42_46=0
.ic qb_42_46=1.8
.ic q_43_46=0
.ic qb_43_46=1.8
.ic q_44_46=0
.ic qb_44_46=1.8
.ic q_45_46=0
.ic qb_45_46=1.8
.ic q_46_46=0
.ic qb_46_46=1.8
.ic q_47_46=0
.ic qb_47_46=1.8
.ic q_48_46=0
.ic qb_48_46=1.8
.ic q_49_46=0
.ic qb_49_46=1.8
.ic q_50_46=0
.ic qb_50_46=1.8
.ic q_51_46=0
.ic qb_51_46=1.8
.ic q_52_46=0
.ic qb_52_46=1.8
.ic q_53_46=0
.ic qb_53_46=1.8
.ic q_54_46=0
.ic qb_54_46=1.8
.ic q_55_46=0
.ic qb_55_46=1.8
.ic q_56_46=0
.ic qb_56_46=1.8
.ic q_57_46=0
.ic qb_57_46=1.8
.ic q_58_46=0
.ic qb_58_46=1.8
.ic q_59_46=0
.ic qb_59_46=1.8
.ic q_60_46=0
.ic qb_60_46=1.8
.ic q_61_46=0
.ic qb_61_46=1.8
.ic q_62_46=0
.ic qb_62_46=1.8
.ic q_63_46=0
.ic qb_63_46=1.8
.ic q_64_46=0
.ic qb_64_46=1.8
.ic q_65_46=0
.ic qb_65_46=1.8
.ic q_66_46=0
.ic qb_66_46=1.8
.ic q_67_46=0
.ic qb_67_46=1.8
.ic q_68_46=0
.ic qb_68_46=1.8
.ic q_69_46=0
.ic qb_69_46=1.8
.ic q_70_46=0
.ic qb_70_46=1.8
.ic q_71_46=0
.ic qb_71_46=1.8
.ic q_72_46=0
.ic qb_72_46=1.8
.ic q_73_46=0
.ic qb_73_46=1.8
.ic q_74_46=0
.ic qb_74_46=1.8
.ic q_75_46=0
.ic qb_75_46=1.8
.ic q_76_46=0
.ic qb_76_46=1.8
.ic q_77_46=0
.ic qb_77_46=1.8
.ic q_78_46=0
.ic qb_78_46=1.8
.ic q_79_46=0
.ic qb_79_46=1.8
.ic q_80_46=0
.ic qb_80_46=1.8
.ic q_81_46=0
.ic qb_81_46=1.8
.ic q_82_46=0
.ic qb_82_46=1.8
.ic q_83_46=0
.ic qb_83_46=1.8
.ic q_84_46=0
.ic qb_84_46=1.8
.ic q_85_46=0
.ic qb_85_46=1.8
.ic q_86_46=0
.ic qb_86_46=1.8
.ic q_87_46=0
.ic qb_87_46=1.8
.ic q_88_46=0
.ic qb_88_46=1.8
.ic q_89_46=0
.ic qb_89_46=1.8
.ic q_90_46=0
.ic qb_90_46=1.8
.ic q_91_46=0
.ic qb_91_46=1.8
.ic q_92_46=0
.ic qb_92_46=1.8
.ic q_93_46=0
.ic qb_93_46=1.8
.ic q_94_46=0
.ic qb_94_46=1.8
.ic q_95_46=0
.ic qb_95_46=1.8
.ic q_96_46=0
.ic qb_96_46=1.8
.ic q_97_46=0
.ic qb_97_46=1.8
.ic q_98_46=0
.ic qb_98_46=1.8
.ic q_99_46=0
.ic qb_99_46=1.8
.ic q_0_47=0
.ic qb_0_47=1.8
.ic q_1_47=0
.ic qb_1_47=1.8
.ic q_2_47=0
.ic qb_2_47=1.8
.ic q_3_47=0
.ic qb_3_47=1.8
.ic q_4_47=0
.ic qb_4_47=1.8
.ic q_5_47=0
.ic qb_5_47=1.8
.ic q_6_47=0
.ic qb_6_47=1.8
.ic q_7_47=0
.ic qb_7_47=1.8
.ic q_8_47=0
.ic qb_8_47=1.8
.ic q_9_47=0
.ic qb_9_47=1.8
.ic q_10_47=0
.ic qb_10_47=1.8
.ic q_11_47=0
.ic qb_11_47=1.8
.ic q_12_47=0
.ic qb_12_47=1.8
.ic q_13_47=0
.ic qb_13_47=1.8
.ic q_14_47=0
.ic qb_14_47=1.8
.ic q_15_47=0
.ic qb_15_47=1.8
.ic q_16_47=0
.ic qb_16_47=1.8
.ic q_17_47=0
.ic qb_17_47=1.8
.ic q_18_47=0
.ic qb_18_47=1.8
.ic q_19_47=0
.ic qb_19_47=1.8
.ic q_20_47=0
.ic qb_20_47=1.8
.ic q_21_47=0
.ic qb_21_47=1.8
.ic q_22_47=0
.ic qb_22_47=1.8
.ic q_23_47=0
.ic qb_23_47=1.8
.ic q_24_47=0
.ic qb_24_47=1.8
.ic q_25_47=0
.ic qb_25_47=1.8
.ic q_26_47=0
.ic qb_26_47=1.8
.ic q_27_47=0
.ic qb_27_47=1.8
.ic q_28_47=0
.ic qb_28_47=1.8
.ic q_29_47=0
.ic qb_29_47=1.8
.ic q_30_47=0
.ic qb_30_47=1.8
.ic q_31_47=0
.ic qb_31_47=1.8
.ic q_32_47=0
.ic qb_32_47=1.8
.ic q_33_47=0
.ic qb_33_47=1.8
.ic q_34_47=0
.ic qb_34_47=1.8
.ic q_35_47=0
.ic qb_35_47=1.8
.ic q_36_47=0
.ic qb_36_47=1.8
.ic q_37_47=0
.ic qb_37_47=1.8
.ic q_38_47=0
.ic qb_38_47=1.8
.ic q_39_47=0
.ic qb_39_47=1.8
.ic q_40_47=0
.ic qb_40_47=1.8
.ic q_41_47=0
.ic qb_41_47=1.8
.ic q_42_47=0
.ic qb_42_47=1.8
.ic q_43_47=0
.ic qb_43_47=1.8
.ic q_44_47=0
.ic qb_44_47=1.8
.ic q_45_47=0
.ic qb_45_47=1.8
.ic q_46_47=0
.ic qb_46_47=1.8
.ic q_47_47=0
.ic qb_47_47=1.8
.ic q_48_47=0
.ic qb_48_47=1.8
.ic q_49_47=0
.ic qb_49_47=1.8
.ic q_50_47=0
.ic qb_50_47=1.8
.ic q_51_47=0
.ic qb_51_47=1.8
.ic q_52_47=0
.ic qb_52_47=1.8
.ic q_53_47=0
.ic qb_53_47=1.8
.ic q_54_47=0
.ic qb_54_47=1.8
.ic q_55_47=0
.ic qb_55_47=1.8
.ic q_56_47=0
.ic qb_56_47=1.8
.ic q_57_47=0
.ic qb_57_47=1.8
.ic q_58_47=0
.ic qb_58_47=1.8
.ic q_59_47=0
.ic qb_59_47=1.8
.ic q_60_47=0
.ic qb_60_47=1.8
.ic q_61_47=0
.ic qb_61_47=1.8
.ic q_62_47=0
.ic qb_62_47=1.8
.ic q_63_47=0
.ic qb_63_47=1.8
.ic q_64_47=0
.ic qb_64_47=1.8
.ic q_65_47=0
.ic qb_65_47=1.8
.ic q_66_47=0
.ic qb_66_47=1.8
.ic q_67_47=0
.ic qb_67_47=1.8
.ic q_68_47=0
.ic qb_68_47=1.8
.ic q_69_47=0
.ic qb_69_47=1.8
.ic q_70_47=0
.ic qb_70_47=1.8
.ic q_71_47=0
.ic qb_71_47=1.8
.ic q_72_47=0
.ic qb_72_47=1.8
.ic q_73_47=0
.ic qb_73_47=1.8
.ic q_74_47=0
.ic qb_74_47=1.8
.ic q_75_47=0
.ic qb_75_47=1.8
.ic q_76_47=0
.ic qb_76_47=1.8
.ic q_77_47=0
.ic qb_77_47=1.8
.ic q_78_47=0
.ic qb_78_47=1.8
.ic q_79_47=0
.ic qb_79_47=1.8
.ic q_80_47=0
.ic qb_80_47=1.8
.ic q_81_47=0
.ic qb_81_47=1.8
.ic q_82_47=0
.ic qb_82_47=1.8
.ic q_83_47=0
.ic qb_83_47=1.8
.ic q_84_47=0
.ic qb_84_47=1.8
.ic q_85_47=0
.ic qb_85_47=1.8
.ic q_86_47=0
.ic qb_86_47=1.8
.ic q_87_47=0
.ic qb_87_47=1.8
.ic q_88_47=0
.ic qb_88_47=1.8
.ic q_89_47=0
.ic qb_89_47=1.8
.ic q_90_47=0
.ic qb_90_47=1.8
.ic q_91_47=0
.ic qb_91_47=1.8
.ic q_92_47=0
.ic qb_92_47=1.8
.ic q_93_47=0
.ic qb_93_47=1.8
.ic q_94_47=0
.ic qb_94_47=1.8
.ic q_95_47=0
.ic qb_95_47=1.8
.ic q_96_47=0
.ic qb_96_47=1.8
.ic q_97_47=0
.ic qb_97_47=1.8
.ic q_98_47=0
.ic qb_98_47=1.8
.ic q_99_47=0
.ic qb_99_47=1.8
.ic q_0_48=0
.ic qb_0_48=1.8
.ic q_1_48=0
.ic qb_1_48=1.8
.ic q_2_48=0
.ic qb_2_48=1.8
.ic q_3_48=0
.ic qb_3_48=1.8
.ic q_4_48=0
.ic qb_4_48=1.8
.ic q_5_48=0
.ic qb_5_48=1.8
.ic q_6_48=0
.ic qb_6_48=1.8
.ic q_7_48=0
.ic qb_7_48=1.8
.ic q_8_48=0
.ic qb_8_48=1.8
.ic q_9_48=0
.ic qb_9_48=1.8
.ic q_10_48=0
.ic qb_10_48=1.8
.ic q_11_48=0
.ic qb_11_48=1.8
.ic q_12_48=0
.ic qb_12_48=1.8
.ic q_13_48=0
.ic qb_13_48=1.8
.ic q_14_48=0
.ic qb_14_48=1.8
.ic q_15_48=0
.ic qb_15_48=1.8
.ic q_16_48=0
.ic qb_16_48=1.8
.ic q_17_48=0
.ic qb_17_48=1.8
.ic q_18_48=0
.ic qb_18_48=1.8
.ic q_19_48=0
.ic qb_19_48=1.8
.ic q_20_48=0
.ic qb_20_48=1.8
.ic q_21_48=0
.ic qb_21_48=1.8
.ic q_22_48=0
.ic qb_22_48=1.8
.ic q_23_48=0
.ic qb_23_48=1.8
.ic q_24_48=0
.ic qb_24_48=1.8
.ic q_25_48=0
.ic qb_25_48=1.8
.ic q_26_48=0
.ic qb_26_48=1.8
.ic q_27_48=0
.ic qb_27_48=1.8
.ic q_28_48=0
.ic qb_28_48=1.8
.ic q_29_48=0
.ic qb_29_48=1.8
.ic q_30_48=0
.ic qb_30_48=1.8
.ic q_31_48=0
.ic qb_31_48=1.8
.ic q_32_48=0
.ic qb_32_48=1.8
.ic q_33_48=0
.ic qb_33_48=1.8
.ic q_34_48=0
.ic qb_34_48=1.8
.ic q_35_48=0
.ic qb_35_48=1.8
.ic q_36_48=0
.ic qb_36_48=1.8
.ic q_37_48=0
.ic qb_37_48=1.8
.ic q_38_48=0
.ic qb_38_48=1.8
.ic q_39_48=0
.ic qb_39_48=1.8
.ic q_40_48=0
.ic qb_40_48=1.8
.ic q_41_48=0
.ic qb_41_48=1.8
.ic q_42_48=0
.ic qb_42_48=1.8
.ic q_43_48=0
.ic qb_43_48=1.8
.ic q_44_48=0
.ic qb_44_48=1.8
.ic q_45_48=0
.ic qb_45_48=1.8
.ic q_46_48=0
.ic qb_46_48=1.8
.ic q_47_48=0
.ic qb_47_48=1.8
.ic q_48_48=0
.ic qb_48_48=1.8
.ic q_49_48=0
.ic qb_49_48=1.8
.ic q_50_48=0
.ic qb_50_48=1.8
.ic q_51_48=0
.ic qb_51_48=1.8
.ic q_52_48=0
.ic qb_52_48=1.8
.ic q_53_48=0
.ic qb_53_48=1.8
.ic q_54_48=0
.ic qb_54_48=1.8
.ic q_55_48=0
.ic qb_55_48=1.8
.ic q_56_48=0
.ic qb_56_48=1.8
.ic q_57_48=0
.ic qb_57_48=1.8
.ic q_58_48=0
.ic qb_58_48=1.8
.ic q_59_48=0
.ic qb_59_48=1.8
.ic q_60_48=0
.ic qb_60_48=1.8
.ic q_61_48=0
.ic qb_61_48=1.8
.ic q_62_48=0
.ic qb_62_48=1.8
.ic q_63_48=0
.ic qb_63_48=1.8
.ic q_64_48=0
.ic qb_64_48=1.8
.ic q_65_48=0
.ic qb_65_48=1.8
.ic q_66_48=0
.ic qb_66_48=1.8
.ic q_67_48=0
.ic qb_67_48=1.8
.ic q_68_48=0
.ic qb_68_48=1.8
.ic q_69_48=0
.ic qb_69_48=1.8
.ic q_70_48=0
.ic qb_70_48=1.8
.ic q_71_48=0
.ic qb_71_48=1.8
.ic q_72_48=0
.ic qb_72_48=1.8
.ic q_73_48=0
.ic qb_73_48=1.8
.ic q_74_48=0
.ic qb_74_48=1.8
.ic q_75_48=0
.ic qb_75_48=1.8
.ic q_76_48=0
.ic qb_76_48=1.8
.ic q_77_48=0
.ic qb_77_48=1.8
.ic q_78_48=0
.ic qb_78_48=1.8
.ic q_79_48=0
.ic qb_79_48=1.8
.ic q_80_48=0
.ic qb_80_48=1.8
.ic q_81_48=0
.ic qb_81_48=1.8
.ic q_82_48=0
.ic qb_82_48=1.8
.ic q_83_48=0
.ic qb_83_48=1.8
.ic q_84_48=0
.ic qb_84_48=1.8
.ic q_85_48=0
.ic qb_85_48=1.8
.ic q_86_48=0
.ic qb_86_48=1.8
.ic q_87_48=0
.ic qb_87_48=1.8
.ic q_88_48=0
.ic qb_88_48=1.8
.ic q_89_48=0
.ic qb_89_48=1.8
.ic q_90_48=0
.ic qb_90_48=1.8
.ic q_91_48=0
.ic qb_91_48=1.8
.ic q_92_48=0
.ic qb_92_48=1.8
.ic q_93_48=0
.ic qb_93_48=1.8
.ic q_94_48=0
.ic qb_94_48=1.8
.ic q_95_48=0
.ic qb_95_48=1.8
.ic q_96_48=0
.ic qb_96_48=1.8
.ic q_97_48=0
.ic qb_97_48=1.8
.ic q_98_48=0
.ic qb_98_48=1.8
.ic q_99_48=0
.ic qb_99_48=1.8
.ic q_0_49=0
.ic qb_0_49=1.8
.ic q_1_49=0
.ic qb_1_49=1.8
.ic q_2_49=0
.ic qb_2_49=1.8
.ic q_3_49=0
.ic qb_3_49=1.8
.ic q_4_49=0
.ic qb_4_49=1.8
.ic q_5_49=0
.ic qb_5_49=1.8
.ic q_6_49=0
.ic qb_6_49=1.8
.ic q_7_49=0
.ic qb_7_49=1.8
.ic q_8_49=0
.ic qb_8_49=1.8
.ic q_9_49=0
.ic qb_9_49=1.8
.ic q_10_49=0
.ic qb_10_49=1.8
.ic q_11_49=0
.ic qb_11_49=1.8
.ic q_12_49=0
.ic qb_12_49=1.8
.ic q_13_49=0
.ic qb_13_49=1.8
.ic q_14_49=0
.ic qb_14_49=1.8
.ic q_15_49=0
.ic qb_15_49=1.8
.ic q_16_49=0
.ic qb_16_49=1.8
.ic q_17_49=0
.ic qb_17_49=1.8
.ic q_18_49=0
.ic qb_18_49=1.8
.ic q_19_49=0
.ic qb_19_49=1.8
.ic q_20_49=0
.ic qb_20_49=1.8
.ic q_21_49=0
.ic qb_21_49=1.8
.ic q_22_49=0
.ic qb_22_49=1.8
.ic q_23_49=0
.ic qb_23_49=1.8
.ic q_24_49=0
.ic qb_24_49=1.8
.ic q_25_49=0
.ic qb_25_49=1.8
.ic q_26_49=0
.ic qb_26_49=1.8
.ic q_27_49=0
.ic qb_27_49=1.8
.ic q_28_49=0
.ic qb_28_49=1.8
.ic q_29_49=0
.ic qb_29_49=1.8
.ic q_30_49=0
.ic qb_30_49=1.8
.ic q_31_49=0
.ic qb_31_49=1.8
.ic q_32_49=0
.ic qb_32_49=1.8
.ic q_33_49=0
.ic qb_33_49=1.8
.ic q_34_49=0
.ic qb_34_49=1.8
.ic q_35_49=0
.ic qb_35_49=1.8
.ic q_36_49=0
.ic qb_36_49=1.8
.ic q_37_49=0
.ic qb_37_49=1.8
.ic q_38_49=0
.ic qb_38_49=1.8
.ic q_39_49=0
.ic qb_39_49=1.8
.ic q_40_49=0
.ic qb_40_49=1.8
.ic q_41_49=0
.ic qb_41_49=1.8
.ic q_42_49=0
.ic qb_42_49=1.8
.ic q_43_49=0
.ic qb_43_49=1.8
.ic q_44_49=0
.ic qb_44_49=1.8
.ic q_45_49=0
.ic qb_45_49=1.8
.ic q_46_49=0
.ic qb_46_49=1.8
.ic q_47_49=0
.ic qb_47_49=1.8
.ic q_48_49=0
.ic qb_48_49=1.8
.ic q_49_49=0
.ic qb_49_49=1.8
.ic q_50_49=0
.ic qb_50_49=1.8
.ic q_51_49=0
.ic qb_51_49=1.8
.ic q_52_49=0
.ic qb_52_49=1.8
.ic q_53_49=0
.ic qb_53_49=1.8
.ic q_54_49=0
.ic qb_54_49=1.8
.ic q_55_49=0
.ic qb_55_49=1.8
.ic q_56_49=0
.ic qb_56_49=1.8
.ic q_57_49=0
.ic qb_57_49=1.8
.ic q_58_49=0
.ic qb_58_49=1.8
.ic q_59_49=0
.ic qb_59_49=1.8
.ic q_60_49=0
.ic qb_60_49=1.8
.ic q_61_49=0
.ic qb_61_49=1.8
.ic q_62_49=0
.ic qb_62_49=1.8
.ic q_63_49=0
.ic qb_63_49=1.8
.ic q_64_49=0
.ic qb_64_49=1.8
.ic q_65_49=0
.ic qb_65_49=1.8
.ic q_66_49=0
.ic qb_66_49=1.8
.ic q_67_49=0
.ic qb_67_49=1.8
.ic q_68_49=0
.ic qb_68_49=1.8
.ic q_69_49=0
.ic qb_69_49=1.8
.ic q_70_49=0
.ic qb_70_49=1.8
.ic q_71_49=0
.ic qb_71_49=1.8
.ic q_72_49=0
.ic qb_72_49=1.8
.ic q_73_49=0
.ic qb_73_49=1.8
.ic q_74_49=0
.ic qb_74_49=1.8
.ic q_75_49=0
.ic qb_75_49=1.8
.ic q_76_49=0
.ic qb_76_49=1.8
.ic q_77_49=0
.ic qb_77_49=1.8
.ic q_78_49=0
.ic qb_78_49=1.8
.ic q_79_49=0
.ic qb_79_49=1.8
.ic q_80_49=0
.ic qb_80_49=1.8
.ic q_81_49=0
.ic qb_81_49=1.8
.ic q_82_49=0
.ic qb_82_49=1.8
.ic q_83_49=0
.ic qb_83_49=1.8
.ic q_84_49=0
.ic qb_84_49=1.8
.ic q_85_49=0
.ic qb_85_49=1.8
.ic q_86_49=0
.ic qb_86_49=1.8
.ic q_87_49=0
.ic qb_87_49=1.8
.ic q_88_49=0
.ic qb_88_49=1.8
.ic q_89_49=0
.ic qb_89_49=1.8
.ic q_90_49=0
.ic qb_90_49=1.8
.ic q_91_49=0
.ic qb_91_49=1.8
.ic q_92_49=0
.ic qb_92_49=1.8
.ic q_93_49=0
.ic qb_93_49=1.8
.ic q_94_49=0
.ic qb_94_49=1.8
.ic q_95_49=0
.ic qb_95_49=1.8
.ic q_96_49=0
.ic qb_96_49=1.8
.ic q_97_49=0
.ic qb_97_49=1.8
.ic q_98_49=0
.ic qb_98_49=1.8
.ic q_99_49=0
.ic qb_99_49=1.8
.ic q_0_50=0
.ic qb_0_50=1.8
.ic q_1_50=0
.ic qb_1_50=1.8
.ic q_2_50=0
.ic qb_2_50=1.8
.ic q_3_50=0
.ic qb_3_50=1.8
.ic q_4_50=0
.ic qb_4_50=1.8
.ic q_5_50=0
.ic qb_5_50=1.8
.ic q_6_50=0
.ic qb_6_50=1.8
.ic q_7_50=0
.ic qb_7_50=1.8
.ic q_8_50=0
.ic qb_8_50=1.8
.ic q_9_50=0
.ic qb_9_50=1.8
.ic q_10_50=0
.ic qb_10_50=1.8
.ic q_11_50=0
.ic qb_11_50=1.8
.ic q_12_50=0
.ic qb_12_50=1.8
.ic q_13_50=0
.ic qb_13_50=1.8
.ic q_14_50=0
.ic qb_14_50=1.8
.ic q_15_50=0
.ic qb_15_50=1.8
.ic q_16_50=0
.ic qb_16_50=1.8
.ic q_17_50=0
.ic qb_17_50=1.8
.ic q_18_50=0
.ic qb_18_50=1.8
.ic q_19_50=0
.ic qb_19_50=1.8
.ic q_20_50=0
.ic qb_20_50=1.8
.ic q_21_50=0
.ic qb_21_50=1.8
.ic q_22_50=0
.ic qb_22_50=1.8
.ic q_23_50=0
.ic qb_23_50=1.8
.ic q_24_50=0
.ic qb_24_50=1.8
.ic q_25_50=0
.ic qb_25_50=1.8
.ic q_26_50=0
.ic qb_26_50=1.8
.ic q_27_50=0
.ic qb_27_50=1.8
.ic q_28_50=0
.ic qb_28_50=1.8
.ic q_29_50=0
.ic qb_29_50=1.8
.ic q_30_50=0
.ic qb_30_50=1.8
.ic q_31_50=0
.ic qb_31_50=1.8
.ic q_32_50=0
.ic qb_32_50=1.8
.ic q_33_50=0
.ic qb_33_50=1.8
.ic q_34_50=0
.ic qb_34_50=1.8
.ic q_35_50=0
.ic qb_35_50=1.8
.ic q_36_50=0
.ic qb_36_50=1.8
.ic q_37_50=0
.ic qb_37_50=1.8
.ic q_38_50=0
.ic qb_38_50=1.8
.ic q_39_50=0
.ic qb_39_50=1.8
.ic q_40_50=0
.ic qb_40_50=1.8
.ic q_41_50=0
.ic qb_41_50=1.8
.ic q_42_50=0
.ic qb_42_50=1.8
.ic q_43_50=0
.ic qb_43_50=1.8
.ic q_44_50=0
.ic qb_44_50=1.8
.ic q_45_50=0
.ic qb_45_50=1.8
.ic q_46_50=0
.ic qb_46_50=1.8
.ic q_47_50=0
.ic qb_47_50=1.8
.ic q_48_50=0
.ic qb_48_50=1.8
.ic q_49_50=0
.ic qb_49_50=1.8
.ic q_50_50=0
.ic qb_50_50=1.8
.ic q_51_50=0
.ic qb_51_50=1.8
.ic q_52_50=0
.ic qb_52_50=1.8
.ic q_53_50=0
.ic qb_53_50=1.8
.ic q_54_50=0
.ic qb_54_50=1.8
.ic q_55_50=0
.ic qb_55_50=1.8
.ic q_56_50=0
.ic qb_56_50=1.8
.ic q_57_50=0
.ic qb_57_50=1.8
.ic q_58_50=0
.ic qb_58_50=1.8
.ic q_59_50=0
.ic qb_59_50=1.8
.ic q_60_50=0
.ic qb_60_50=1.8
.ic q_61_50=0
.ic qb_61_50=1.8
.ic q_62_50=0
.ic qb_62_50=1.8
.ic q_63_50=0
.ic qb_63_50=1.8
.ic q_64_50=0
.ic qb_64_50=1.8
.ic q_65_50=0
.ic qb_65_50=1.8
.ic q_66_50=0
.ic qb_66_50=1.8
.ic q_67_50=0
.ic qb_67_50=1.8
.ic q_68_50=0
.ic qb_68_50=1.8
.ic q_69_50=0
.ic qb_69_50=1.8
.ic q_70_50=0
.ic qb_70_50=1.8
.ic q_71_50=0
.ic qb_71_50=1.8
.ic q_72_50=0
.ic qb_72_50=1.8
.ic q_73_50=0
.ic qb_73_50=1.8
.ic q_74_50=0
.ic qb_74_50=1.8
.ic q_75_50=0
.ic qb_75_50=1.8
.ic q_76_50=0
.ic qb_76_50=1.8
.ic q_77_50=0
.ic qb_77_50=1.8
.ic q_78_50=0
.ic qb_78_50=1.8
.ic q_79_50=0
.ic qb_79_50=1.8
.ic q_80_50=0
.ic qb_80_50=1.8
.ic q_81_50=0
.ic qb_81_50=1.8
.ic q_82_50=0
.ic qb_82_50=1.8
.ic q_83_50=0
.ic qb_83_50=1.8
.ic q_84_50=0
.ic qb_84_50=1.8
.ic q_85_50=0
.ic qb_85_50=1.8
.ic q_86_50=0
.ic qb_86_50=1.8
.ic q_87_50=0
.ic qb_87_50=1.8
.ic q_88_50=0
.ic qb_88_50=1.8
.ic q_89_50=0
.ic qb_89_50=1.8
.ic q_90_50=0
.ic qb_90_50=1.8
.ic q_91_50=0
.ic qb_91_50=1.8
.ic q_92_50=0
.ic qb_92_50=1.8
.ic q_93_50=0
.ic qb_93_50=1.8
.ic q_94_50=0
.ic qb_94_50=1.8
.ic q_95_50=0
.ic qb_95_50=1.8
.ic q_96_50=0
.ic qb_96_50=1.8
.ic q_97_50=0
.ic qb_97_50=1.8
.ic q_98_50=0
.ic qb_98_50=1.8
.ic q_99_50=0
.ic qb_99_50=1.8
.ic q_0_51=0
.ic qb_0_51=1.8
.ic q_1_51=0
.ic qb_1_51=1.8
.ic q_2_51=0
.ic qb_2_51=1.8
.ic q_3_51=0
.ic qb_3_51=1.8
.ic q_4_51=0
.ic qb_4_51=1.8
.ic q_5_51=0
.ic qb_5_51=1.8
.ic q_6_51=0
.ic qb_6_51=1.8
.ic q_7_51=0
.ic qb_7_51=1.8
.ic q_8_51=0
.ic qb_8_51=1.8
.ic q_9_51=0
.ic qb_9_51=1.8
.ic q_10_51=0
.ic qb_10_51=1.8
.ic q_11_51=0
.ic qb_11_51=1.8
.ic q_12_51=0
.ic qb_12_51=1.8
.ic q_13_51=0
.ic qb_13_51=1.8
.ic q_14_51=0
.ic qb_14_51=1.8
.ic q_15_51=0
.ic qb_15_51=1.8
.ic q_16_51=0
.ic qb_16_51=1.8
.ic q_17_51=0
.ic qb_17_51=1.8
.ic q_18_51=0
.ic qb_18_51=1.8
.ic q_19_51=0
.ic qb_19_51=1.8
.ic q_20_51=0
.ic qb_20_51=1.8
.ic q_21_51=0
.ic qb_21_51=1.8
.ic q_22_51=0
.ic qb_22_51=1.8
.ic q_23_51=0
.ic qb_23_51=1.8
.ic q_24_51=0
.ic qb_24_51=1.8
.ic q_25_51=0
.ic qb_25_51=1.8
.ic q_26_51=0
.ic qb_26_51=1.8
.ic q_27_51=0
.ic qb_27_51=1.8
.ic q_28_51=0
.ic qb_28_51=1.8
.ic q_29_51=0
.ic qb_29_51=1.8
.ic q_30_51=0
.ic qb_30_51=1.8
.ic q_31_51=0
.ic qb_31_51=1.8
.ic q_32_51=0
.ic qb_32_51=1.8
.ic q_33_51=0
.ic qb_33_51=1.8
.ic q_34_51=0
.ic qb_34_51=1.8
.ic q_35_51=0
.ic qb_35_51=1.8
.ic q_36_51=0
.ic qb_36_51=1.8
.ic q_37_51=0
.ic qb_37_51=1.8
.ic q_38_51=0
.ic qb_38_51=1.8
.ic q_39_51=0
.ic qb_39_51=1.8
.ic q_40_51=0
.ic qb_40_51=1.8
.ic q_41_51=0
.ic qb_41_51=1.8
.ic q_42_51=0
.ic qb_42_51=1.8
.ic q_43_51=0
.ic qb_43_51=1.8
.ic q_44_51=0
.ic qb_44_51=1.8
.ic q_45_51=0
.ic qb_45_51=1.8
.ic q_46_51=0
.ic qb_46_51=1.8
.ic q_47_51=0
.ic qb_47_51=1.8
.ic q_48_51=0
.ic qb_48_51=1.8
.ic q_49_51=0
.ic qb_49_51=1.8
.ic q_50_51=0
.ic qb_50_51=1.8
.ic q_51_51=0
.ic qb_51_51=1.8
.ic q_52_51=0
.ic qb_52_51=1.8
.ic q_53_51=0
.ic qb_53_51=1.8
.ic q_54_51=0
.ic qb_54_51=1.8
.ic q_55_51=0
.ic qb_55_51=1.8
.ic q_56_51=0
.ic qb_56_51=1.8
.ic q_57_51=0
.ic qb_57_51=1.8
.ic q_58_51=0
.ic qb_58_51=1.8
.ic q_59_51=0
.ic qb_59_51=1.8
.ic q_60_51=0
.ic qb_60_51=1.8
.ic q_61_51=0
.ic qb_61_51=1.8
.ic q_62_51=0
.ic qb_62_51=1.8
.ic q_63_51=0
.ic qb_63_51=1.8
.ic q_64_51=0
.ic qb_64_51=1.8
.ic q_65_51=0
.ic qb_65_51=1.8
.ic q_66_51=0
.ic qb_66_51=1.8
.ic q_67_51=0
.ic qb_67_51=1.8
.ic q_68_51=0
.ic qb_68_51=1.8
.ic q_69_51=0
.ic qb_69_51=1.8
.ic q_70_51=0
.ic qb_70_51=1.8
.ic q_71_51=0
.ic qb_71_51=1.8
.ic q_72_51=0
.ic qb_72_51=1.8
.ic q_73_51=0
.ic qb_73_51=1.8
.ic q_74_51=0
.ic qb_74_51=1.8
.ic q_75_51=0
.ic qb_75_51=1.8
.ic q_76_51=0
.ic qb_76_51=1.8
.ic q_77_51=0
.ic qb_77_51=1.8
.ic q_78_51=0
.ic qb_78_51=1.8
.ic q_79_51=0
.ic qb_79_51=1.8
.ic q_80_51=0
.ic qb_80_51=1.8
.ic q_81_51=0
.ic qb_81_51=1.8
.ic q_82_51=0
.ic qb_82_51=1.8
.ic q_83_51=0
.ic qb_83_51=1.8
.ic q_84_51=0
.ic qb_84_51=1.8
.ic q_85_51=0
.ic qb_85_51=1.8
.ic q_86_51=0
.ic qb_86_51=1.8
.ic q_87_51=0
.ic qb_87_51=1.8
.ic q_88_51=0
.ic qb_88_51=1.8
.ic q_89_51=0
.ic qb_89_51=1.8
.ic q_90_51=0
.ic qb_90_51=1.8
.ic q_91_51=0
.ic qb_91_51=1.8
.ic q_92_51=0
.ic qb_92_51=1.8
.ic q_93_51=0
.ic qb_93_51=1.8
.ic q_94_51=0
.ic qb_94_51=1.8
.ic q_95_51=0
.ic qb_95_51=1.8
.ic q_96_51=0
.ic qb_96_51=1.8
.ic q_97_51=0
.ic qb_97_51=1.8
.ic q_98_51=0
.ic qb_98_51=1.8
.ic q_99_51=0
.ic qb_99_51=1.8
.ic q_0_52=0
.ic qb_0_52=1.8
.ic q_1_52=0
.ic qb_1_52=1.8
.ic q_2_52=0
.ic qb_2_52=1.8
.ic q_3_52=0
.ic qb_3_52=1.8
.ic q_4_52=0
.ic qb_4_52=1.8
.ic q_5_52=0
.ic qb_5_52=1.8
.ic q_6_52=0
.ic qb_6_52=1.8
.ic q_7_52=0
.ic qb_7_52=1.8
.ic q_8_52=0
.ic qb_8_52=1.8
.ic q_9_52=0
.ic qb_9_52=1.8
.ic q_10_52=0
.ic qb_10_52=1.8
.ic q_11_52=0
.ic qb_11_52=1.8
.ic q_12_52=0
.ic qb_12_52=1.8
.ic q_13_52=0
.ic qb_13_52=1.8
.ic q_14_52=0
.ic qb_14_52=1.8
.ic q_15_52=0
.ic qb_15_52=1.8
.ic q_16_52=0
.ic qb_16_52=1.8
.ic q_17_52=0
.ic qb_17_52=1.8
.ic q_18_52=0
.ic qb_18_52=1.8
.ic q_19_52=0
.ic qb_19_52=1.8
.ic q_20_52=0
.ic qb_20_52=1.8
.ic q_21_52=0
.ic qb_21_52=1.8
.ic q_22_52=0
.ic qb_22_52=1.8
.ic q_23_52=0
.ic qb_23_52=1.8
.ic q_24_52=0
.ic qb_24_52=1.8
.ic q_25_52=0
.ic qb_25_52=1.8
.ic q_26_52=0
.ic qb_26_52=1.8
.ic q_27_52=0
.ic qb_27_52=1.8
.ic q_28_52=0
.ic qb_28_52=1.8
.ic q_29_52=0
.ic qb_29_52=1.8
.ic q_30_52=0
.ic qb_30_52=1.8
.ic q_31_52=0
.ic qb_31_52=1.8
.ic q_32_52=0
.ic qb_32_52=1.8
.ic q_33_52=0
.ic qb_33_52=1.8
.ic q_34_52=0
.ic qb_34_52=1.8
.ic q_35_52=0
.ic qb_35_52=1.8
.ic q_36_52=0
.ic qb_36_52=1.8
.ic q_37_52=0
.ic qb_37_52=1.8
.ic q_38_52=0
.ic qb_38_52=1.8
.ic q_39_52=0
.ic qb_39_52=1.8
.ic q_40_52=0
.ic qb_40_52=1.8
.ic q_41_52=0
.ic qb_41_52=1.8
.ic q_42_52=0
.ic qb_42_52=1.8
.ic q_43_52=0
.ic qb_43_52=1.8
.ic q_44_52=0
.ic qb_44_52=1.8
.ic q_45_52=0
.ic qb_45_52=1.8
.ic q_46_52=0
.ic qb_46_52=1.8
.ic q_47_52=0
.ic qb_47_52=1.8
.ic q_48_52=0
.ic qb_48_52=1.8
.ic q_49_52=0
.ic qb_49_52=1.8
.ic q_50_52=0
.ic qb_50_52=1.8
.ic q_51_52=0
.ic qb_51_52=1.8
.ic q_52_52=0
.ic qb_52_52=1.8
.ic q_53_52=0
.ic qb_53_52=1.8
.ic q_54_52=0
.ic qb_54_52=1.8
.ic q_55_52=0
.ic qb_55_52=1.8
.ic q_56_52=0
.ic qb_56_52=1.8
.ic q_57_52=0
.ic qb_57_52=1.8
.ic q_58_52=0
.ic qb_58_52=1.8
.ic q_59_52=0
.ic qb_59_52=1.8
.ic q_60_52=0
.ic qb_60_52=1.8
.ic q_61_52=0
.ic qb_61_52=1.8
.ic q_62_52=0
.ic qb_62_52=1.8
.ic q_63_52=0
.ic qb_63_52=1.8
.ic q_64_52=0
.ic qb_64_52=1.8
.ic q_65_52=0
.ic qb_65_52=1.8
.ic q_66_52=0
.ic qb_66_52=1.8
.ic q_67_52=0
.ic qb_67_52=1.8
.ic q_68_52=0
.ic qb_68_52=1.8
.ic q_69_52=0
.ic qb_69_52=1.8
.ic q_70_52=0
.ic qb_70_52=1.8
.ic q_71_52=0
.ic qb_71_52=1.8
.ic q_72_52=0
.ic qb_72_52=1.8
.ic q_73_52=0
.ic qb_73_52=1.8
.ic q_74_52=0
.ic qb_74_52=1.8
.ic q_75_52=0
.ic qb_75_52=1.8
.ic q_76_52=0
.ic qb_76_52=1.8
.ic q_77_52=0
.ic qb_77_52=1.8
.ic q_78_52=0
.ic qb_78_52=1.8
.ic q_79_52=0
.ic qb_79_52=1.8
.ic q_80_52=0
.ic qb_80_52=1.8
.ic q_81_52=0
.ic qb_81_52=1.8
.ic q_82_52=0
.ic qb_82_52=1.8
.ic q_83_52=0
.ic qb_83_52=1.8
.ic q_84_52=0
.ic qb_84_52=1.8
.ic q_85_52=0
.ic qb_85_52=1.8
.ic q_86_52=0
.ic qb_86_52=1.8
.ic q_87_52=0
.ic qb_87_52=1.8
.ic q_88_52=0
.ic qb_88_52=1.8
.ic q_89_52=0
.ic qb_89_52=1.8
.ic q_90_52=0
.ic qb_90_52=1.8
.ic q_91_52=0
.ic qb_91_52=1.8
.ic q_92_52=0
.ic qb_92_52=1.8
.ic q_93_52=0
.ic qb_93_52=1.8
.ic q_94_52=0
.ic qb_94_52=1.8
.ic q_95_52=0
.ic qb_95_52=1.8
.ic q_96_52=0
.ic qb_96_52=1.8
.ic q_97_52=0
.ic qb_97_52=1.8
.ic q_98_52=0
.ic qb_98_52=1.8
.ic q_99_52=0
.ic qb_99_52=1.8
.ic q_0_53=0
.ic qb_0_53=1.8
.ic q_1_53=0
.ic qb_1_53=1.8
.ic q_2_53=0
.ic qb_2_53=1.8
.ic q_3_53=0
.ic qb_3_53=1.8
.ic q_4_53=0
.ic qb_4_53=1.8
.ic q_5_53=0
.ic qb_5_53=1.8
.ic q_6_53=0
.ic qb_6_53=1.8
.ic q_7_53=0
.ic qb_7_53=1.8
.ic q_8_53=0
.ic qb_8_53=1.8
.ic q_9_53=0
.ic qb_9_53=1.8
.ic q_10_53=0
.ic qb_10_53=1.8
.ic q_11_53=0
.ic qb_11_53=1.8
.ic q_12_53=0
.ic qb_12_53=1.8
.ic q_13_53=0
.ic qb_13_53=1.8
.ic q_14_53=0
.ic qb_14_53=1.8
.ic q_15_53=0
.ic qb_15_53=1.8
.ic q_16_53=0
.ic qb_16_53=1.8
.ic q_17_53=0
.ic qb_17_53=1.8
.ic q_18_53=0
.ic qb_18_53=1.8
.ic q_19_53=0
.ic qb_19_53=1.8
.ic q_20_53=0
.ic qb_20_53=1.8
.ic q_21_53=0
.ic qb_21_53=1.8
.ic q_22_53=0
.ic qb_22_53=1.8
.ic q_23_53=0
.ic qb_23_53=1.8
.ic q_24_53=0
.ic qb_24_53=1.8
.ic q_25_53=0
.ic qb_25_53=1.8
.ic q_26_53=0
.ic qb_26_53=1.8
.ic q_27_53=0
.ic qb_27_53=1.8
.ic q_28_53=0
.ic qb_28_53=1.8
.ic q_29_53=0
.ic qb_29_53=1.8
.ic q_30_53=0
.ic qb_30_53=1.8
.ic q_31_53=0
.ic qb_31_53=1.8
.ic q_32_53=0
.ic qb_32_53=1.8
.ic q_33_53=0
.ic qb_33_53=1.8
.ic q_34_53=0
.ic qb_34_53=1.8
.ic q_35_53=0
.ic qb_35_53=1.8
.ic q_36_53=0
.ic qb_36_53=1.8
.ic q_37_53=0
.ic qb_37_53=1.8
.ic q_38_53=0
.ic qb_38_53=1.8
.ic q_39_53=0
.ic qb_39_53=1.8
.ic q_40_53=0
.ic qb_40_53=1.8
.ic q_41_53=0
.ic qb_41_53=1.8
.ic q_42_53=0
.ic qb_42_53=1.8
.ic q_43_53=0
.ic qb_43_53=1.8
.ic q_44_53=0
.ic qb_44_53=1.8
.ic q_45_53=0
.ic qb_45_53=1.8
.ic q_46_53=0
.ic qb_46_53=1.8
.ic q_47_53=0
.ic qb_47_53=1.8
.ic q_48_53=0
.ic qb_48_53=1.8
.ic q_49_53=0
.ic qb_49_53=1.8
.ic q_50_53=0
.ic qb_50_53=1.8
.ic q_51_53=0
.ic qb_51_53=1.8
.ic q_52_53=0
.ic qb_52_53=1.8
.ic q_53_53=0
.ic qb_53_53=1.8
.ic q_54_53=0
.ic qb_54_53=1.8
.ic q_55_53=0
.ic qb_55_53=1.8
.ic q_56_53=0
.ic qb_56_53=1.8
.ic q_57_53=0
.ic qb_57_53=1.8
.ic q_58_53=0
.ic qb_58_53=1.8
.ic q_59_53=0
.ic qb_59_53=1.8
.ic q_60_53=0
.ic qb_60_53=1.8
.ic q_61_53=0
.ic qb_61_53=1.8
.ic q_62_53=0
.ic qb_62_53=1.8
.ic q_63_53=0
.ic qb_63_53=1.8
.ic q_64_53=0
.ic qb_64_53=1.8
.ic q_65_53=0
.ic qb_65_53=1.8
.ic q_66_53=0
.ic qb_66_53=1.8
.ic q_67_53=0
.ic qb_67_53=1.8
.ic q_68_53=0
.ic qb_68_53=1.8
.ic q_69_53=0
.ic qb_69_53=1.8
.ic q_70_53=0
.ic qb_70_53=1.8
.ic q_71_53=0
.ic qb_71_53=1.8
.ic q_72_53=0
.ic qb_72_53=1.8
.ic q_73_53=0
.ic qb_73_53=1.8
.ic q_74_53=0
.ic qb_74_53=1.8
.ic q_75_53=0
.ic qb_75_53=1.8
.ic q_76_53=0
.ic qb_76_53=1.8
.ic q_77_53=0
.ic qb_77_53=1.8
.ic q_78_53=0
.ic qb_78_53=1.8
.ic q_79_53=0
.ic qb_79_53=1.8
.ic q_80_53=0
.ic qb_80_53=1.8
.ic q_81_53=0
.ic qb_81_53=1.8
.ic q_82_53=0
.ic qb_82_53=1.8
.ic q_83_53=0
.ic qb_83_53=1.8
.ic q_84_53=0
.ic qb_84_53=1.8
.ic q_85_53=0
.ic qb_85_53=1.8
.ic q_86_53=0
.ic qb_86_53=1.8
.ic q_87_53=0
.ic qb_87_53=1.8
.ic q_88_53=0
.ic qb_88_53=1.8
.ic q_89_53=0
.ic qb_89_53=1.8
.ic q_90_53=0
.ic qb_90_53=1.8
.ic q_91_53=0
.ic qb_91_53=1.8
.ic q_92_53=0
.ic qb_92_53=1.8
.ic q_93_53=0
.ic qb_93_53=1.8
.ic q_94_53=0
.ic qb_94_53=1.8
.ic q_95_53=0
.ic qb_95_53=1.8
.ic q_96_53=0
.ic qb_96_53=1.8
.ic q_97_53=0
.ic qb_97_53=1.8
.ic q_98_53=0
.ic qb_98_53=1.8
.ic q_99_53=0
.ic qb_99_53=1.8
.ic q_0_54=0
.ic qb_0_54=1.8
.ic q_1_54=0
.ic qb_1_54=1.8
.ic q_2_54=0
.ic qb_2_54=1.8
.ic q_3_54=0
.ic qb_3_54=1.8
.ic q_4_54=0
.ic qb_4_54=1.8
.ic q_5_54=0
.ic qb_5_54=1.8
.ic q_6_54=0
.ic qb_6_54=1.8
.ic q_7_54=0
.ic qb_7_54=1.8
.ic q_8_54=0
.ic qb_8_54=1.8
.ic q_9_54=0
.ic qb_9_54=1.8
.ic q_10_54=0
.ic qb_10_54=1.8
.ic q_11_54=0
.ic qb_11_54=1.8
.ic q_12_54=0
.ic qb_12_54=1.8
.ic q_13_54=0
.ic qb_13_54=1.8
.ic q_14_54=0
.ic qb_14_54=1.8
.ic q_15_54=0
.ic qb_15_54=1.8
.ic q_16_54=0
.ic qb_16_54=1.8
.ic q_17_54=0
.ic qb_17_54=1.8
.ic q_18_54=0
.ic qb_18_54=1.8
.ic q_19_54=0
.ic qb_19_54=1.8
.ic q_20_54=0
.ic qb_20_54=1.8
.ic q_21_54=0
.ic qb_21_54=1.8
.ic q_22_54=0
.ic qb_22_54=1.8
.ic q_23_54=0
.ic qb_23_54=1.8
.ic q_24_54=0
.ic qb_24_54=1.8
.ic q_25_54=0
.ic qb_25_54=1.8
.ic q_26_54=0
.ic qb_26_54=1.8
.ic q_27_54=0
.ic qb_27_54=1.8
.ic q_28_54=0
.ic qb_28_54=1.8
.ic q_29_54=0
.ic qb_29_54=1.8
.ic q_30_54=0
.ic qb_30_54=1.8
.ic q_31_54=0
.ic qb_31_54=1.8
.ic q_32_54=0
.ic qb_32_54=1.8
.ic q_33_54=0
.ic qb_33_54=1.8
.ic q_34_54=0
.ic qb_34_54=1.8
.ic q_35_54=0
.ic qb_35_54=1.8
.ic q_36_54=0
.ic qb_36_54=1.8
.ic q_37_54=0
.ic qb_37_54=1.8
.ic q_38_54=0
.ic qb_38_54=1.8
.ic q_39_54=0
.ic qb_39_54=1.8
.ic q_40_54=0
.ic qb_40_54=1.8
.ic q_41_54=0
.ic qb_41_54=1.8
.ic q_42_54=0
.ic qb_42_54=1.8
.ic q_43_54=0
.ic qb_43_54=1.8
.ic q_44_54=0
.ic qb_44_54=1.8
.ic q_45_54=0
.ic qb_45_54=1.8
.ic q_46_54=0
.ic qb_46_54=1.8
.ic q_47_54=0
.ic qb_47_54=1.8
.ic q_48_54=0
.ic qb_48_54=1.8
.ic q_49_54=0
.ic qb_49_54=1.8
.ic q_50_54=0
.ic qb_50_54=1.8
.ic q_51_54=0
.ic qb_51_54=1.8
.ic q_52_54=0
.ic qb_52_54=1.8
.ic q_53_54=0
.ic qb_53_54=1.8
.ic q_54_54=0
.ic qb_54_54=1.8
.ic q_55_54=0
.ic qb_55_54=1.8
.ic q_56_54=0
.ic qb_56_54=1.8
.ic q_57_54=0
.ic qb_57_54=1.8
.ic q_58_54=0
.ic qb_58_54=1.8
.ic q_59_54=0
.ic qb_59_54=1.8
.ic q_60_54=0
.ic qb_60_54=1.8
.ic q_61_54=0
.ic qb_61_54=1.8
.ic q_62_54=0
.ic qb_62_54=1.8
.ic q_63_54=0
.ic qb_63_54=1.8
.ic q_64_54=0
.ic qb_64_54=1.8
.ic q_65_54=0
.ic qb_65_54=1.8
.ic q_66_54=0
.ic qb_66_54=1.8
.ic q_67_54=0
.ic qb_67_54=1.8
.ic q_68_54=0
.ic qb_68_54=1.8
.ic q_69_54=0
.ic qb_69_54=1.8
.ic q_70_54=0
.ic qb_70_54=1.8
.ic q_71_54=0
.ic qb_71_54=1.8
.ic q_72_54=0
.ic qb_72_54=1.8
.ic q_73_54=0
.ic qb_73_54=1.8
.ic q_74_54=0
.ic qb_74_54=1.8
.ic q_75_54=0
.ic qb_75_54=1.8
.ic q_76_54=0
.ic qb_76_54=1.8
.ic q_77_54=0
.ic qb_77_54=1.8
.ic q_78_54=0
.ic qb_78_54=1.8
.ic q_79_54=0
.ic qb_79_54=1.8
.ic q_80_54=0
.ic qb_80_54=1.8
.ic q_81_54=0
.ic qb_81_54=1.8
.ic q_82_54=0
.ic qb_82_54=1.8
.ic q_83_54=0
.ic qb_83_54=1.8
.ic q_84_54=0
.ic qb_84_54=1.8
.ic q_85_54=0
.ic qb_85_54=1.8
.ic q_86_54=0
.ic qb_86_54=1.8
.ic q_87_54=0
.ic qb_87_54=1.8
.ic q_88_54=0
.ic qb_88_54=1.8
.ic q_89_54=0
.ic qb_89_54=1.8
.ic q_90_54=0
.ic qb_90_54=1.8
.ic q_91_54=0
.ic qb_91_54=1.8
.ic q_92_54=0
.ic qb_92_54=1.8
.ic q_93_54=0
.ic qb_93_54=1.8
.ic q_94_54=0
.ic qb_94_54=1.8
.ic q_95_54=0
.ic qb_95_54=1.8
.ic q_96_54=0
.ic qb_96_54=1.8
.ic q_97_54=0
.ic qb_97_54=1.8
.ic q_98_54=0
.ic qb_98_54=1.8
.ic q_99_54=0
.ic qb_99_54=1.8
.ic q_0_55=0
.ic qb_0_55=1.8
.ic q_1_55=0
.ic qb_1_55=1.8
.ic q_2_55=0
.ic qb_2_55=1.8
.ic q_3_55=0
.ic qb_3_55=1.8
.ic q_4_55=0
.ic qb_4_55=1.8
.ic q_5_55=0
.ic qb_5_55=1.8
.ic q_6_55=0
.ic qb_6_55=1.8
.ic q_7_55=0
.ic qb_7_55=1.8
.ic q_8_55=0
.ic qb_8_55=1.8
.ic q_9_55=0
.ic qb_9_55=1.8
.ic q_10_55=0
.ic qb_10_55=1.8
.ic q_11_55=0
.ic qb_11_55=1.8
.ic q_12_55=0
.ic qb_12_55=1.8
.ic q_13_55=0
.ic qb_13_55=1.8
.ic q_14_55=0
.ic qb_14_55=1.8
.ic q_15_55=0
.ic qb_15_55=1.8
.ic q_16_55=0
.ic qb_16_55=1.8
.ic q_17_55=0
.ic qb_17_55=1.8
.ic q_18_55=0
.ic qb_18_55=1.8
.ic q_19_55=0
.ic qb_19_55=1.8
.ic q_20_55=0
.ic qb_20_55=1.8
.ic q_21_55=0
.ic qb_21_55=1.8
.ic q_22_55=0
.ic qb_22_55=1.8
.ic q_23_55=0
.ic qb_23_55=1.8
.ic q_24_55=0
.ic qb_24_55=1.8
.ic q_25_55=0
.ic qb_25_55=1.8
.ic q_26_55=0
.ic qb_26_55=1.8
.ic q_27_55=0
.ic qb_27_55=1.8
.ic q_28_55=0
.ic qb_28_55=1.8
.ic q_29_55=0
.ic qb_29_55=1.8
.ic q_30_55=0
.ic qb_30_55=1.8
.ic q_31_55=0
.ic qb_31_55=1.8
.ic q_32_55=0
.ic qb_32_55=1.8
.ic q_33_55=0
.ic qb_33_55=1.8
.ic q_34_55=0
.ic qb_34_55=1.8
.ic q_35_55=0
.ic qb_35_55=1.8
.ic q_36_55=0
.ic qb_36_55=1.8
.ic q_37_55=0
.ic qb_37_55=1.8
.ic q_38_55=0
.ic qb_38_55=1.8
.ic q_39_55=0
.ic qb_39_55=1.8
.ic q_40_55=0
.ic qb_40_55=1.8
.ic q_41_55=0
.ic qb_41_55=1.8
.ic q_42_55=0
.ic qb_42_55=1.8
.ic q_43_55=0
.ic qb_43_55=1.8
.ic q_44_55=0
.ic qb_44_55=1.8
.ic q_45_55=0
.ic qb_45_55=1.8
.ic q_46_55=0
.ic qb_46_55=1.8
.ic q_47_55=0
.ic qb_47_55=1.8
.ic q_48_55=0
.ic qb_48_55=1.8
.ic q_49_55=0
.ic qb_49_55=1.8
.ic q_50_55=0
.ic qb_50_55=1.8
.ic q_51_55=0
.ic qb_51_55=1.8
.ic q_52_55=0
.ic qb_52_55=1.8
.ic q_53_55=0
.ic qb_53_55=1.8
.ic q_54_55=0
.ic qb_54_55=1.8
.ic q_55_55=0
.ic qb_55_55=1.8
.ic q_56_55=0
.ic qb_56_55=1.8
.ic q_57_55=0
.ic qb_57_55=1.8
.ic q_58_55=0
.ic qb_58_55=1.8
.ic q_59_55=0
.ic qb_59_55=1.8
.ic q_60_55=0
.ic qb_60_55=1.8
.ic q_61_55=0
.ic qb_61_55=1.8
.ic q_62_55=0
.ic qb_62_55=1.8
.ic q_63_55=0
.ic qb_63_55=1.8
.ic q_64_55=0
.ic qb_64_55=1.8
.ic q_65_55=0
.ic qb_65_55=1.8
.ic q_66_55=0
.ic qb_66_55=1.8
.ic q_67_55=0
.ic qb_67_55=1.8
.ic q_68_55=0
.ic qb_68_55=1.8
.ic q_69_55=0
.ic qb_69_55=1.8
.ic q_70_55=0
.ic qb_70_55=1.8
.ic q_71_55=0
.ic qb_71_55=1.8
.ic q_72_55=0
.ic qb_72_55=1.8
.ic q_73_55=0
.ic qb_73_55=1.8
.ic q_74_55=0
.ic qb_74_55=1.8
.ic q_75_55=0
.ic qb_75_55=1.8
.ic q_76_55=0
.ic qb_76_55=1.8
.ic q_77_55=0
.ic qb_77_55=1.8
.ic q_78_55=0
.ic qb_78_55=1.8
.ic q_79_55=0
.ic qb_79_55=1.8
.ic q_80_55=0
.ic qb_80_55=1.8
.ic q_81_55=0
.ic qb_81_55=1.8
.ic q_82_55=0
.ic qb_82_55=1.8
.ic q_83_55=0
.ic qb_83_55=1.8
.ic q_84_55=0
.ic qb_84_55=1.8
.ic q_85_55=0
.ic qb_85_55=1.8
.ic q_86_55=0
.ic qb_86_55=1.8
.ic q_87_55=0
.ic qb_87_55=1.8
.ic q_88_55=0
.ic qb_88_55=1.8
.ic q_89_55=0
.ic qb_89_55=1.8
.ic q_90_55=0
.ic qb_90_55=1.8
.ic q_91_55=0
.ic qb_91_55=1.8
.ic q_92_55=0
.ic qb_92_55=1.8
.ic q_93_55=0
.ic qb_93_55=1.8
.ic q_94_55=0
.ic qb_94_55=1.8
.ic q_95_55=0
.ic qb_95_55=1.8
.ic q_96_55=0
.ic qb_96_55=1.8
.ic q_97_55=0
.ic qb_97_55=1.8
.ic q_98_55=0
.ic qb_98_55=1.8
.ic q_99_55=0
.ic qb_99_55=1.8
.ic q_0_56=0
.ic qb_0_56=1.8
.ic q_1_56=0
.ic qb_1_56=1.8
.ic q_2_56=0
.ic qb_2_56=1.8
.ic q_3_56=0
.ic qb_3_56=1.8
.ic q_4_56=0
.ic qb_4_56=1.8
.ic q_5_56=0
.ic qb_5_56=1.8
.ic q_6_56=0
.ic qb_6_56=1.8
.ic q_7_56=0
.ic qb_7_56=1.8
.ic q_8_56=0
.ic qb_8_56=1.8
.ic q_9_56=0
.ic qb_9_56=1.8
.ic q_10_56=0
.ic qb_10_56=1.8
.ic q_11_56=0
.ic qb_11_56=1.8
.ic q_12_56=0
.ic qb_12_56=1.8
.ic q_13_56=0
.ic qb_13_56=1.8
.ic q_14_56=0
.ic qb_14_56=1.8
.ic q_15_56=0
.ic qb_15_56=1.8
.ic q_16_56=0
.ic qb_16_56=1.8
.ic q_17_56=0
.ic qb_17_56=1.8
.ic q_18_56=0
.ic qb_18_56=1.8
.ic q_19_56=0
.ic qb_19_56=1.8
.ic q_20_56=0
.ic qb_20_56=1.8
.ic q_21_56=0
.ic qb_21_56=1.8
.ic q_22_56=0
.ic qb_22_56=1.8
.ic q_23_56=0
.ic qb_23_56=1.8
.ic q_24_56=0
.ic qb_24_56=1.8
.ic q_25_56=0
.ic qb_25_56=1.8
.ic q_26_56=0
.ic qb_26_56=1.8
.ic q_27_56=0
.ic qb_27_56=1.8
.ic q_28_56=0
.ic qb_28_56=1.8
.ic q_29_56=0
.ic qb_29_56=1.8
.ic q_30_56=0
.ic qb_30_56=1.8
.ic q_31_56=0
.ic qb_31_56=1.8
.ic q_32_56=0
.ic qb_32_56=1.8
.ic q_33_56=0
.ic qb_33_56=1.8
.ic q_34_56=0
.ic qb_34_56=1.8
.ic q_35_56=0
.ic qb_35_56=1.8
.ic q_36_56=0
.ic qb_36_56=1.8
.ic q_37_56=0
.ic qb_37_56=1.8
.ic q_38_56=0
.ic qb_38_56=1.8
.ic q_39_56=0
.ic qb_39_56=1.8
.ic q_40_56=0
.ic qb_40_56=1.8
.ic q_41_56=0
.ic qb_41_56=1.8
.ic q_42_56=0
.ic qb_42_56=1.8
.ic q_43_56=0
.ic qb_43_56=1.8
.ic q_44_56=0
.ic qb_44_56=1.8
.ic q_45_56=0
.ic qb_45_56=1.8
.ic q_46_56=0
.ic qb_46_56=1.8
.ic q_47_56=0
.ic qb_47_56=1.8
.ic q_48_56=0
.ic qb_48_56=1.8
.ic q_49_56=0
.ic qb_49_56=1.8
.ic q_50_56=0
.ic qb_50_56=1.8
.ic q_51_56=0
.ic qb_51_56=1.8
.ic q_52_56=0
.ic qb_52_56=1.8
.ic q_53_56=0
.ic qb_53_56=1.8
.ic q_54_56=0
.ic qb_54_56=1.8
.ic q_55_56=0
.ic qb_55_56=1.8
.ic q_56_56=0
.ic qb_56_56=1.8
.ic q_57_56=0
.ic qb_57_56=1.8
.ic q_58_56=0
.ic qb_58_56=1.8
.ic q_59_56=0
.ic qb_59_56=1.8
.ic q_60_56=0
.ic qb_60_56=1.8
.ic q_61_56=0
.ic qb_61_56=1.8
.ic q_62_56=0
.ic qb_62_56=1.8
.ic q_63_56=0
.ic qb_63_56=1.8
.ic q_64_56=0
.ic qb_64_56=1.8
.ic q_65_56=0
.ic qb_65_56=1.8
.ic q_66_56=0
.ic qb_66_56=1.8
.ic q_67_56=0
.ic qb_67_56=1.8
.ic q_68_56=0
.ic qb_68_56=1.8
.ic q_69_56=0
.ic qb_69_56=1.8
.ic q_70_56=0
.ic qb_70_56=1.8
.ic q_71_56=0
.ic qb_71_56=1.8
.ic q_72_56=0
.ic qb_72_56=1.8
.ic q_73_56=0
.ic qb_73_56=1.8
.ic q_74_56=0
.ic qb_74_56=1.8
.ic q_75_56=0
.ic qb_75_56=1.8
.ic q_76_56=0
.ic qb_76_56=1.8
.ic q_77_56=0
.ic qb_77_56=1.8
.ic q_78_56=0
.ic qb_78_56=1.8
.ic q_79_56=0
.ic qb_79_56=1.8
.ic q_80_56=0
.ic qb_80_56=1.8
.ic q_81_56=0
.ic qb_81_56=1.8
.ic q_82_56=0
.ic qb_82_56=1.8
.ic q_83_56=0
.ic qb_83_56=1.8
.ic q_84_56=0
.ic qb_84_56=1.8
.ic q_85_56=0
.ic qb_85_56=1.8
.ic q_86_56=0
.ic qb_86_56=1.8
.ic q_87_56=0
.ic qb_87_56=1.8
.ic q_88_56=0
.ic qb_88_56=1.8
.ic q_89_56=0
.ic qb_89_56=1.8
.ic q_90_56=0
.ic qb_90_56=1.8
.ic q_91_56=0
.ic qb_91_56=1.8
.ic q_92_56=0
.ic qb_92_56=1.8
.ic q_93_56=0
.ic qb_93_56=1.8
.ic q_94_56=0
.ic qb_94_56=1.8
.ic q_95_56=0
.ic qb_95_56=1.8
.ic q_96_56=0
.ic qb_96_56=1.8
.ic q_97_56=0
.ic qb_97_56=1.8
.ic q_98_56=0
.ic qb_98_56=1.8
.ic q_99_56=0
.ic qb_99_56=1.8
.ic q_0_57=0
.ic qb_0_57=1.8
.ic q_1_57=0
.ic qb_1_57=1.8
.ic q_2_57=0
.ic qb_2_57=1.8
.ic q_3_57=0
.ic qb_3_57=1.8
.ic q_4_57=0
.ic qb_4_57=1.8
.ic q_5_57=0
.ic qb_5_57=1.8
.ic q_6_57=0
.ic qb_6_57=1.8
.ic q_7_57=0
.ic qb_7_57=1.8
.ic q_8_57=0
.ic qb_8_57=1.8
.ic q_9_57=0
.ic qb_9_57=1.8
.ic q_10_57=0
.ic qb_10_57=1.8
.ic q_11_57=0
.ic qb_11_57=1.8
.ic q_12_57=0
.ic qb_12_57=1.8
.ic q_13_57=0
.ic qb_13_57=1.8
.ic q_14_57=0
.ic qb_14_57=1.8
.ic q_15_57=0
.ic qb_15_57=1.8
.ic q_16_57=0
.ic qb_16_57=1.8
.ic q_17_57=0
.ic qb_17_57=1.8
.ic q_18_57=0
.ic qb_18_57=1.8
.ic q_19_57=0
.ic qb_19_57=1.8
.ic q_20_57=0
.ic qb_20_57=1.8
.ic q_21_57=0
.ic qb_21_57=1.8
.ic q_22_57=0
.ic qb_22_57=1.8
.ic q_23_57=0
.ic qb_23_57=1.8
.ic q_24_57=0
.ic qb_24_57=1.8
.ic q_25_57=0
.ic qb_25_57=1.8
.ic q_26_57=0
.ic qb_26_57=1.8
.ic q_27_57=0
.ic qb_27_57=1.8
.ic q_28_57=0
.ic qb_28_57=1.8
.ic q_29_57=0
.ic qb_29_57=1.8
.ic q_30_57=0
.ic qb_30_57=1.8
.ic q_31_57=0
.ic qb_31_57=1.8
.ic q_32_57=0
.ic qb_32_57=1.8
.ic q_33_57=0
.ic qb_33_57=1.8
.ic q_34_57=0
.ic qb_34_57=1.8
.ic q_35_57=0
.ic qb_35_57=1.8
.ic q_36_57=0
.ic qb_36_57=1.8
.ic q_37_57=0
.ic qb_37_57=1.8
.ic q_38_57=0
.ic qb_38_57=1.8
.ic q_39_57=0
.ic qb_39_57=1.8
.ic q_40_57=0
.ic qb_40_57=1.8
.ic q_41_57=0
.ic qb_41_57=1.8
.ic q_42_57=0
.ic qb_42_57=1.8
.ic q_43_57=0
.ic qb_43_57=1.8
.ic q_44_57=0
.ic qb_44_57=1.8
.ic q_45_57=0
.ic qb_45_57=1.8
.ic q_46_57=0
.ic qb_46_57=1.8
.ic q_47_57=0
.ic qb_47_57=1.8
.ic q_48_57=0
.ic qb_48_57=1.8
.ic q_49_57=0
.ic qb_49_57=1.8
.ic q_50_57=0
.ic qb_50_57=1.8
.ic q_51_57=0
.ic qb_51_57=1.8
.ic q_52_57=0
.ic qb_52_57=1.8
.ic q_53_57=0
.ic qb_53_57=1.8
.ic q_54_57=0
.ic qb_54_57=1.8
.ic q_55_57=0
.ic qb_55_57=1.8
.ic q_56_57=0
.ic qb_56_57=1.8
.ic q_57_57=0
.ic qb_57_57=1.8
.ic q_58_57=0
.ic qb_58_57=1.8
.ic q_59_57=0
.ic qb_59_57=1.8
.ic q_60_57=0
.ic qb_60_57=1.8
.ic q_61_57=0
.ic qb_61_57=1.8
.ic q_62_57=0
.ic qb_62_57=1.8
.ic q_63_57=0
.ic qb_63_57=1.8
.ic q_64_57=0
.ic qb_64_57=1.8
.ic q_65_57=0
.ic qb_65_57=1.8
.ic q_66_57=0
.ic qb_66_57=1.8
.ic q_67_57=0
.ic qb_67_57=1.8
.ic q_68_57=0
.ic qb_68_57=1.8
.ic q_69_57=0
.ic qb_69_57=1.8
.ic q_70_57=0
.ic qb_70_57=1.8
.ic q_71_57=0
.ic qb_71_57=1.8
.ic q_72_57=0
.ic qb_72_57=1.8
.ic q_73_57=0
.ic qb_73_57=1.8
.ic q_74_57=0
.ic qb_74_57=1.8
.ic q_75_57=0
.ic qb_75_57=1.8
.ic q_76_57=0
.ic qb_76_57=1.8
.ic q_77_57=0
.ic qb_77_57=1.8
.ic q_78_57=0
.ic qb_78_57=1.8
.ic q_79_57=0
.ic qb_79_57=1.8
.ic q_80_57=0
.ic qb_80_57=1.8
.ic q_81_57=0
.ic qb_81_57=1.8
.ic q_82_57=0
.ic qb_82_57=1.8
.ic q_83_57=0
.ic qb_83_57=1.8
.ic q_84_57=0
.ic qb_84_57=1.8
.ic q_85_57=0
.ic qb_85_57=1.8
.ic q_86_57=0
.ic qb_86_57=1.8
.ic q_87_57=0
.ic qb_87_57=1.8
.ic q_88_57=0
.ic qb_88_57=1.8
.ic q_89_57=0
.ic qb_89_57=1.8
.ic q_90_57=0
.ic qb_90_57=1.8
.ic q_91_57=0
.ic qb_91_57=1.8
.ic q_92_57=0
.ic qb_92_57=1.8
.ic q_93_57=0
.ic qb_93_57=1.8
.ic q_94_57=0
.ic qb_94_57=1.8
.ic q_95_57=0
.ic qb_95_57=1.8
.ic q_96_57=0
.ic qb_96_57=1.8
.ic q_97_57=0
.ic qb_97_57=1.8
.ic q_98_57=0
.ic qb_98_57=1.8
.ic q_99_57=0
.ic qb_99_57=1.8
.ic q_0_58=0
.ic qb_0_58=1.8
.ic q_1_58=0
.ic qb_1_58=1.8
.ic q_2_58=0
.ic qb_2_58=1.8
.ic q_3_58=0
.ic qb_3_58=1.8
.ic q_4_58=0
.ic qb_4_58=1.8
.ic q_5_58=0
.ic qb_5_58=1.8
.ic q_6_58=0
.ic qb_6_58=1.8
.ic q_7_58=0
.ic qb_7_58=1.8
.ic q_8_58=0
.ic qb_8_58=1.8
.ic q_9_58=0
.ic qb_9_58=1.8
.ic q_10_58=0
.ic qb_10_58=1.8
.ic q_11_58=0
.ic qb_11_58=1.8
.ic q_12_58=0
.ic qb_12_58=1.8
.ic q_13_58=0
.ic qb_13_58=1.8
.ic q_14_58=0
.ic qb_14_58=1.8
.ic q_15_58=0
.ic qb_15_58=1.8
.ic q_16_58=0
.ic qb_16_58=1.8
.ic q_17_58=0
.ic qb_17_58=1.8
.ic q_18_58=0
.ic qb_18_58=1.8
.ic q_19_58=0
.ic qb_19_58=1.8
.ic q_20_58=0
.ic qb_20_58=1.8
.ic q_21_58=0
.ic qb_21_58=1.8
.ic q_22_58=0
.ic qb_22_58=1.8
.ic q_23_58=0
.ic qb_23_58=1.8
.ic q_24_58=0
.ic qb_24_58=1.8
.ic q_25_58=0
.ic qb_25_58=1.8
.ic q_26_58=0
.ic qb_26_58=1.8
.ic q_27_58=0
.ic qb_27_58=1.8
.ic q_28_58=0
.ic qb_28_58=1.8
.ic q_29_58=0
.ic qb_29_58=1.8
.ic q_30_58=0
.ic qb_30_58=1.8
.ic q_31_58=0
.ic qb_31_58=1.8
.ic q_32_58=0
.ic qb_32_58=1.8
.ic q_33_58=0
.ic qb_33_58=1.8
.ic q_34_58=0
.ic qb_34_58=1.8
.ic q_35_58=0
.ic qb_35_58=1.8
.ic q_36_58=0
.ic qb_36_58=1.8
.ic q_37_58=0
.ic qb_37_58=1.8
.ic q_38_58=0
.ic qb_38_58=1.8
.ic q_39_58=0
.ic qb_39_58=1.8
.ic q_40_58=0
.ic qb_40_58=1.8
.ic q_41_58=0
.ic qb_41_58=1.8
.ic q_42_58=0
.ic qb_42_58=1.8
.ic q_43_58=0
.ic qb_43_58=1.8
.ic q_44_58=0
.ic qb_44_58=1.8
.ic q_45_58=0
.ic qb_45_58=1.8
.ic q_46_58=0
.ic qb_46_58=1.8
.ic q_47_58=0
.ic qb_47_58=1.8
.ic q_48_58=0
.ic qb_48_58=1.8
.ic q_49_58=0
.ic qb_49_58=1.8
.ic q_50_58=0
.ic qb_50_58=1.8
.ic q_51_58=0
.ic qb_51_58=1.8
.ic q_52_58=0
.ic qb_52_58=1.8
.ic q_53_58=0
.ic qb_53_58=1.8
.ic q_54_58=0
.ic qb_54_58=1.8
.ic q_55_58=0
.ic qb_55_58=1.8
.ic q_56_58=0
.ic qb_56_58=1.8
.ic q_57_58=0
.ic qb_57_58=1.8
.ic q_58_58=0
.ic qb_58_58=1.8
.ic q_59_58=0
.ic qb_59_58=1.8
.ic q_60_58=0
.ic qb_60_58=1.8
.ic q_61_58=0
.ic qb_61_58=1.8
.ic q_62_58=0
.ic qb_62_58=1.8
.ic q_63_58=0
.ic qb_63_58=1.8
.ic q_64_58=0
.ic qb_64_58=1.8
.ic q_65_58=0
.ic qb_65_58=1.8
.ic q_66_58=0
.ic qb_66_58=1.8
.ic q_67_58=0
.ic qb_67_58=1.8
.ic q_68_58=0
.ic qb_68_58=1.8
.ic q_69_58=0
.ic qb_69_58=1.8
.ic q_70_58=0
.ic qb_70_58=1.8
.ic q_71_58=0
.ic qb_71_58=1.8
.ic q_72_58=0
.ic qb_72_58=1.8
.ic q_73_58=0
.ic qb_73_58=1.8
.ic q_74_58=0
.ic qb_74_58=1.8
.ic q_75_58=0
.ic qb_75_58=1.8
.ic q_76_58=0
.ic qb_76_58=1.8
.ic q_77_58=0
.ic qb_77_58=1.8
.ic q_78_58=0
.ic qb_78_58=1.8
.ic q_79_58=0
.ic qb_79_58=1.8
.ic q_80_58=0
.ic qb_80_58=1.8
.ic q_81_58=0
.ic qb_81_58=1.8
.ic q_82_58=0
.ic qb_82_58=1.8
.ic q_83_58=0
.ic qb_83_58=1.8
.ic q_84_58=0
.ic qb_84_58=1.8
.ic q_85_58=0
.ic qb_85_58=1.8
.ic q_86_58=0
.ic qb_86_58=1.8
.ic q_87_58=0
.ic qb_87_58=1.8
.ic q_88_58=0
.ic qb_88_58=1.8
.ic q_89_58=0
.ic qb_89_58=1.8
.ic q_90_58=0
.ic qb_90_58=1.8
.ic q_91_58=0
.ic qb_91_58=1.8
.ic q_92_58=0
.ic qb_92_58=1.8
.ic q_93_58=0
.ic qb_93_58=1.8
.ic q_94_58=0
.ic qb_94_58=1.8
.ic q_95_58=0
.ic qb_95_58=1.8
.ic q_96_58=0
.ic qb_96_58=1.8
.ic q_97_58=0
.ic qb_97_58=1.8
.ic q_98_58=0
.ic qb_98_58=1.8
.ic q_99_58=0
.ic qb_99_58=1.8
.ic q_0_59=0
.ic qb_0_59=1.8
.ic q_1_59=0
.ic qb_1_59=1.8
.ic q_2_59=0
.ic qb_2_59=1.8
.ic q_3_59=0
.ic qb_3_59=1.8
.ic q_4_59=0
.ic qb_4_59=1.8
.ic q_5_59=0
.ic qb_5_59=1.8
.ic q_6_59=0
.ic qb_6_59=1.8
.ic q_7_59=0
.ic qb_7_59=1.8
.ic q_8_59=0
.ic qb_8_59=1.8
.ic q_9_59=0
.ic qb_9_59=1.8
.ic q_10_59=0
.ic qb_10_59=1.8
.ic q_11_59=0
.ic qb_11_59=1.8
.ic q_12_59=0
.ic qb_12_59=1.8
.ic q_13_59=0
.ic qb_13_59=1.8
.ic q_14_59=0
.ic qb_14_59=1.8
.ic q_15_59=0
.ic qb_15_59=1.8
.ic q_16_59=0
.ic qb_16_59=1.8
.ic q_17_59=0
.ic qb_17_59=1.8
.ic q_18_59=0
.ic qb_18_59=1.8
.ic q_19_59=0
.ic qb_19_59=1.8
.ic q_20_59=0
.ic qb_20_59=1.8
.ic q_21_59=0
.ic qb_21_59=1.8
.ic q_22_59=0
.ic qb_22_59=1.8
.ic q_23_59=0
.ic qb_23_59=1.8
.ic q_24_59=0
.ic qb_24_59=1.8
.ic q_25_59=0
.ic qb_25_59=1.8
.ic q_26_59=0
.ic qb_26_59=1.8
.ic q_27_59=0
.ic qb_27_59=1.8
.ic q_28_59=0
.ic qb_28_59=1.8
.ic q_29_59=0
.ic qb_29_59=1.8
.ic q_30_59=0
.ic qb_30_59=1.8
.ic q_31_59=0
.ic qb_31_59=1.8
.ic q_32_59=0
.ic qb_32_59=1.8
.ic q_33_59=0
.ic qb_33_59=1.8
.ic q_34_59=0
.ic qb_34_59=1.8
.ic q_35_59=0
.ic qb_35_59=1.8
.ic q_36_59=0
.ic qb_36_59=1.8
.ic q_37_59=0
.ic qb_37_59=1.8
.ic q_38_59=0
.ic qb_38_59=1.8
.ic q_39_59=0
.ic qb_39_59=1.8
.ic q_40_59=0
.ic qb_40_59=1.8
.ic q_41_59=0
.ic qb_41_59=1.8
.ic q_42_59=0
.ic qb_42_59=1.8
.ic q_43_59=0
.ic qb_43_59=1.8
.ic q_44_59=0
.ic qb_44_59=1.8
.ic q_45_59=0
.ic qb_45_59=1.8
.ic q_46_59=0
.ic qb_46_59=1.8
.ic q_47_59=0
.ic qb_47_59=1.8
.ic q_48_59=0
.ic qb_48_59=1.8
.ic q_49_59=0
.ic qb_49_59=1.8
.ic q_50_59=0
.ic qb_50_59=1.8
.ic q_51_59=0
.ic qb_51_59=1.8
.ic q_52_59=0
.ic qb_52_59=1.8
.ic q_53_59=0
.ic qb_53_59=1.8
.ic q_54_59=0
.ic qb_54_59=1.8
.ic q_55_59=0
.ic qb_55_59=1.8
.ic q_56_59=0
.ic qb_56_59=1.8
.ic q_57_59=0
.ic qb_57_59=1.8
.ic q_58_59=0
.ic qb_58_59=1.8
.ic q_59_59=0
.ic qb_59_59=1.8
.ic q_60_59=0
.ic qb_60_59=1.8
.ic q_61_59=0
.ic qb_61_59=1.8
.ic q_62_59=0
.ic qb_62_59=1.8
.ic q_63_59=0
.ic qb_63_59=1.8
.ic q_64_59=0
.ic qb_64_59=1.8
.ic q_65_59=0
.ic qb_65_59=1.8
.ic q_66_59=0
.ic qb_66_59=1.8
.ic q_67_59=0
.ic qb_67_59=1.8
.ic q_68_59=0
.ic qb_68_59=1.8
.ic q_69_59=0
.ic qb_69_59=1.8
.ic q_70_59=0
.ic qb_70_59=1.8
.ic q_71_59=0
.ic qb_71_59=1.8
.ic q_72_59=0
.ic qb_72_59=1.8
.ic q_73_59=0
.ic qb_73_59=1.8
.ic q_74_59=0
.ic qb_74_59=1.8
.ic q_75_59=0
.ic qb_75_59=1.8
.ic q_76_59=0
.ic qb_76_59=1.8
.ic q_77_59=0
.ic qb_77_59=1.8
.ic q_78_59=0
.ic qb_78_59=1.8
.ic q_79_59=0
.ic qb_79_59=1.8
.ic q_80_59=0
.ic qb_80_59=1.8
.ic q_81_59=0
.ic qb_81_59=1.8
.ic q_82_59=0
.ic qb_82_59=1.8
.ic q_83_59=0
.ic qb_83_59=1.8
.ic q_84_59=0
.ic qb_84_59=1.8
.ic q_85_59=0
.ic qb_85_59=1.8
.ic q_86_59=0
.ic qb_86_59=1.8
.ic q_87_59=0
.ic qb_87_59=1.8
.ic q_88_59=0
.ic qb_88_59=1.8
.ic q_89_59=0
.ic qb_89_59=1.8
.ic q_90_59=0
.ic qb_90_59=1.8
.ic q_91_59=0
.ic qb_91_59=1.8
.ic q_92_59=0
.ic qb_92_59=1.8
.ic q_93_59=0
.ic qb_93_59=1.8
.ic q_94_59=0
.ic qb_94_59=1.8
.ic q_95_59=0
.ic qb_95_59=1.8
.ic q_96_59=0
.ic qb_96_59=1.8
.ic q_97_59=0
.ic qb_97_59=1.8
.ic q_98_59=0
.ic qb_98_59=1.8
.ic q_99_59=0
.ic qb_99_59=1.8
.ic q_0_60=0
.ic qb_0_60=1.8
.ic q_1_60=0
.ic qb_1_60=1.8
.ic q_2_60=0
.ic qb_2_60=1.8
.ic q_3_60=0
.ic qb_3_60=1.8
.ic q_4_60=0
.ic qb_4_60=1.8
.ic q_5_60=0
.ic qb_5_60=1.8
.ic q_6_60=0
.ic qb_6_60=1.8
.ic q_7_60=0
.ic qb_7_60=1.8
.ic q_8_60=0
.ic qb_8_60=1.8
.ic q_9_60=0
.ic qb_9_60=1.8
.ic q_10_60=0
.ic qb_10_60=1.8
.ic q_11_60=0
.ic qb_11_60=1.8
.ic q_12_60=0
.ic qb_12_60=1.8
.ic q_13_60=0
.ic qb_13_60=1.8
.ic q_14_60=0
.ic qb_14_60=1.8
.ic q_15_60=0
.ic qb_15_60=1.8
.ic q_16_60=0
.ic qb_16_60=1.8
.ic q_17_60=0
.ic qb_17_60=1.8
.ic q_18_60=0
.ic qb_18_60=1.8
.ic q_19_60=0
.ic qb_19_60=1.8
.ic q_20_60=0
.ic qb_20_60=1.8
.ic q_21_60=0
.ic qb_21_60=1.8
.ic q_22_60=0
.ic qb_22_60=1.8
.ic q_23_60=0
.ic qb_23_60=1.8
.ic q_24_60=0
.ic qb_24_60=1.8
.ic q_25_60=0
.ic qb_25_60=1.8
.ic q_26_60=0
.ic qb_26_60=1.8
.ic q_27_60=0
.ic qb_27_60=1.8
.ic q_28_60=0
.ic qb_28_60=1.8
.ic q_29_60=0
.ic qb_29_60=1.8
.ic q_30_60=0
.ic qb_30_60=1.8
.ic q_31_60=0
.ic qb_31_60=1.8
.ic q_32_60=0
.ic qb_32_60=1.8
.ic q_33_60=0
.ic qb_33_60=1.8
.ic q_34_60=0
.ic qb_34_60=1.8
.ic q_35_60=0
.ic qb_35_60=1.8
.ic q_36_60=0
.ic qb_36_60=1.8
.ic q_37_60=0
.ic qb_37_60=1.8
.ic q_38_60=0
.ic qb_38_60=1.8
.ic q_39_60=0
.ic qb_39_60=1.8
.ic q_40_60=0
.ic qb_40_60=1.8
.ic q_41_60=0
.ic qb_41_60=1.8
.ic q_42_60=0
.ic qb_42_60=1.8
.ic q_43_60=0
.ic qb_43_60=1.8
.ic q_44_60=0
.ic qb_44_60=1.8
.ic q_45_60=0
.ic qb_45_60=1.8
.ic q_46_60=0
.ic qb_46_60=1.8
.ic q_47_60=0
.ic qb_47_60=1.8
.ic q_48_60=0
.ic qb_48_60=1.8
.ic q_49_60=0
.ic qb_49_60=1.8
.ic q_50_60=0
.ic qb_50_60=1.8
.ic q_51_60=0
.ic qb_51_60=1.8
.ic q_52_60=0
.ic qb_52_60=1.8
.ic q_53_60=0
.ic qb_53_60=1.8
.ic q_54_60=0
.ic qb_54_60=1.8
.ic q_55_60=0
.ic qb_55_60=1.8
.ic q_56_60=0
.ic qb_56_60=1.8
.ic q_57_60=0
.ic qb_57_60=1.8
.ic q_58_60=0
.ic qb_58_60=1.8
.ic q_59_60=0
.ic qb_59_60=1.8
.ic q_60_60=0
.ic qb_60_60=1.8
.ic q_61_60=0
.ic qb_61_60=1.8
.ic q_62_60=0
.ic qb_62_60=1.8
.ic q_63_60=0
.ic qb_63_60=1.8
.ic q_64_60=0
.ic qb_64_60=1.8
.ic q_65_60=0
.ic qb_65_60=1.8
.ic q_66_60=0
.ic qb_66_60=1.8
.ic q_67_60=0
.ic qb_67_60=1.8
.ic q_68_60=0
.ic qb_68_60=1.8
.ic q_69_60=0
.ic qb_69_60=1.8
.ic q_70_60=0
.ic qb_70_60=1.8
.ic q_71_60=0
.ic qb_71_60=1.8
.ic q_72_60=0
.ic qb_72_60=1.8
.ic q_73_60=0
.ic qb_73_60=1.8
.ic q_74_60=0
.ic qb_74_60=1.8
.ic q_75_60=0
.ic qb_75_60=1.8
.ic q_76_60=0
.ic qb_76_60=1.8
.ic q_77_60=0
.ic qb_77_60=1.8
.ic q_78_60=0
.ic qb_78_60=1.8
.ic q_79_60=0
.ic qb_79_60=1.8
.ic q_80_60=0
.ic qb_80_60=1.8
.ic q_81_60=0
.ic qb_81_60=1.8
.ic q_82_60=0
.ic qb_82_60=1.8
.ic q_83_60=0
.ic qb_83_60=1.8
.ic q_84_60=0
.ic qb_84_60=1.8
.ic q_85_60=0
.ic qb_85_60=1.8
.ic q_86_60=0
.ic qb_86_60=1.8
.ic q_87_60=0
.ic qb_87_60=1.8
.ic q_88_60=0
.ic qb_88_60=1.8
.ic q_89_60=0
.ic qb_89_60=1.8
.ic q_90_60=0
.ic qb_90_60=1.8
.ic q_91_60=0
.ic qb_91_60=1.8
.ic q_92_60=0
.ic qb_92_60=1.8
.ic q_93_60=0
.ic qb_93_60=1.8
.ic q_94_60=0
.ic qb_94_60=1.8
.ic q_95_60=0
.ic qb_95_60=1.8
.ic q_96_60=0
.ic qb_96_60=1.8
.ic q_97_60=0
.ic qb_97_60=1.8
.ic q_98_60=0
.ic qb_98_60=1.8
.ic q_99_60=0
.ic qb_99_60=1.8
.ic q_0_61=0
.ic qb_0_61=1.8
.ic q_1_61=0
.ic qb_1_61=1.8
.ic q_2_61=0
.ic qb_2_61=1.8
.ic q_3_61=0
.ic qb_3_61=1.8
.ic q_4_61=0
.ic qb_4_61=1.8
.ic q_5_61=0
.ic qb_5_61=1.8
.ic q_6_61=0
.ic qb_6_61=1.8
.ic q_7_61=0
.ic qb_7_61=1.8
.ic q_8_61=0
.ic qb_8_61=1.8
.ic q_9_61=0
.ic qb_9_61=1.8
.ic q_10_61=0
.ic qb_10_61=1.8
.ic q_11_61=0
.ic qb_11_61=1.8
.ic q_12_61=0
.ic qb_12_61=1.8
.ic q_13_61=0
.ic qb_13_61=1.8
.ic q_14_61=0
.ic qb_14_61=1.8
.ic q_15_61=0
.ic qb_15_61=1.8
.ic q_16_61=0
.ic qb_16_61=1.8
.ic q_17_61=0
.ic qb_17_61=1.8
.ic q_18_61=0
.ic qb_18_61=1.8
.ic q_19_61=0
.ic qb_19_61=1.8
.ic q_20_61=0
.ic qb_20_61=1.8
.ic q_21_61=0
.ic qb_21_61=1.8
.ic q_22_61=0
.ic qb_22_61=1.8
.ic q_23_61=0
.ic qb_23_61=1.8
.ic q_24_61=0
.ic qb_24_61=1.8
.ic q_25_61=0
.ic qb_25_61=1.8
.ic q_26_61=0
.ic qb_26_61=1.8
.ic q_27_61=0
.ic qb_27_61=1.8
.ic q_28_61=0
.ic qb_28_61=1.8
.ic q_29_61=0
.ic qb_29_61=1.8
.ic q_30_61=0
.ic qb_30_61=1.8
.ic q_31_61=0
.ic qb_31_61=1.8
.ic q_32_61=0
.ic qb_32_61=1.8
.ic q_33_61=0
.ic qb_33_61=1.8
.ic q_34_61=0
.ic qb_34_61=1.8
.ic q_35_61=0
.ic qb_35_61=1.8
.ic q_36_61=0
.ic qb_36_61=1.8
.ic q_37_61=0
.ic qb_37_61=1.8
.ic q_38_61=0
.ic qb_38_61=1.8
.ic q_39_61=0
.ic qb_39_61=1.8
.ic q_40_61=0
.ic qb_40_61=1.8
.ic q_41_61=0
.ic qb_41_61=1.8
.ic q_42_61=0
.ic qb_42_61=1.8
.ic q_43_61=0
.ic qb_43_61=1.8
.ic q_44_61=0
.ic qb_44_61=1.8
.ic q_45_61=0
.ic qb_45_61=1.8
.ic q_46_61=0
.ic qb_46_61=1.8
.ic q_47_61=0
.ic qb_47_61=1.8
.ic q_48_61=0
.ic qb_48_61=1.8
.ic q_49_61=0
.ic qb_49_61=1.8
.ic q_50_61=0
.ic qb_50_61=1.8
.ic q_51_61=0
.ic qb_51_61=1.8
.ic q_52_61=0
.ic qb_52_61=1.8
.ic q_53_61=0
.ic qb_53_61=1.8
.ic q_54_61=0
.ic qb_54_61=1.8
.ic q_55_61=0
.ic qb_55_61=1.8
.ic q_56_61=0
.ic qb_56_61=1.8
.ic q_57_61=0
.ic qb_57_61=1.8
.ic q_58_61=0
.ic qb_58_61=1.8
.ic q_59_61=0
.ic qb_59_61=1.8
.ic q_60_61=0
.ic qb_60_61=1.8
.ic q_61_61=0
.ic qb_61_61=1.8
.ic q_62_61=0
.ic qb_62_61=1.8
.ic q_63_61=0
.ic qb_63_61=1.8
.ic q_64_61=0
.ic qb_64_61=1.8
.ic q_65_61=0
.ic qb_65_61=1.8
.ic q_66_61=0
.ic qb_66_61=1.8
.ic q_67_61=0
.ic qb_67_61=1.8
.ic q_68_61=0
.ic qb_68_61=1.8
.ic q_69_61=0
.ic qb_69_61=1.8
.ic q_70_61=0
.ic qb_70_61=1.8
.ic q_71_61=0
.ic qb_71_61=1.8
.ic q_72_61=0
.ic qb_72_61=1.8
.ic q_73_61=0
.ic qb_73_61=1.8
.ic q_74_61=0
.ic qb_74_61=1.8
.ic q_75_61=0
.ic qb_75_61=1.8
.ic q_76_61=0
.ic qb_76_61=1.8
.ic q_77_61=0
.ic qb_77_61=1.8
.ic q_78_61=0
.ic qb_78_61=1.8
.ic q_79_61=0
.ic qb_79_61=1.8
.ic q_80_61=0
.ic qb_80_61=1.8
.ic q_81_61=0
.ic qb_81_61=1.8
.ic q_82_61=0
.ic qb_82_61=1.8
.ic q_83_61=0
.ic qb_83_61=1.8
.ic q_84_61=0
.ic qb_84_61=1.8
.ic q_85_61=0
.ic qb_85_61=1.8
.ic q_86_61=0
.ic qb_86_61=1.8
.ic q_87_61=0
.ic qb_87_61=1.8
.ic q_88_61=0
.ic qb_88_61=1.8
.ic q_89_61=0
.ic qb_89_61=1.8
.ic q_90_61=0
.ic qb_90_61=1.8
.ic q_91_61=0
.ic qb_91_61=1.8
.ic q_92_61=0
.ic qb_92_61=1.8
.ic q_93_61=0
.ic qb_93_61=1.8
.ic q_94_61=0
.ic qb_94_61=1.8
.ic q_95_61=0
.ic qb_95_61=1.8
.ic q_96_61=0
.ic qb_96_61=1.8
.ic q_97_61=0
.ic qb_97_61=1.8
.ic q_98_61=0
.ic qb_98_61=1.8
.ic q_99_61=0
.ic qb_99_61=1.8
.ic q_0_62=0
.ic qb_0_62=1.8
.ic q_1_62=0
.ic qb_1_62=1.8
.ic q_2_62=0
.ic qb_2_62=1.8
.ic q_3_62=0
.ic qb_3_62=1.8
.ic q_4_62=0
.ic qb_4_62=1.8
.ic q_5_62=0
.ic qb_5_62=1.8
.ic q_6_62=0
.ic qb_6_62=1.8
.ic q_7_62=0
.ic qb_7_62=1.8
.ic q_8_62=0
.ic qb_8_62=1.8
.ic q_9_62=0
.ic qb_9_62=1.8
.ic q_10_62=0
.ic qb_10_62=1.8
.ic q_11_62=0
.ic qb_11_62=1.8
.ic q_12_62=0
.ic qb_12_62=1.8
.ic q_13_62=0
.ic qb_13_62=1.8
.ic q_14_62=0
.ic qb_14_62=1.8
.ic q_15_62=0
.ic qb_15_62=1.8
.ic q_16_62=0
.ic qb_16_62=1.8
.ic q_17_62=0
.ic qb_17_62=1.8
.ic q_18_62=0
.ic qb_18_62=1.8
.ic q_19_62=0
.ic qb_19_62=1.8
.ic q_20_62=0
.ic qb_20_62=1.8
.ic q_21_62=0
.ic qb_21_62=1.8
.ic q_22_62=0
.ic qb_22_62=1.8
.ic q_23_62=0
.ic qb_23_62=1.8
.ic q_24_62=0
.ic qb_24_62=1.8
.ic q_25_62=0
.ic qb_25_62=1.8
.ic q_26_62=0
.ic qb_26_62=1.8
.ic q_27_62=0
.ic qb_27_62=1.8
.ic q_28_62=0
.ic qb_28_62=1.8
.ic q_29_62=0
.ic qb_29_62=1.8
.ic q_30_62=0
.ic qb_30_62=1.8
.ic q_31_62=0
.ic qb_31_62=1.8
.ic q_32_62=0
.ic qb_32_62=1.8
.ic q_33_62=0
.ic qb_33_62=1.8
.ic q_34_62=0
.ic qb_34_62=1.8
.ic q_35_62=0
.ic qb_35_62=1.8
.ic q_36_62=0
.ic qb_36_62=1.8
.ic q_37_62=0
.ic qb_37_62=1.8
.ic q_38_62=0
.ic qb_38_62=1.8
.ic q_39_62=0
.ic qb_39_62=1.8
.ic q_40_62=0
.ic qb_40_62=1.8
.ic q_41_62=0
.ic qb_41_62=1.8
.ic q_42_62=0
.ic qb_42_62=1.8
.ic q_43_62=0
.ic qb_43_62=1.8
.ic q_44_62=0
.ic qb_44_62=1.8
.ic q_45_62=0
.ic qb_45_62=1.8
.ic q_46_62=0
.ic qb_46_62=1.8
.ic q_47_62=0
.ic qb_47_62=1.8
.ic q_48_62=0
.ic qb_48_62=1.8
.ic q_49_62=0
.ic qb_49_62=1.8
.ic q_50_62=0
.ic qb_50_62=1.8
.ic q_51_62=0
.ic qb_51_62=1.8
.ic q_52_62=0
.ic qb_52_62=1.8
.ic q_53_62=0
.ic qb_53_62=1.8
.ic q_54_62=0
.ic qb_54_62=1.8
.ic q_55_62=0
.ic qb_55_62=1.8
.ic q_56_62=0
.ic qb_56_62=1.8
.ic q_57_62=0
.ic qb_57_62=1.8
.ic q_58_62=0
.ic qb_58_62=1.8
.ic q_59_62=0
.ic qb_59_62=1.8
.ic q_60_62=0
.ic qb_60_62=1.8
.ic q_61_62=0
.ic qb_61_62=1.8
.ic q_62_62=0
.ic qb_62_62=1.8
.ic q_63_62=0
.ic qb_63_62=1.8
.ic q_64_62=0
.ic qb_64_62=1.8
.ic q_65_62=0
.ic qb_65_62=1.8
.ic q_66_62=0
.ic qb_66_62=1.8
.ic q_67_62=0
.ic qb_67_62=1.8
.ic q_68_62=0
.ic qb_68_62=1.8
.ic q_69_62=0
.ic qb_69_62=1.8
.ic q_70_62=0
.ic qb_70_62=1.8
.ic q_71_62=0
.ic qb_71_62=1.8
.ic q_72_62=0
.ic qb_72_62=1.8
.ic q_73_62=0
.ic qb_73_62=1.8
.ic q_74_62=0
.ic qb_74_62=1.8
.ic q_75_62=0
.ic qb_75_62=1.8
.ic q_76_62=0
.ic qb_76_62=1.8
.ic q_77_62=0
.ic qb_77_62=1.8
.ic q_78_62=0
.ic qb_78_62=1.8
.ic q_79_62=0
.ic qb_79_62=1.8
.ic q_80_62=0
.ic qb_80_62=1.8
.ic q_81_62=0
.ic qb_81_62=1.8
.ic q_82_62=0
.ic qb_82_62=1.8
.ic q_83_62=0
.ic qb_83_62=1.8
.ic q_84_62=0
.ic qb_84_62=1.8
.ic q_85_62=0
.ic qb_85_62=1.8
.ic q_86_62=0
.ic qb_86_62=1.8
.ic q_87_62=0
.ic qb_87_62=1.8
.ic q_88_62=0
.ic qb_88_62=1.8
.ic q_89_62=0
.ic qb_89_62=1.8
.ic q_90_62=0
.ic qb_90_62=1.8
.ic q_91_62=0
.ic qb_91_62=1.8
.ic q_92_62=0
.ic qb_92_62=1.8
.ic q_93_62=0
.ic qb_93_62=1.8
.ic q_94_62=0
.ic qb_94_62=1.8
.ic q_95_62=0
.ic qb_95_62=1.8
.ic q_96_62=0
.ic qb_96_62=1.8
.ic q_97_62=0
.ic qb_97_62=1.8
.ic q_98_62=0
.ic qb_98_62=1.8
.ic q_99_62=0
.ic qb_99_62=1.8
.ic q_0_63=0
.ic qb_0_63=1.8
.ic q_1_63=0
.ic qb_1_63=1.8
.ic q_2_63=0
.ic qb_2_63=1.8
.ic q_3_63=0
.ic qb_3_63=1.8
.ic q_4_63=0
.ic qb_4_63=1.8
.ic q_5_63=0
.ic qb_5_63=1.8
.ic q_6_63=0
.ic qb_6_63=1.8
.ic q_7_63=0
.ic qb_7_63=1.8
.ic q_8_63=0
.ic qb_8_63=1.8
.ic q_9_63=0
.ic qb_9_63=1.8
.ic q_10_63=0
.ic qb_10_63=1.8
.ic q_11_63=0
.ic qb_11_63=1.8
.ic q_12_63=0
.ic qb_12_63=1.8
.ic q_13_63=0
.ic qb_13_63=1.8
.ic q_14_63=0
.ic qb_14_63=1.8
.ic q_15_63=0
.ic qb_15_63=1.8
.ic q_16_63=0
.ic qb_16_63=1.8
.ic q_17_63=0
.ic qb_17_63=1.8
.ic q_18_63=0
.ic qb_18_63=1.8
.ic q_19_63=0
.ic qb_19_63=1.8
.ic q_20_63=0
.ic qb_20_63=1.8
.ic q_21_63=0
.ic qb_21_63=1.8
.ic q_22_63=0
.ic qb_22_63=1.8
.ic q_23_63=0
.ic qb_23_63=1.8
.ic q_24_63=0
.ic qb_24_63=1.8
.ic q_25_63=0
.ic qb_25_63=1.8
.ic q_26_63=0
.ic qb_26_63=1.8
.ic q_27_63=0
.ic qb_27_63=1.8
.ic q_28_63=0
.ic qb_28_63=1.8
.ic q_29_63=0
.ic qb_29_63=1.8
.ic q_30_63=0
.ic qb_30_63=1.8
.ic q_31_63=0
.ic qb_31_63=1.8
.ic q_32_63=0
.ic qb_32_63=1.8
.ic q_33_63=0
.ic qb_33_63=1.8
.ic q_34_63=0
.ic qb_34_63=1.8
.ic q_35_63=0
.ic qb_35_63=1.8
.ic q_36_63=0
.ic qb_36_63=1.8
.ic q_37_63=0
.ic qb_37_63=1.8
.ic q_38_63=0
.ic qb_38_63=1.8
.ic q_39_63=0
.ic qb_39_63=1.8
.ic q_40_63=0
.ic qb_40_63=1.8
.ic q_41_63=0
.ic qb_41_63=1.8
.ic q_42_63=0
.ic qb_42_63=1.8
.ic q_43_63=0
.ic qb_43_63=1.8
.ic q_44_63=0
.ic qb_44_63=1.8
.ic q_45_63=0
.ic qb_45_63=1.8
.ic q_46_63=0
.ic qb_46_63=1.8
.ic q_47_63=0
.ic qb_47_63=1.8
.ic q_48_63=0
.ic qb_48_63=1.8
.ic q_49_63=0
.ic qb_49_63=1.8
.ic q_50_63=0
.ic qb_50_63=1.8
.ic q_51_63=0
.ic qb_51_63=1.8
.ic q_52_63=0
.ic qb_52_63=1.8
.ic q_53_63=0
.ic qb_53_63=1.8
.ic q_54_63=0
.ic qb_54_63=1.8
.ic q_55_63=0
.ic qb_55_63=1.8
.ic q_56_63=0
.ic qb_56_63=1.8
.ic q_57_63=0
.ic qb_57_63=1.8
.ic q_58_63=0
.ic qb_58_63=1.8
.ic q_59_63=0
.ic qb_59_63=1.8
.ic q_60_63=0
.ic qb_60_63=1.8
.ic q_61_63=0
.ic qb_61_63=1.8
.ic q_62_63=0
.ic qb_62_63=1.8
.ic q_63_63=0
.ic qb_63_63=1.8
.ic q_64_63=0
.ic qb_64_63=1.8
.ic q_65_63=0
.ic qb_65_63=1.8
.ic q_66_63=0
.ic qb_66_63=1.8
.ic q_67_63=0
.ic qb_67_63=1.8
.ic q_68_63=0
.ic qb_68_63=1.8
.ic q_69_63=0
.ic qb_69_63=1.8
.ic q_70_63=0
.ic qb_70_63=1.8
.ic q_71_63=0
.ic qb_71_63=1.8
.ic q_72_63=0
.ic qb_72_63=1.8
.ic q_73_63=0
.ic qb_73_63=1.8
.ic q_74_63=0
.ic qb_74_63=1.8
.ic q_75_63=0
.ic qb_75_63=1.8
.ic q_76_63=0
.ic qb_76_63=1.8
.ic q_77_63=0
.ic qb_77_63=1.8
.ic q_78_63=0
.ic qb_78_63=1.8
.ic q_79_63=0
.ic qb_79_63=1.8
.ic q_80_63=0
.ic qb_80_63=1.8
.ic q_81_63=0
.ic qb_81_63=1.8
.ic q_82_63=0
.ic qb_82_63=1.8
.ic q_83_63=0
.ic qb_83_63=1.8
.ic q_84_63=0
.ic qb_84_63=1.8
.ic q_85_63=0
.ic qb_85_63=1.8
.ic q_86_63=0
.ic qb_86_63=1.8
.ic q_87_63=0
.ic qb_87_63=1.8
.ic q_88_63=0
.ic qb_88_63=1.8
.ic q_89_63=0
.ic qb_89_63=1.8
.ic q_90_63=0
.ic qb_90_63=1.8
.ic q_91_63=0
.ic qb_91_63=1.8
.ic q_92_63=0
.ic qb_92_63=1.8
.ic q_93_63=0
.ic qb_93_63=1.8
.ic q_94_63=0
.ic qb_94_63=1.8
.ic q_95_63=0
.ic qb_95_63=1.8
.ic q_96_63=0
.ic qb_96_63=1.8
.ic q_97_63=0
.ic qb_97_63=1.8
.ic q_98_63=0
.ic qb_98_63=1.8
.ic q_99_63=0
.ic qb_99_63=1.8
.ic q_0_64=0
.ic qb_0_64=1.8
.ic q_1_64=0
.ic qb_1_64=1.8
.ic q_2_64=0
.ic qb_2_64=1.8
.ic q_3_64=0
.ic qb_3_64=1.8
.ic q_4_64=0
.ic qb_4_64=1.8
.ic q_5_64=0
.ic qb_5_64=1.8
.ic q_6_64=0
.ic qb_6_64=1.8
.ic q_7_64=0
.ic qb_7_64=1.8
.ic q_8_64=0
.ic qb_8_64=1.8
.ic q_9_64=0
.ic qb_9_64=1.8
.ic q_10_64=0
.ic qb_10_64=1.8
.ic q_11_64=0
.ic qb_11_64=1.8
.ic q_12_64=0
.ic qb_12_64=1.8
.ic q_13_64=0
.ic qb_13_64=1.8
.ic q_14_64=0
.ic qb_14_64=1.8
.ic q_15_64=0
.ic qb_15_64=1.8
.ic q_16_64=0
.ic qb_16_64=1.8
.ic q_17_64=0
.ic qb_17_64=1.8
.ic q_18_64=0
.ic qb_18_64=1.8
.ic q_19_64=0
.ic qb_19_64=1.8
.ic q_20_64=0
.ic qb_20_64=1.8
.ic q_21_64=0
.ic qb_21_64=1.8
.ic q_22_64=0
.ic qb_22_64=1.8
.ic q_23_64=0
.ic qb_23_64=1.8
.ic q_24_64=0
.ic qb_24_64=1.8
.ic q_25_64=0
.ic qb_25_64=1.8
.ic q_26_64=0
.ic qb_26_64=1.8
.ic q_27_64=0
.ic qb_27_64=1.8
.ic q_28_64=0
.ic qb_28_64=1.8
.ic q_29_64=0
.ic qb_29_64=1.8
.ic q_30_64=0
.ic qb_30_64=1.8
.ic q_31_64=0
.ic qb_31_64=1.8
.ic q_32_64=0
.ic qb_32_64=1.8
.ic q_33_64=0
.ic qb_33_64=1.8
.ic q_34_64=0
.ic qb_34_64=1.8
.ic q_35_64=0
.ic qb_35_64=1.8
.ic q_36_64=0
.ic qb_36_64=1.8
.ic q_37_64=0
.ic qb_37_64=1.8
.ic q_38_64=0
.ic qb_38_64=1.8
.ic q_39_64=0
.ic qb_39_64=1.8
.ic q_40_64=0
.ic qb_40_64=1.8
.ic q_41_64=0
.ic qb_41_64=1.8
.ic q_42_64=0
.ic qb_42_64=1.8
.ic q_43_64=0
.ic qb_43_64=1.8
.ic q_44_64=0
.ic qb_44_64=1.8
.ic q_45_64=0
.ic qb_45_64=1.8
.ic q_46_64=0
.ic qb_46_64=1.8
.ic q_47_64=0
.ic qb_47_64=1.8
.ic q_48_64=0
.ic qb_48_64=1.8
.ic q_49_64=0
.ic qb_49_64=1.8
.ic q_50_64=0
.ic qb_50_64=1.8
.ic q_51_64=0
.ic qb_51_64=1.8
.ic q_52_64=0
.ic qb_52_64=1.8
.ic q_53_64=0
.ic qb_53_64=1.8
.ic q_54_64=0
.ic qb_54_64=1.8
.ic q_55_64=0
.ic qb_55_64=1.8
.ic q_56_64=0
.ic qb_56_64=1.8
.ic q_57_64=0
.ic qb_57_64=1.8
.ic q_58_64=0
.ic qb_58_64=1.8
.ic q_59_64=0
.ic qb_59_64=1.8
.ic q_60_64=0
.ic qb_60_64=1.8
.ic q_61_64=0
.ic qb_61_64=1.8
.ic q_62_64=0
.ic qb_62_64=1.8
.ic q_63_64=0
.ic qb_63_64=1.8
.ic q_64_64=0
.ic qb_64_64=1.8
.ic q_65_64=0
.ic qb_65_64=1.8
.ic q_66_64=0
.ic qb_66_64=1.8
.ic q_67_64=0
.ic qb_67_64=1.8
.ic q_68_64=0
.ic qb_68_64=1.8
.ic q_69_64=0
.ic qb_69_64=1.8
.ic q_70_64=0
.ic qb_70_64=1.8
.ic q_71_64=0
.ic qb_71_64=1.8
.ic q_72_64=0
.ic qb_72_64=1.8
.ic q_73_64=0
.ic qb_73_64=1.8
.ic q_74_64=0
.ic qb_74_64=1.8
.ic q_75_64=0
.ic qb_75_64=1.8
.ic q_76_64=0
.ic qb_76_64=1.8
.ic q_77_64=0
.ic qb_77_64=1.8
.ic q_78_64=0
.ic qb_78_64=1.8
.ic q_79_64=0
.ic qb_79_64=1.8
.ic q_80_64=0
.ic qb_80_64=1.8
.ic q_81_64=0
.ic qb_81_64=1.8
.ic q_82_64=0
.ic qb_82_64=1.8
.ic q_83_64=0
.ic qb_83_64=1.8
.ic q_84_64=0
.ic qb_84_64=1.8
.ic q_85_64=0
.ic qb_85_64=1.8
.ic q_86_64=0
.ic qb_86_64=1.8
.ic q_87_64=0
.ic qb_87_64=1.8
.ic q_88_64=0
.ic qb_88_64=1.8
.ic q_89_64=0
.ic qb_89_64=1.8
.ic q_90_64=0
.ic qb_90_64=1.8
.ic q_91_64=0
.ic qb_91_64=1.8
.ic q_92_64=0
.ic qb_92_64=1.8
.ic q_93_64=0
.ic qb_93_64=1.8
.ic q_94_64=0
.ic qb_94_64=1.8
.ic q_95_64=0
.ic qb_95_64=1.8
.ic q_96_64=0
.ic qb_96_64=1.8
.ic q_97_64=0
.ic qb_97_64=1.8
.ic q_98_64=0
.ic qb_98_64=1.8
.ic q_99_64=0
.ic qb_99_64=1.8
.ic q_0_65=0
.ic qb_0_65=1.8
.ic q_1_65=0
.ic qb_1_65=1.8
.ic q_2_65=0
.ic qb_2_65=1.8
.ic q_3_65=0
.ic qb_3_65=1.8
.ic q_4_65=0
.ic qb_4_65=1.8
.ic q_5_65=0
.ic qb_5_65=1.8
.ic q_6_65=0
.ic qb_6_65=1.8
.ic q_7_65=0
.ic qb_7_65=1.8
.ic q_8_65=0
.ic qb_8_65=1.8
.ic q_9_65=0
.ic qb_9_65=1.8
.ic q_10_65=0
.ic qb_10_65=1.8
.ic q_11_65=0
.ic qb_11_65=1.8
.ic q_12_65=0
.ic qb_12_65=1.8
.ic q_13_65=0
.ic qb_13_65=1.8
.ic q_14_65=0
.ic qb_14_65=1.8
.ic q_15_65=0
.ic qb_15_65=1.8
.ic q_16_65=0
.ic qb_16_65=1.8
.ic q_17_65=0
.ic qb_17_65=1.8
.ic q_18_65=0
.ic qb_18_65=1.8
.ic q_19_65=0
.ic qb_19_65=1.8
.ic q_20_65=0
.ic qb_20_65=1.8
.ic q_21_65=0
.ic qb_21_65=1.8
.ic q_22_65=0
.ic qb_22_65=1.8
.ic q_23_65=0
.ic qb_23_65=1.8
.ic q_24_65=0
.ic qb_24_65=1.8
.ic q_25_65=0
.ic qb_25_65=1.8
.ic q_26_65=0
.ic qb_26_65=1.8
.ic q_27_65=0
.ic qb_27_65=1.8
.ic q_28_65=0
.ic qb_28_65=1.8
.ic q_29_65=0
.ic qb_29_65=1.8
.ic q_30_65=0
.ic qb_30_65=1.8
.ic q_31_65=0
.ic qb_31_65=1.8
.ic q_32_65=0
.ic qb_32_65=1.8
.ic q_33_65=0
.ic qb_33_65=1.8
.ic q_34_65=0
.ic qb_34_65=1.8
.ic q_35_65=0
.ic qb_35_65=1.8
.ic q_36_65=0
.ic qb_36_65=1.8
.ic q_37_65=0
.ic qb_37_65=1.8
.ic q_38_65=0
.ic qb_38_65=1.8
.ic q_39_65=0
.ic qb_39_65=1.8
.ic q_40_65=0
.ic qb_40_65=1.8
.ic q_41_65=0
.ic qb_41_65=1.8
.ic q_42_65=0
.ic qb_42_65=1.8
.ic q_43_65=0
.ic qb_43_65=1.8
.ic q_44_65=0
.ic qb_44_65=1.8
.ic q_45_65=0
.ic qb_45_65=1.8
.ic q_46_65=0
.ic qb_46_65=1.8
.ic q_47_65=0
.ic qb_47_65=1.8
.ic q_48_65=0
.ic qb_48_65=1.8
.ic q_49_65=0
.ic qb_49_65=1.8
.ic q_50_65=0
.ic qb_50_65=1.8
.ic q_51_65=0
.ic qb_51_65=1.8
.ic q_52_65=0
.ic qb_52_65=1.8
.ic q_53_65=0
.ic qb_53_65=1.8
.ic q_54_65=0
.ic qb_54_65=1.8
.ic q_55_65=0
.ic qb_55_65=1.8
.ic q_56_65=0
.ic qb_56_65=1.8
.ic q_57_65=0
.ic qb_57_65=1.8
.ic q_58_65=0
.ic qb_58_65=1.8
.ic q_59_65=0
.ic qb_59_65=1.8
.ic q_60_65=0
.ic qb_60_65=1.8
.ic q_61_65=0
.ic qb_61_65=1.8
.ic q_62_65=0
.ic qb_62_65=1.8
.ic q_63_65=0
.ic qb_63_65=1.8
.ic q_64_65=0
.ic qb_64_65=1.8
.ic q_65_65=0
.ic qb_65_65=1.8
.ic q_66_65=0
.ic qb_66_65=1.8
.ic q_67_65=0
.ic qb_67_65=1.8
.ic q_68_65=0
.ic qb_68_65=1.8
.ic q_69_65=0
.ic qb_69_65=1.8
.ic q_70_65=0
.ic qb_70_65=1.8
.ic q_71_65=0
.ic qb_71_65=1.8
.ic q_72_65=0
.ic qb_72_65=1.8
.ic q_73_65=0
.ic qb_73_65=1.8
.ic q_74_65=0
.ic qb_74_65=1.8
.ic q_75_65=0
.ic qb_75_65=1.8
.ic q_76_65=0
.ic qb_76_65=1.8
.ic q_77_65=0
.ic qb_77_65=1.8
.ic q_78_65=0
.ic qb_78_65=1.8
.ic q_79_65=0
.ic qb_79_65=1.8
.ic q_80_65=0
.ic qb_80_65=1.8
.ic q_81_65=0
.ic qb_81_65=1.8
.ic q_82_65=0
.ic qb_82_65=1.8
.ic q_83_65=0
.ic qb_83_65=1.8
.ic q_84_65=0
.ic qb_84_65=1.8
.ic q_85_65=0
.ic qb_85_65=1.8
.ic q_86_65=0
.ic qb_86_65=1.8
.ic q_87_65=0
.ic qb_87_65=1.8
.ic q_88_65=0
.ic qb_88_65=1.8
.ic q_89_65=0
.ic qb_89_65=1.8
.ic q_90_65=0
.ic qb_90_65=1.8
.ic q_91_65=0
.ic qb_91_65=1.8
.ic q_92_65=0
.ic qb_92_65=1.8
.ic q_93_65=0
.ic qb_93_65=1.8
.ic q_94_65=0
.ic qb_94_65=1.8
.ic q_95_65=0
.ic qb_95_65=1.8
.ic q_96_65=0
.ic qb_96_65=1.8
.ic q_97_65=0
.ic qb_97_65=1.8
.ic q_98_65=0
.ic qb_98_65=1.8
.ic q_99_65=0
.ic qb_99_65=1.8
.ic q_0_66=0
.ic qb_0_66=1.8
.ic q_1_66=0
.ic qb_1_66=1.8
.ic q_2_66=0
.ic qb_2_66=1.8
.ic q_3_66=0
.ic qb_3_66=1.8
.ic q_4_66=0
.ic qb_4_66=1.8
.ic q_5_66=0
.ic qb_5_66=1.8
.ic q_6_66=0
.ic qb_6_66=1.8
.ic q_7_66=0
.ic qb_7_66=1.8
.ic q_8_66=0
.ic qb_8_66=1.8
.ic q_9_66=0
.ic qb_9_66=1.8
.ic q_10_66=0
.ic qb_10_66=1.8
.ic q_11_66=0
.ic qb_11_66=1.8
.ic q_12_66=0
.ic qb_12_66=1.8
.ic q_13_66=0
.ic qb_13_66=1.8
.ic q_14_66=0
.ic qb_14_66=1.8
.ic q_15_66=0
.ic qb_15_66=1.8
.ic q_16_66=0
.ic qb_16_66=1.8
.ic q_17_66=0
.ic qb_17_66=1.8
.ic q_18_66=0
.ic qb_18_66=1.8
.ic q_19_66=0
.ic qb_19_66=1.8
.ic q_20_66=0
.ic qb_20_66=1.8
.ic q_21_66=0
.ic qb_21_66=1.8
.ic q_22_66=0
.ic qb_22_66=1.8
.ic q_23_66=0
.ic qb_23_66=1.8
.ic q_24_66=0
.ic qb_24_66=1.8
.ic q_25_66=0
.ic qb_25_66=1.8
.ic q_26_66=0
.ic qb_26_66=1.8
.ic q_27_66=0
.ic qb_27_66=1.8
.ic q_28_66=0
.ic qb_28_66=1.8
.ic q_29_66=0
.ic qb_29_66=1.8
.ic q_30_66=0
.ic qb_30_66=1.8
.ic q_31_66=0
.ic qb_31_66=1.8
.ic q_32_66=0
.ic qb_32_66=1.8
.ic q_33_66=0
.ic qb_33_66=1.8
.ic q_34_66=0
.ic qb_34_66=1.8
.ic q_35_66=0
.ic qb_35_66=1.8
.ic q_36_66=0
.ic qb_36_66=1.8
.ic q_37_66=0
.ic qb_37_66=1.8
.ic q_38_66=0
.ic qb_38_66=1.8
.ic q_39_66=0
.ic qb_39_66=1.8
.ic q_40_66=0
.ic qb_40_66=1.8
.ic q_41_66=0
.ic qb_41_66=1.8
.ic q_42_66=0
.ic qb_42_66=1.8
.ic q_43_66=0
.ic qb_43_66=1.8
.ic q_44_66=0
.ic qb_44_66=1.8
.ic q_45_66=0
.ic qb_45_66=1.8
.ic q_46_66=0
.ic qb_46_66=1.8
.ic q_47_66=0
.ic qb_47_66=1.8
.ic q_48_66=0
.ic qb_48_66=1.8
.ic q_49_66=0
.ic qb_49_66=1.8
.ic q_50_66=0
.ic qb_50_66=1.8
.ic q_51_66=0
.ic qb_51_66=1.8
.ic q_52_66=0
.ic qb_52_66=1.8
.ic q_53_66=0
.ic qb_53_66=1.8
.ic q_54_66=0
.ic qb_54_66=1.8
.ic q_55_66=0
.ic qb_55_66=1.8
.ic q_56_66=0
.ic qb_56_66=1.8
.ic q_57_66=0
.ic qb_57_66=1.8
.ic q_58_66=0
.ic qb_58_66=1.8
.ic q_59_66=0
.ic qb_59_66=1.8
.ic q_60_66=0
.ic qb_60_66=1.8
.ic q_61_66=0
.ic qb_61_66=1.8
.ic q_62_66=0
.ic qb_62_66=1.8
.ic q_63_66=0
.ic qb_63_66=1.8
.ic q_64_66=0
.ic qb_64_66=1.8
.ic q_65_66=0
.ic qb_65_66=1.8
.ic q_66_66=0
.ic qb_66_66=1.8
.ic q_67_66=0
.ic qb_67_66=1.8
.ic q_68_66=0
.ic qb_68_66=1.8
.ic q_69_66=0
.ic qb_69_66=1.8
.ic q_70_66=0
.ic qb_70_66=1.8
.ic q_71_66=0
.ic qb_71_66=1.8
.ic q_72_66=0
.ic qb_72_66=1.8
.ic q_73_66=0
.ic qb_73_66=1.8
.ic q_74_66=0
.ic qb_74_66=1.8
.ic q_75_66=0
.ic qb_75_66=1.8
.ic q_76_66=0
.ic qb_76_66=1.8
.ic q_77_66=0
.ic qb_77_66=1.8
.ic q_78_66=0
.ic qb_78_66=1.8
.ic q_79_66=0
.ic qb_79_66=1.8
.ic q_80_66=0
.ic qb_80_66=1.8
.ic q_81_66=0
.ic qb_81_66=1.8
.ic q_82_66=0
.ic qb_82_66=1.8
.ic q_83_66=0
.ic qb_83_66=1.8
.ic q_84_66=0
.ic qb_84_66=1.8
.ic q_85_66=0
.ic qb_85_66=1.8
.ic q_86_66=0
.ic qb_86_66=1.8
.ic q_87_66=0
.ic qb_87_66=1.8
.ic q_88_66=0
.ic qb_88_66=1.8
.ic q_89_66=0
.ic qb_89_66=1.8
.ic q_90_66=0
.ic qb_90_66=1.8
.ic q_91_66=0
.ic qb_91_66=1.8
.ic q_92_66=0
.ic qb_92_66=1.8
.ic q_93_66=0
.ic qb_93_66=1.8
.ic q_94_66=0
.ic qb_94_66=1.8
.ic q_95_66=0
.ic qb_95_66=1.8
.ic q_96_66=0
.ic qb_96_66=1.8
.ic q_97_66=0
.ic qb_97_66=1.8
.ic q_98_66=0
.ic qb_98_66=1.8
.ic q_99_66=0
.ic qb_99_66=1.8
.ic q_0_67=0
.ic qb_0_67=1.8
.ic q_1_67=0
.ic qb_1_67=1.8
.ic q_2_67=0
.ic qb_2_67=1.8
.ic q_3_67=0
.ic qb_3_67=1.8
.ic q_4_67=0
.ic qb_4_67=1.8
.ic q_5_67=0
.ic qb_5_67=1.8
.ic q_6_67=0
.ic qb_6_67=1.8
.ic q_7_67=0
.ic qb_7_67=1.8
.ic q_8_67=0
.ic qb_8_67=1.8
.ic q_9_67=0
.ic qb_9_67=1.8
.ic q_10_67=0
.ic qb_10_67=1.8
.ic q_11_67=0
.ic qb_11_67=1.8
.ic q_12_67=0
.ic qb_12_67=1.8
.ic q_13_67=0
.ic qb_13_67=1.8
.ic q_14_67=0
.ic qb_14_67=1.8
.ic q_15_67=0
.ic qb_15_67=1.8
.ic q_16_67=0
.ic qb_16_67=1.8
.ic q_17_67=0
.ic qb_17_67=1.8
.ic q_18_67=0
.ic qb_18_67=1.8
.ic q_19_67=0
.ic qb_19_67=1.8
.ic q_20_67=0
.ic qb_20_67=1.8
.ic q_21_67=0
.ic qb_21_67=1.8
.ic q_22_67=0
.ic qb_22_67=1.8
.ic q_23_67=0
.ic qb_23_67=1.8
.ic q_24_67=0
.ic qb_24_67=1.8
.ic q_25_67=0
.ic qb_25_67=1.8
.ic q_26_67=0
.ic qb_26_67=1.8
.ic q_27_67=0
.ic qb_27_67=1.8
.ic q_28_67=0
.ic qb_28_67=1.8
.ic q_29_67=0
.ic qb_29_67=1.8
.ic q_30_67=0
.ic qb_30_67=1.8
.ic q_31_67=0
.ic qb_31_67=1.8
.ic q_32_67=0
.ic qb_32_67=1.8
.ic q_33_67=0
.ic qb_33_67=1.8
.ic q_34_67=0
.ic qb_34_67=1.8
.ic q_35_67=0
.ic qb_35_67=1.8
.ic q_36_67=0
.ic qb_36_67=1.8
.ic q_37_67=0
.ic qb_37_67=1.8
.ic q_38_67=0
.ic qb_38_67=1.8
.ic q_39_67=0
.ic qb_39_67=1.8
.ic q_40_67=0
.ic qb_40_67=1.8
.ic q_41_67=0
.ic qb_41_67=1.8
.ic q_42_67=0
.ic qb_42_67=1.8
.ic q_43_67=0
.ic qb_43_67=1.8
.ic q_44_67=0
.ic qb_44_67=1.8
.ic q_45_67=0
.ic qb_45_67=1.8
.ic q_46_67=0
.ic qb_46_67=1.8
.ic q_47_67=0
.ic qb_47_67=1.8
.ic q_48_67=0
.ic qb_48_67=1.8
.ic q_49_67=0
.ic qb_49_67=1.8
.ic q_50_67=0
.ic qb_50_67=1.8
.ic q_51_67=0
.ic qb_51_67=1.8
.ic q_52_67=0
.ic qb_52_67=1.8
.ic q_53_67=0
.ic qb_53_67=1.8
.ic q_54_67=0
.ic qb_54_67=1.8
.ic q_55_67=0
.ic qb_55_67=1.8
.ic q_56_67=0
.ic qb_56_67=1.8
.ic q_57_67=0
.ic qb_57_67=1.8
.ic q_58_67=0
.ic qb_58_67=1.8
.ic q_59_67=0
.ic qb_59_67=1.8
.ic q_60_67=0
.ic qb_60_67=1.8
.ic q_61_67=0
.ic qb_61_67=1.8
.ic q_62_67=0
.ic qb_62_67=1.8
.ic q_63_67=0
.ic qb_63_67=1.8
.ic q_64_67=0
.ic qb_64_67=1.8
.ic q_65_67=0
.ic qb_65_67=1.8
.ic q_66_67=0
.ic qb_66_67=1.8
.ic q_67_67=0
.ic qb_67_67=1.8
.ic q_68_67=0
.ic qb_68_67=1.8
.ic q_69_67=0
.ic qb_69_67=1.8
.ic q_70_67=0
.ic qb_70_67=1.8
.ic q_71_67=0
.ic qb_71_67=1.8
.ic q_72_67=0
.ic qb_72_67=1.8
.ic q_73_67=0
.ic qb_73_67=1.8
.ic q_74_67=0
.ic qb_74_67=1.8
.ic q_75_67=0
.ic qb_75_67=1.8
.ic q_76_67=0
.ic qb_76_67=1.8
.ic q_77_67=0
.ic qb_77_67=1.8
.ic q_78_67=0
.ic qb_78_67=1.8
.ic q_79_67=0
.ic qb_79_67=1.8
.ic q_80_67=0
.ic qb_80_67=1.8
.ic q_81_67=0
.ic qb_81_67=1.8
.ic q_82_67=0
.ic qb_82_67=1.8
.ic q_83_67=0
.ic qb_83_67=1.8
.ic q_84_67=0
.ic qb_84_67=1.8
.ic q_85_67=0
.ic qb_85_67=1.8
.ic q_86_67=0
.ic qb_86_67=1.8
.ic q_87_67=0
.ic qb_87_67=1.8
.ic q_88_67=0
.ic qb_88_67=1.8
.ic q_89_67=0
.ic qb_89_67=1.8
.ic q_90_67=0
.ic qb_90_67=1.8
.ic q_91_67=0
.ic qb_91_67=1.8
.ic q_92_67=0
.ic qb_92_67=1.8
.ic q_93_67=0
.ic qb_93_67=1.8
.ic q_94_67=0
.ic qb_94_67=1.8
.ic q_95_67=0
.ic qb_95_67=1.8
.ic q_96_67=0
.ic qb_96_67=1.8
.ic q_97_67=0
.ic qb_97_67=1.8
.ic q_98_67=0
.ic qb_98_67=1.8
.ic q_99_67=0
.ic qb_99_67=1.8
.ic q_0_68=0
.ic qb_0_68=1.8
.ic q_1_68=0
.ic qb_1_68=1.8
.ic q_2_68=0
.ic qb_2_68=1.8
.ic q_3_68=0
.ic qb_3_68=1.8
.ic q_4_68=0
.ic qb_4_68=1.8
.ic q_5_68=0
.ic qb_5_68=1.8
.ic q_6_68=0
.ic qb_6_68=1.8
.ic q_7_68=0
.ic qb_7_68=1.8
.ic q_8_68=0
.ic qb_8_68=1.8
.ic q_9_68=0
.ic qb_9_68=1.8
.ic q_10_68=0
.ic qb_10_68=1.8
.ic q_11_68=0
.ic qb_11_68=1.8
.ic q_12_68=0
.ic qb_12_68=1.8
.ic q_13_68=0
.ic qb_13_68=1.8
.ic q_14_68=0
.ic qb_14_68=1.8
.ic q_15_68=0
.ic qb_15_68=1.8
.ic q_16_68=0
.ic qb_16_68=1.8
.ic q_17_68=0
.ic qb_17_68=1.8
.ic q_18_68=0
.ic qb_18_68=1.8
.ic q_19_68=0
.ic qb_19_68=1.8
.ic q_20_68=0
.ic qb_20_68=1.8
.ic q_21_68=0
.ic qb_21_68=1.8
.ic q_22_68=0
.ic qb_22_68=1.8
.ic q_23_68=0
.ic qb_23_68=1.8
.ic q_24_68=0
.ic qb_24_68=1.8
.ic q_25_68=0
.ic qb_25_68=1.8
.ic q_26_68=0
.ic qb_26_68=1.8
.ic q_27_68=0
.ic qb_27_68=1.8
.ic q_28_68=0
.ic qb_28_68=1.8
.ic q_29_68=0
.ic qb_29_68=1.8
.ic q_30_68=0
.ic qb_30_68=1.8
.ic q_31_68=0
.ic qb_31_68=1.8
.ic q_32_68=0
.ic qb_32_68=1.8
.ic q_33_68=0
.ic qb_33_68=1.8
.ic q_34_68=0
.ic qb_34_68=1.8
.ic q_35_68=0
.ic qb_35_68=1.8
.ic q_36_68=0
.ic qb_36_68=1.8
.ic q_37_68=0
.ic qb_37_68=1.8
.ic q_38_68=0
.ic qb_38_68=1.8
.ic q_39_68=0
.ic qb_39_68=1.8
.ic q_40_68=0
.ic qb_40_68=1.8
.ic q_41_68=0
.ic qb_41_68=1.8
.ic q_42_68=0
.ic qb_42_68=1.8
.ic q_43_68=0
.ic qb_43_68=1.8
.ic q_44_68=0
.ic qb_44_68=1.8
.ic q_45_68=0
.ic qb_45_68=1.8
.ic q_46_68=0
.ic qb_46_68=1.8
.ic q_47_68=0
.ic qb_47_68=1.8
.ic q_48_68=0
.ic qb_48_68=1.8
.ic q_49_68=0
.ic qb_49_68=1.8
.ic q_50_68=0
.ic qb_50_68=1.8
.ic q_51_68=0
.ic qb_51_68=1.8
.ic q_52_68=0
.ic qb_52_68=1.8
.ic q_53_68=0
.ic qb_53_68=1.8
.ic q_54_68=0
.ic qb_54_68=1.8
.ic q_55_68=0
.ic qb_55_68=1.8
.ic q_56_68=0
.ic qb_56_68=1.8
.ic q_57_68=0
.ic qb_57_68=1.8
.ic q_58_68=0
.ic qb_58_68=1.8
.ic q_59_68=0
.ic qb_59_68=1.8
.ic q_60_68=0
.ic qb_60_68=1.8
.ic q_61_68=0
.ic qb_61_68=1.8
.ic q_62_68=0
.ic qb_62_68=1.8
.ic q_63_68=0
.ic qb_63_68=1.8
.ic q_64_68=0
.ic qb_64_68=1.8
.ic q_65_68=0
.ic qb_65_68=1.8
.ic q_66_68=0
.ic qb_66_68=1.8
.ic q_67_68=0
.ic qb_67_68=1.8
.ic q_68_68=0
.ic qb_68_68=1.8
.ic q_69_68=0
.ic qb_69_68=1.8
.ic q_70_68=0
.ic qb_70_68=1.8
.ic q_71_68=0
.ic qb_71_68=1.8
.ic q_72_68=0
.ic qb_72_68=1.8
.ic q_73_68=0
.ic qb_73_68=1.8
.ic q_74_68=0
.ic qb_74_68=1.8
.ic q_75_68=0
.ic qb_75_68=1.8
.ic q_76_68=0
.ic qb_76_68=1.8
.ic q_77_68=0
.ic qb_77_68=1.8
.ic q_78_68=0
.ic qb_78_68=1.8
.ic q_79_68=0
.ic qb_79_68=1.8
.ic q_80_68=0
.ic qb_80_68=1.8
.ic q_81_68=0
.ic qb_81_68=1.8
.ic q_82_68=0
.ic qb_82_68=1.8
.ic q_83_68=0
.ic qb_83_68=1.8
.ic q_84_68=0
.ic qb_84_68=1.8
.ic q_85_68=0
.ic qb_85_68=1.8
.ic q_86_68=0
.ic qb_86_68=1.8
.ic q_87_68=0
.ic qb_87_68=1.8
.ic q_88_68=0
.ic qb_88_68=1.8
.ic q_89_68=0
.ic qb_89_68=1.8
.ic q_90_68=0
.ic qb_90_68=1.8
.ic q_91_68=0
.ic qb_91_68=1.8
.ic q_92_68=0
.ic qb_92_68=1.8
.ic q_93_68=0
.ic qb_93_68=1.8
.ic q_94_68=0
.ic qb_94_68=1.8
.ic q_95_68=0
.ic qb_95_68=1.8
.ic q_96_68=0
.ic qb_96_68=1.8
.ic q_97_68=0
.ic qb_97_68=1.8
.ic q_98_68=0
.ic qb_98_68=1.8
.ic q_99_68=0
.ic qb_99_68=1.8
.ic q_0_69=0
.ic qb_0_69=1.8
.ic q_1_69=0
.ic qb_1_69=1.8
.ic q_2_69=0
.ic qb_2_69=1.8
.ic q_3_69=0
.ic qb_3_69=1.8
.ic q_4_69=0
.ic qb_4_69=1.8
.ic q_5_69=0
.ic qb_5_69=1.8
.ic q_6_69=0
.ic qb_6_69=1.8
.ic q_7_69=0
.ic qb_7_69=1.8
.ic q_8_69=0
.ic qb_8_69=1.8
.ic q_9_69=0
.ic qb_9_69=1.8
.ic q_10_69=0
.ic qb_10_69=1.8
.ic q_11_69=0
.ic qb_11_69=1.8
.ic q_12_69=0
.ic qb_12_69=1.8
.ic q_13_69=0
.ic qb_13_69=1.8
.ic q_14_69=0
.ic qb_14_69=1.8
.ic q_15_69=0
.ic qb_15_69=1.8
.ic q_16_69=0
.ic qb_16_69=1.8
.ic q_17_69=0
.ic qb_17_69=1.8
.ic q_18_69=0
.ic qb_18_69=1.8
.ic q_19_69=0
.ic qb_19_69=1.8
.ic q_20_69=0
.ic qb_20_69=1.8
.ic q_21_69=0
.ic qb_21_69=1.8
.ic q_22_69=0
.ic qb_22_69=1.8
.ic q_23_69=0
.ic qb_23_69=1.8
.ic q_24_69=0
.ic qb_24_69=1.8
.ic q_25_69=0
.ic qb_25_69=1.8
.ic q_26_69=0
.ic qb_26_69=1.8
.ic q_27_69=0
.ic qb_27_69=1.8
.ic q_28_69=0
.ic qb_28_69=1.8
.ic q_29_69=0
.ic qb_29_69=1.8
.ic q_30_69=0
.ic qb_30_69=1.8
.ic q_31_69=0
.ic qb_31_69=1.8
.ic q_32_69=0
.ic qb_32_69=1.8
.ic q_33_69=0
.ic qb_33_69=1.8
.ic q_34_69=0
.ic qb_34_69=1.8
.ic q_35_69=0
.ic qb_35_69=1.8
.ic q_36_69=0
.ic qb_36_69=1.8
.ic q_37_69=0
.ic qb_37_69=1.8
.ic q_38_69=0
.ic qb_38_69=1.8
.ic q_39_69=0
.ic qb_39_69=1.8
.ic q_40_69=0
.ic qb_40_69=1.8
.ic q_41_69=0
.ic qb_41_69=1.8
.ic q_42_69=0
.ic qb_42_69=1.8
.ic q_43_69=0
.ic qb_43_69=1.8
.ic q_44_69=0
.ic qb_44_69=1.8
.ic q_45_69=0
.ic qb_45_69=1.8
.ic q_46_69=0
.ic qb_46_69=1.8
.ic q_47_69=0
.ic qb_47_69=1.8
.ic q_48_69=0
.ic qb_48_69=1.8
.ic q_49_69=0
.ic qb_49_69=1.8
.ic q_50_69=0
.ic qb_50_69=1.8
.ic q_51_69=0
.ic qb_51_69=1.8
.ic q_52_69=0
.ic qb_52_69=1.8
.ic q_53_69=0
.ic qb_53_69=1.8
.ic q_54_69=0
.ic qb_54_69=1.8
.ic q_55_69=0
.ic qb_55_69=1.8
.ic q_56_69=0
.ic qb_56_69=1.8
.ic q_57_69=0
.ic qb_57_69=1.8
.ic q_58_69=0
.ic qb_58_69=1.8
.ic q_59_69=0
.ic qb_59_69=1.8
.ic q_60_69=0
.ic qb_60_69=1.8
.ic q_61_69=0
.ic qb_61_69=1.8
.ic q_62_69=0
.ic qb_62_69=1.8
.ic q_63_69=0
.ic qb_63_69=1.8
.ic q_64_69=0
.ic qb_64_69=1.8
.ic q_65_69=0
.ic qb_65_69=1.8
.ic q_66_69=0
.ic qb_66_69=1.8
.ic q_67_69=0
.ic qb_67_69=1.8
.ic q_68_69=0
.ic qb_68_69=1.8
.ic q_69_69=0
.ic qb_69_69=1.8
.ic q_70_69=0
.ic qb_70_69=1.8
.ic q_71_69=0
.ic qb_71_69=1.8
.ic q_72_69=0
.ic qb_72_69=1.8
.ic q_73_69=0
.ic qb_73_69=1.8
.ic q_74_69=0
.ic qb_74_69=1.8
.ic q_75_69=0
.ic qb_75_69=1.8
.ic q_76_69=0
.ic qb_76_69=1.8
.ic q_77_69=0
.ic qb_77_69=1.8
.ic q_78_69=0
.ic qb_78_69=1.8
.ic q_79_69=0
.ic qb_79_69=1.8
.ic q_80_69=0
.ic qb_80_69=1.8
.ic q_81_69=0
.ic qb_81_69=1.8
.ic q_82_69=0
.ic qb_82_69=1.8
.ic q_83_69=0
.ic qb_83_69=1.8
.ic q_84_69=0
.ic qb_84_69=1.8
.ic q_85_69=0
.ic qb_85_69=1.8
.ic q_86_69=0
.ic qb_86_69=1.8
.ic q_87_69=0
.ic qb_87_69=1.8
.ic q_88_69=0
.ic qb_88_69=1.8
.ic q_89_69=0
.ic qb_89_69=1.8
.ic q_90_69=0
.ic qb_90_69=1.8
.ic q_91_69=0
.ic qb_91_69=1.8
.ic q_92_69=0
.ic qb_92_69=1.8
.ic q_93_69=0
.ic qb_93_69=1.8
.ic q_94_69=0
.ic qb_94_69=1.8
.ic q_95_69=0
.ic qb_95_69=1.8
.ic q_96_69=0
.ic qb_96_69=1.8
.ic q_97_69=0
.ic qb_97_69=1.8
.ic q_98_69=0
.ic qb_98_69=1.8
.ic q_99_69=0
.ic qb_99_69=1.8
.ic q_0_70=0
.ic qb_0_70=1.8
.ic q_1_70=0
.ic qb_1_70=1.8
.ic q_2_70=0
.ic qb_2_70=1.8
.ic q_3_70=0
.ic qb_3_70=1.8
.ic q_4_70=0
.ic qb_4_70=1.8
.ic q_5_70=0
.ic qb_5_70=1.8
.ic q_6_70=0
.ic qb_6_70=1.8
.ic q_7_70=0
.ic qb_7_70=1.8
.ic q_8_70=0
.ic qb_8_70=1.8
.ic q_9_70=0
.ic qb_9_70=1.8
.ic q_10_70=0
.ic qb_10_70=1.8
.ic q_11_70=0
.ic qb_11_70=1.8
.ic q_12_70=0
.ic qb_12_70=1.8
.ic q_13_70=0
.ic qb_13_70=1.8
.ic q_14_70=0
.ic qb_14_70=1.8
.ic q_15_70=0
.ic qb_15_70=1.8
.ic q_16_70=0
.ic qb_16_70=1.8
.ic q_17_70=0
.ic qb_17_70=1.8
.ic q_18_70=0
.ic qb_18_70=1.8
.ic q_19_70=0
.ic qb_19_70=1.8
.ic q_20_70=0
.ic qb_20_70=1.8
.ic q_21_70=0
.ic qb_21_70=1.8
.ic q_22_70=0
.ic qb_22_70=1.8
.ic q_23_70=0
.ic qb_23_70=1.8
.ic q_24_70=0
.ic qb_24_70=1.8
.ic q_25_70=0
.ic qb_25_70=1.8
.ic q_26_70=0
.ic qb_26_70=1.8
.ic q_27_70=0
.ic qb_27_70=1.8
.ic q_28_70=0
.ic qb_28_70=1.8
.ic q_29_70=0
.ic qb_29_70=1.8
.ic q_30_70=0
.ic qb_30_70=1.8
.ic q_31_70=0
.ic qb_31_70=1.8
.ic q_32_70=0
.ic qb_32_70=1.8
.ic q_33_70=0
.ic qb_33_70=1.8
.ic q_34_70=0
.ic qb_34_70=1.8
.ic q_35_70=0
.ic qb_35_70=1.8
.ic q_36_70=0
.ic qb_36_70=1.8
.ic q_37_70=0
.ic qb_37_70=1.8
.ic q_38_70=0
.ic qb_38_70=1.8
.ic q_39_70=0
.ic qb_39_70=1.8
.ic q_40_70=0
.ic qb_40_70=1.8
.ic q_41_70=0
.ic qb_41_70=1.8
.ic q_42_70=0
.ic qb_42_70=1.8
.ic q_43_70=0
.ic qb_43_70=1.8
.ic q_44_70=0
.ic qb_44_70=1.8
.ic q_45_70=0
.ic qb_45_70=1.8
.ic q_46_70=0
.ic qb_46_70=1.8
.ic q_47_70=0
.ic qb_47_70=1.8
.ic q_48_70=0
.ic qb_48_70=1.8
.ic q_49_70=0
.ic qb_49_70=1.8
.ic q_50_70=0
.ic qb_50_70=1.8
.ic q_51_70=0
.ic qb_51_70=1.8
.ic q_52_70=0
.ic qb_52_70=1.8
.ic q_53_70=0
.ic qb_53_70=1.8
.ic q_54_70=0
.ic qb_54_70=1.8
.ic q_55_70=0
.ic qb_55_70=1.8
.ic q_56_70=0
.ic qb_56_70=1.8
.ic q_57_70=0
.ic qb_57_70=1.8
.ic q_58_70=0
.ic qb_58_70=1.8
.ic q_59_70=0
.ic qb_59_70=1.8
.ic q_60_70=0
.ic qb_60_70=1.8
.ic q_61_70=0
.ic qb_61_70=1.8
.ic q_62_70=0
.ic qb_62_70=1.8
.ic q_63_70=0
.ic qb_63_70=1.8
.ic q_64_70=0
.ic qb_64_70=1.8
.ic q_65_70=0
.ic qb_65_70=1.8
.ic q_66_70=0
.ic qb_66_70=1.8
.ic q_67_70=0
.ic qb_67_70=1.8
.ic q_68_70=0
.ic qb_68_70=1.8
.ic q_69_70=0
.ic qb_69_70=1.8
.ic q_70_70=0
.ic qb_70_70=1.8
.ic q_71_70=0
.ic qb_71_70=1.8
.ic q_72_70=0
.ic qb_72_70=1.8
.ic q_73_70=0
.ic qb_73_70=1.8
.ic q_74_70=0
.ic qb_74_70=1.8
.ic q_75_70=0
.ic qb_75_70=1.8
.ic q_76_70=0
.ic qb_76_70=1.8
.ic q_77_70=0
.ic qb_77_70=1.8
.ic q_78_70=0
.ic qb_78_70=1.8
.ic q_79_70=0
.ic qb_79_70=1.8
.ic q_80_70=0
.ic qb_80_70=1.8
.ic q_81_70=0
.ic qb_81_70=1.8
.ic q_82_70=0
.ic qb_82_70=1.8
.ic q_83_70=0
.ic qb_83_70=1.8
.ic q_84_70=0
.ic qb_84_70=1.8
.ic q_85_70=0
.ic qb_85_70=1.8
.ic q_86_70=0
.ic qb_86_70=1.8
.ic q_87_70=0
.ic qb_87_70=1.8
.ic q_88_70=0
.ic qb_88_70=1.8
.ic q_89_70=0
.ic qb_89_70=1.8
.ic q_90_70=0
.ic qb_90_70=1.8
.ic q_91_70=0
.ic qb_91_70=1.8
.ic q_92_70=0
.ic qb_92_70=1.8
.ic q_93_70=0
.ic qb_93_70=1.8
.ic q_94_70=0
.ic qb_94_70=1.8
.ic q_95_70=0
.ic qb_95_70=1.8
.ic q_96_70=0
.ic qb_96_70=1.8
.ic q_97_70=0
.ic qb_97_70=1.8
.ic q_98_70=0
.ic qb_98_70=1.8
.ic q_99_70=0
.ic qb_99_70=1.8
.ic q_0_71=0
.ic qb_0_71=1.8
.ic q_1_71=0
.ic qb_1_71=1.8
.ic q_2_71=0
.ic qb_2_71=1.8
.ic q_3_71=0
.ic qb_3_71=1.8
.ic q_4_71=0
.ic qb_4_71=1.8
.ic q_5_71=0
.ic qb_5_71=1.8
.ic q_6_71=0
.ic qb_6_71=1.8
.ic q_7_71=0
.ic qb_7_71=1.8
.ic q_8_71=0
.ic qb_8_71=1.8
.ic q_9_71=0
.ic qb_9_71=1.8
.ic q_10_71=0
.ic qb_10_71=1.8
.ic q_11_71=0
.ic qb_11_71=1.8
.ic q_12_71=0
.ic qb_12_71=1.8
.ic q_13_71=0
.ic qb_13_71=1.8
.ic q_14_71=0
.ic qb_14_71=1.8
.ic q_15_71=0
.ic qb_15_71=1.8
.ic q_16_71=0
.ic qb_16_71=1.8
.ic q_17_71=0
.ic qb_17_71=1.8
.ic q_18_71=0
.ic qb_18_71=1.8
.ic q_19_71=0
.ic qb_19_71=1.8
.ic q_20_71=0
.ic qb_20_71=1.8
.ic q_21_71=0
.ic qb_21_71=1.8
.ic q_22_71=0
.ic qb_22_71=1.8
.ic q_23_71=0
.ic qb_23_71=1.8
.ic q_24_71=0
.ic qb_24_71=1.8
.ic q_25_71=0
.ic qb_25_71=1.8
.ic q_26_71=0
.ic qb_26_71=1.8
.ic q_27_71=0
.ic qb_27_71=1.8
.ic q_28_71=0
.ic qb_28_71=1.8
.ic q_29_71=0
.ic qb_29_71=1.8
.ic q_30_71=0
.ic qb_30_71=1.8
.ic q_31_71=0
.ic qb_31_71=1.8
.ic q_32_71=0
.ic qb_32_71=1.8
.ic q_33_71=0
.ic qb_33_71=1.8
.ic q_34_71=0
.ic qb_34_71=1.8
.ic q_35_71=0
.ic qb_35_71=1.8
.ic q_36_71=0
.ic qb_36_71=1.8
.ic q_37_71=0
.ic qb_37_71=1.8
.ic q_38_71=0
.ic qb_38_71=1.8
.ic q_39_71=0
.ic qb_39_71=1.8
.ic q_40_71=0
.ic qb_40_71=1.8
.ic q_41_71=0
.ic qb_41_71=1.8
.ic q_42_71=0
.ic qb_42_71=1.8
.ic q_43_71=0
.ic qb_43_71=1.8
.ic q_44_71=0
.ic qb_44_71=1.8
.ic q_45_71=0
.ic qb_45_71=1.8
.ic q_46_71=0
.ic qb_46_71=1.8
.ic q_47_71=0
.ic qb_47_71=1.8
.ic q_48_71=0
.ic qb_48_71=1.8
.ic q_49_71=0
.ic qb_49_71=1.8
.ic q_50_71=0
.ic qb_50_71=1.8
.ic q_51_71=0
.ic qb_51_71=1.8
.ic q_52_71=0
.ic qb_52_71=1.8
.ic q_53_71=0
.ic qb_53_71=1.8
.ic q_54_71=0
.ic qb_54_71=1.8
.ic q_55_71=0
.ic qb_55_71=1.8
.ic q_56_71=0
.ic qb_56_71=1.8
.ic q_57_71=0
.ic qb_57_71=1.8
.ic q_58_71=0
.ic qb_58_71=1.8
.ic q_59_71=0
.ic qb_59_71=1.8
.ic q_60_71=0
.ic qb_60_71=1.8
.ic q_61_71=0
.ic qb_61_71=1.8
.ic q_62_71=0
.ic qb_62_71=1.8
.ic q_63_71=0
.ic qb_63_71=1.8
.ic q_64_71=0
.ic qb_64_71=1.8
.ic q_65_71=0
.ic qb_65_71=1.8
.ic q_66_71=0
.ic qb_66_71=1.8
.ic q_67_71=0
.ic qb_67_71=1.8
.ic q_68_71=0
.ic qb_68_71=1.8
.ic q_69_71=0
.ic qb_69_71=1.8
.ic q_70_71=0
.ic qb_70_71=1.8
.ic q_71_71=0
.ic qb_71_71=1.8
.ic q_72_71=0
.ic qb_72_71=1.8
.ic q_73_71=0
.ic qb_73_71=1.8
.ic q_74_71=0
.ic qb_74_71=1.8
.ic q_75_71=0
.ic qb_75_71=1.8
.ic q_76_71=0
.ic qb_76_71=1.8
.ic q_77_71=0
.ic qb_77_71=1.8
.ic q_78_71=0
.ic qb_78_71=1.8
.ic q_79_71=0
.ic qb_79_71=1.8
.ic q_80_71=0
.ic qb_80_71=1.8
.ic q_81_71=0
.ic qb_81_71=1.8
.ic q_82_71=0
.ic qb_82_71=1.8
.ic q_83_71=0
.ic qb_83_71=1.8
.ic q_84_71=0
.ic qb_84_71=1.8
.ic q_85_71=0
.ic qb_85_71=1.8
.ic q_86_71=0
.ic qb_86_71=1.8
.ic q_87_71=0
.ic qb_87_71=1.8
.ic q_88_71=0
.ic qb_88_71=1.8
.ic q_89_71=0
.ic qb_89_71=1.8
.ic q_90_71=0
.ic qb_90_71=1.8
.ic q_91_71=0
.ic qb_91_71=1.8
.ic q_92_71=0
.ic qb_92_71=1.8
.ic q_93_71=0
.ic qb_93_71=1.8
.ic q_94_71=0
.ic qb_94_71=1.8
.ic q_95_71=0
.ic qb_95_71=1.8
.ic q_96_71=0
.ic qb_96_71=1.8
.ic q_97_71=0
.ic qb_97_71=1.8
.ic q_98_71=0
.ic qb_98_71=1.8
.ic q_99_71=0
.ic qb_99_71=1.8
.ic q_0_72=0
.ic qb_0_72=1.8
.ic q_1_72=0
.ic qb_1_72=1.8
.ic q_2_72=0
.ic qb_2_72=1.8
.ic q_3_72=0
.ic qb_3_72=1.8
.ic q_4_72=0
.ic qb_4_72=1.8
.ic q_5_72=0
.ic qb_5_72=1.8
.ic q_6_72=0
.ic qb_6_72=1.8
.ic q_7_72=0
.ic qb_7_72=1.8
.ic q_8_72=0
.ic qb_8_72=1.8
.ic q_9_72=0
.ic qb_9_72=1.8
.ic q_10_72=0
.ic qb_10_72=1.8
.ic q_11_72=0
.ic qb_11_72=1.8
.ic q_12_72=0
.ic qb_12_72=1.8
.ic q_13_72=0
.ic qb_13_72=1.8
.ic q_14_72=0
.ic qb_14_72=1.8
.ic q_15_72=0
.ic qb_15_72=1.8
.ic q_16_72=0
.ic qb_16_72=1.8
.ic q_17_72=0
.ic qb_17_72=1.8
.ic q_18_72=0
.ic qb_18_72=1.8
.ic q_19_72=0
.ic qb_19_72=1.8
.ic q_20_72=0
.ic qb_20_72=1.8
.ic q_21_72=0
.ic qb_21_72=1.8
.ic q_22_72=0
.ic qb_22_72=1.8
.ic q_23_72=0
.ic qb_23_72=1.8
.ic q_24_72=0
.ic qb_24_72=1.8
.ic q_25_72=0
.ic qb_25_72=1.8
.ic q_26_72=0
.ic qb_26_72=1.8
.ic q_27_72=0
.ic qb_27_72=1.8
.ic q_28_72=0
.ic qb_28_72=1.8
.ic q_29_72=0
.ic qb_29_72=1.8
.ic q_30_72=0
.ic qb_30_72=1.8
.ic q_31_72=0
.ic qb_31_72=1.8
.ic q_32_72=0
.ic qb_32_72=1.8
.ic q_33_72=0
.ic qb_33_72=1.8
.ic q_34_72=0
.ic qb_34_72=1.8
.ic q_35_72=0
.ic qb_35_72=1.8
.ic q_36_72=0
.ic qb_36_72=1.8
.ic q_37_72=0
.ic qb_37_72=1.8
.ic q_38_72=0
.ic qb_38_72=1.8
.ic q_39_72=0
.ic qb_39_72=1.8
.ic q_40_72=0
.ic qb_40_72=1.8
.ic q_41_72=0
.ic qb_41_72=1.8
.ic q_42_72=0
.ic qb_42_72=1.8
.ic q_43_72=0
.ic qb_43_72=1.8
.ic q_44_72=0
.ic qb_44_72=1.8
.ic q_45_72=0
.ic qb_45_72=1.8
.ic q_46_72=0
.ic qb_46_72=1.8
.ic q_47_72=0
.ic qb_47_72=1.8
.ic q_48_72=0
.ic qb_48_72=1.8
.ic q_49_72=0
.ic qb_49_72=1.8
.ic q_50_72=0
.ic qb_50_72=1.8
.ic q_51_72=0
.ic qb_51_72=1.8
.ic q_52_72=0
.ic qb_52_72=1.8
.ic q_53_72=0
.ic qb_53_72=1.8
.ic q_54_72=0
.ic qb_54_72=1.8
.ic q_55_72=0
.ic qb_55_72=1.8
.ic q_56_72=0
.ic qb_56_72=1.8
.ic q_57_72=0
.ic qb_57_72=1.8
.ic q_58_72=0
.ic qb_58_72=1.8
.ic q_59_72=0
.ic qb_59_72=1.8
.ic q_60_72=0
.ic qb_60_72=1.8
.ic q_61_72=0
.ic qb_61_72=1.8
.ic q_62_72=0
.ic qb_62_72=1.8
.ic q_63_72=0
.ic qb_63_72=1.8
.ic q_64_72=0
.ic qb_64_72=1.8
.ic q_65_72=0
.ic qb_65_72=1.8
.ic q_66_72=0
.ic qb_66_72=1.8
.ic q_67_72=0
.ic qb_67_72=1.8
.ic q_68_72=0
.ic qb_68_72=1.8
.ic q_69_72=0
.ic qb_69_72=1.8
.ic q_70_72=0
.ic qb_70_72=1.8
.ic q_71_72=0
.ic qb_71_72=1.8
.ic q_72_72=0
.ic qb_72_72=1.8
.ic q_73_72=0
.ic qb_73_72=1.8
.ic q_74_72=0
.ic qb_74_72=1.8
.ic q_75_72=0
.ic qb_75_72=1.8
.ic q_76_72=0
.ic qb_76_72=1.8
.ic q_77_72=0
.ic qb_77_72=1.8
.ic q_78_72=0
.ic qb_78_72=1.8
.ic q_79_72=0
.ic qb_79_72=1.8
.ic q_80_72=0
.ic qb_80_72=1.8
.ic q_81_72=0
.ic qb_81_72=1.8
.ic q_82_72=0
.ic qb_82_72=1.8
.ic q_83_72=0
.ic qb_83_72=1.8
.ic q_84_72=0
.ic qb_84_72=1.8
.ic q_85_72=0
.ic qb_85_72=1.8
.ic q_86_72=0
.ic qb_86_72=1.8
.ic q_87_72=0
.ic qb_87_72=1.8
.ic q_88_72=0
.ic qb_88_72=1.8
.ic q_89_72=0
.ic qb_89_72=1.8
.ic q_90_72=0
.ic qb_90_72=1.8
.ic q_91_72=0
.ic qb_91_72=1.8
.ic q_92_72=0
.ic qb_92_72=1.8
.ic q_93_72=0
.ic qb_93_72=1.8
.ic q_94_72=0
.ic qb_94_72=1.8
.ic q_95_72=0
.ic qb_95_72=1.8
.ic q_96_72=0
.ic qb_96_72=1.8
.ic q_97_72=0
.ic qb_97_72=1.8
.ic q_98_72=0
.ic qb_98_72=1.8
.ic q_99_72=0
.ic qb_99_72=1.8
.ic q_0_73=0
.ic qb_0_73=1.8
.ic q_1_73=0
.ic qb_1_73=1.8
.ic q_2_73=0
.ic qb_2_73=1.8
.ic q_3_73=0
.ic qb_3_73=1.8
.ic q_4_73=0
.ic qb_4_73=1.8
.ic q_5_73=0
.ic qb_5_73=1.8
.ic q_6_73=0
.ic qb_6_73=1.8
.ic q_7_73=0
.ic qb_7_73=1.8
.ic q_8_73=0
.ic qb_8_73=1.8
.ic q_9_73=0
.ic qb_9_73=1.8
.ic q_10_73=0
.ic qb_10_73=1.8
.ic q_11_73=0
.ic qb_11_73=1.8
.ic q_12_73=0
.ic qb_12_73=1.8
.ic q_13_73=0
.ic qb_13_73=1.8
.ic q_14_73=0
.ic qb_14_73=1.8
.ic q_15_73=0
.ic qb_15_73=1.8
.ic q_16_73=0
.ic qb_16_73=1.8
.ic q_17_73=0
.ic qb_17_73=1.8
.ic q_18_73=0
.ic qb_18_73=1.8
.ic q_19_73=0
.ic qb_19_73=1.8
.ic q_20_73=0
.ic qb_20_73=1.8
.ic q_21_73=0
.ic qb_21_73=1.8
.ic q_22_73=0
.ic qb_22_73=1.8
.ic q_23_73=0
.ic qb_23_73=1.8
.ic q_24_73=0
.ic qb_24_73=1.8
.ic q_25_73=0
.ic qb_25_73=1.8
.ic q_26_73=0
.ic qb_26_73=1.8
.ic q_27_73=0
.ic qb_27_73=1.8
.ic q_28_73=0
.ic qb_28_73=1.8
.ic q_29_73=0
.ic qb_29_73=1.8
.ic q_30_73=0
.ic qb_30_73=1.8
.ic q_31_73=0
.ic qb_31_73=1.8
.ic q_32_73=0
.ic qb_32_73=1.8
.ic q_33_73=0
.ic qb_33_73=1.8
.ic q_34_73=0
.ic qb_34_73=1.8
.ic q_35_73=0
.ic qb_35_73=1.8
.ic q_36_73=0
.ic qb_36_73=1.8
.ic q_37_73=0
.ic qb_37_73=1.8
.ic q_38_73=0
.ic qb_38_73=1.8
.ic q_39_73=0
.ic qb_39_73=1.8
.ic q_40_73=0
.ic qb_40_73=1.8
.ic q_41_73=0
.ic qb_41_73=1.8
.ic q_42_73=0
.ic qb_42_73=1.8
.ic q_43_73=0
.ic qb_43_73=1.8
.ic q_44_73=0
.ic qb_44_73=1.8
.ic q_45_73=0
.ic qb_45_73=1.8
.ic q_46_73=0
.ic qb_46_73=1.8
.ic q_47_73=0
.ic qb_47_73=1.8
.ic q_48_73=0
.ic qb_48_73=1.8
.ic q_49_73=0
.ic qb_49_73=1.8
.ic q_50_73=0
.ic qb_50_73=1.8
.ic q_51_73=0
.ic qb_51_73=1.8
.ic q_52_73=0
.ic qb_52_73=1.8
.ic q_53_73=0
.ic qb_53_73=1.8
.ic q_54_73=0
.ic qb_54_73=1.8
.ic q_55_73=0
.ic qb_55_73=1.8
.ic q_56_73=0
.ic qb_56_73=1.8
.ic q_57_73=0
.ic qb_57_73=1.8
.ic q_58_73=0
.ic qb_58_73=1.8
.ic q_59_73=0
.ic qb_59_73=1.8
.ic q_60_73=0
.ic qb_60_73=1.8
.ic q_61_73=0
.ic qb_61_73=1.8
.ic q_62_73=0
.ic qb_62_73=1.8
.ic q_63_73=0
.ic qb_63_73=1.8
.ic q_64_73=0
.ic qb_64_73=1.8
.ic q_65_73=0
.ic qb_65_73=1.8
.ic q_66_73=0
.ic qb_66_73=1.8
.ic q_67_73=0
.ic qb_67_73=1.8
.ic q_68_73=0
.ic qb_68_73=1.8
.ic q_69_73=0
.ic qb_69_73=1.8
.ic q_70_73=0
.ic qb_70_73=1.8
.ic q_71_73=0
.ic qb_71_73=1.8
.ic q_72_73=0
.ic qb_72_73=1.8
.ic q_73_73=0
.ic qb_73_73=1.8
.ic q_74_73=0
.ic qb_74_73=1.8
.ic q_75_73=0
.ic qb_75_73=1.8
.ic q_76_73=0
.ic qb_76_73=1.8
.ic q_77_73=0
.ic qb_77_73=1.8
.ic q_78_73=0
.ic qb_78_73=1.8
.ic q_79_73=0
.ic qb_79_73=1.8
.ic q_80_73=0
.ic qb_80_73=1.8
.ic q_81_73=0
.ic qb_81_73=1.8
.ic q_82_73=0
.ic qb_82_73=1.8
.ic q_83_73=0
.ic qb_83_73=1.8
.ic q_84_73=0
.ic qb_84_73=1.8
.ic q_85_73=0
.ic qb_85_73=1.8
.ic q_86_73=0
.ic qb_86_73=1.8
.ic q_87_73=0
.ic qb_87_73=1.8
.ic q_88_73=0
.ic qb_88_73=1.8
.ic q_89_73=0
.ic qb_89_73=1.8
.ic q_90_73=0
.ic qb_90_73=1.8
.ic q_91_73=0
.ic qb_91_73=1.8
.ic q_92_73=0
.ic qb_92_73=1.8
.ic q_93_73=0
.ic qb_93_73=1.8
.ic q_94_73=0
.ic qb_94_73=1.8
.ic q_95_73=0
.ic qb_95_73=1.8
.ic q_96_73=0
.ic qb_96_73=1.8
.ic q_97_73=0
.ic qb_97_73=1.8
.ic q_98_73=0
.ic qb_98_73=1.8
.ic q_99_73=0
.ic qb_99_73=1.8
.ic q_0_74=0
.ic qb_0_74=1.8
.ic q_1_74=0
.ic qb_1_74=1.8
.ic q_2_74=0
.ic qb_2_74=1.8
.ic q_3_74=0
.ic qb_3_74=1.8
.ic q_4_74=0
.ic qb_4_74=1.8
.ic q_5_74=0
.ic qb_5_74=1.8
.ic q_6_74=0
.ic qb_6_74=1.8
.ic q_7_74=0
.ic qb_7_74=1.8
.ic q_8_74=0
.ic qb_8_74=1.8
.ic q_9_74=0
.ic qb_9_74=1.8
.ic q_10_74=0
.ic qb_10_74=1.8
.ic q_11_74=0
.ic qb_11_74=1.8
.ic q_12_74=0
.ic qb_12_74=1.8
.ic q_13_74=0
.ic qb_13_74=1.8
.ic q_14_74=0
.ic qb_14_74=1.8
.ic q_15_74=0
.ic qb_15_74=1.8
.ic q_16_74=0
.ic qb_16_74=1.8
.ic q_17_74=0
.ic qb_17_74=1.8
.ic q_18_74=0
.ic qb_18_74=1.8
.ic q_19_74=0
.ic qb_19_74=1.8
.ic q_20_74=0
.ic qb_20_74=1.8
.ic q_21_74=0
.ic qb_21_74=1.8
.ic q_22_74=0
.ic qb_22_74=1.8
.ic q_23_74=0
.ic qb_23_74=1.8
.ic q_24_74=0
.ic qb_24_74=1.8
.ic q_25_74=0
.ic qb_25_74=1.8
.ic q_26_74=0
.ic qb_26_74=1.8
.ic q_27_74=0
.ic qb_27_74=1.8
.ic q_28_74=0
.ic qb_28_74=1.8
.ic q_29_74=0
.ic qb_29_74=1.8
.ic q_30_74=0
.ic qb_30_74=1.8
.ic q_31_74=0
.ic qb_31_74=1.8
.ic q_32_74=0
.ic qb_32_74=1.8
.ic q_33_74=0
.ic qb_33_74=1.8
.ic q_34_74=0
.ic qb_34_74=1.8
.ic q_35_74=0
.ic qb_35_74=1.8
.ic q_36_74=0
.ic qb_36_74=1.8
.ic q_37_74=0
.ic qb_37_74=1.8
.ic q_38_74=0
.ic qb_38_74=1.8
.ic q_39_74=0
.ic qb_39_74=1.8
.ic q_40_74=0
.ic qb_40_74=1.8
.ic q_41_74=0
.ic qb_41_74=1.8
.ic q_42_74=0
.ic qb_42_74=1.8
.ic q_43_74=0
.ic qb_43_74=1.8
.ic q_44_74=0
.ic qb_44_74=1.8
.ic q_45_74=0
.ic qb_45_74=1.8
.ic q_46_74=0
.ic qb_46_74=1.8
.ic q_47_74=0
.ic qb_47_74=1.8
.ic q_48_74=0
.ic qb_48_74=1.8
.ic q_49_74=0
.ic qb_49_74=1.8
.ic q_50_74=0
.ic qb_50_74=1.8
.ic q_51_74=0
.ic qb_51_74=1.8
.ic q_52_74=0
.ic qb_52_74=1.8
.ic q_53_74=0
.ic qb_53_74=1.8
.ic q_54_74=0
.ic qb_54_74=1.8
.ic q_55_74=0
.ic qb_55_74=1.8
.ic q_56_74=0
.ic qb_56_74=1.8
.ic q_57_74=0
.ic qb_57_74=1.8
.ic q_58_74=0
.ic qb_58_74=1.8
.ic q_59_74=0
.ic qb_59_74=1.8
.ic q_60_74=0
.ic qb_60_74=1.8
.ic q_61_74=0
.ic qb_61_74=1.8
.ic q_62_74=0
.ic qb_62_74=1.8
.ic q_63_74=0
.ic qb_63_74=1.8
.ic q_64_74=0
.ic qb_64_74=1.8
.ic q_65_74=0
.ic qb_65_74=1.8
.ic q_66_74=0
.ic qb_66_74=1.8
.ic q_67_74=0
.ic qb_67_74=1.8
.ic q_68_74=0
.ic qb_68_74=1.8
.ic q_69_74=0
.ic qb_69_74=1.8
.ic q_70_74=0
.ic qb_70_74=1.8
.ic q_71_74=0
.ic qb_71_74=1.8
.ic q_72_74=0
.ic qb_72_74=1.8
.ic q_73_74=0
.ic qb_73_74=1.8
.ic q_74_74=0
.ic qb_74_74=1.8
.ic q_75_74=0
.ic qb_75_74=1.8
.ic q_76_74=0
.ic qb_76_74=1.8
.ic q_77_74=0
.ic qb_77_74=1.8
.ic q_78_74=0
.ic qb_78_74=1.8
.ic q_79_74=0
.ic qb_79_74=1.8
.ic q_80_74=0
.ic qb_80_74=1.8
.ic q_81_74=0
.ic qb_81_74=1.8
.ic q_82_74=0
.ic qb_82_74=1.8
.ic q_83_74=0
.ic qb_83_74=1.8
.ic q_84_74=0
.ic qb_84_74=1.8
.ic q_85_74=0
.ic qb_85_74=1.8
.ic q_86_74=0
.ic qb_86_74=1.8
.ic q_87_74=0
.ic qb_87_74=1.8
.ic q_88_74=0
.ic qb_88_74=1.8
.ic q_89_74=0
.ic qb_89_74=1.8
.ic q_90_74=0
.ic qb_90_74=1.8
.ic q_91_74=0
.ic qb_91_74=1.8
.ic q_92_74=0
.ic qb_92_74=1.8
.ic q_93_74=0
.ic qb_93_74=1.8
.ic q_94_74=0
.ic qb_94_74=1.8
.ic q_95_74=0
.ic qb_95_74=1.8
.ic q_96_74=0
.ic qb_96_74=1.8
.ic q_97_74=0
.ic qb_97_74=1.8
.ic q_98_74=0
.ic qb_98_74=1.8
.ic q_99_74=0
.ic qb_99_74=1.8
.ic q_0_75=0
.ic qb_0_75=1.8
.ic q_1_75=0
.ic qb_1_75=1.8
.ic q_2_75=0
.ic qb_2_75=1.8
.ic q_3_75=0
.ic qb_3_75=1.8
.ic q_4_75=0
.ic qb_4_75=1.8
.ic q_5_75=0
.ic qb_5_75=1.8
.ic q_6_75=0
.ic qb_6_75=1.8
.ic q_7_75=0
.ic qb_7_75=1.8
.ic q_8_75=0
.ic qb_8_75=1.8
.ic q_9_75=0
.ic qb_9_75=1.8
.ic q_10_75=0
.ic qb_10_75=1.8
.ic q_11_75=0
.ic qb_11_75=1.8
.ic q_12_75=0
.ic qb_12_75=1.8
.ic q_13_75=0
.ic qb_13_75=1.8
.ic q_14_75=0
.ic qb_14_75=1.8
.ic q_15_75=0
.ic qb_15_75=1.8
.ic q_16_75=0
.ic qb_16_75=1.8
.ic q_17_75=0
.ic qb_17_75=1.8
.ic q_18_75=0
.ic qb_18_75=1.8
.ic q_19_75=0
.ic qb_19_75=1.8
.ic q_20_75=0
.ic qb_20_75=1.8
.ic q_21_75=0
.ic qb_21_75=1.8
.ic q_22_75=0
.ic qb_22_75=1.8
.ic q_23_75=0
.ic qb_23_75=1.8
.ic q_24_75=0
.ic qb_24_75=1.8
.ic q_25_75=0
.ic qb_25_75=1.8
.ic q_26_75=0
.ic qb_26_75=1.8
.ic q_27_75=0
.ic qb_27_75=1.8
.ic q_28_75=0
.ic qb_28_75=1.8
.ic q_29_75=0
.ic qb_29_75=1.8
.ic q_30_75=0
.ic qb_30_75=1.8
.ic q_31_75=0
.ic qb_31_75=1.8
.ic q_32_75=0
.ic qb_32_75=1.8
.ic q_33_75=0
.ic qb_33_75=1.8
.ic q_34_75=0
.ic qb_34_75=1.8
.ic q_35_75=0
.ic qb_35_75=1.8
.ic q_36_75=0
.ic qb_36_75=1.8
.ic q_37_75=0
.ic qb_37_75=1.8
.ic q_38_75=0
.ic qb_38_75=1.8
.ic q_39_75=0
.ic qb_39_75=1.8
.ic q_40_75=0
.ic qb_40_75=1.8
.ic q_41_75=0
.ic qb_41_75=1.8
.ic q_42_75=0
.ic qb_42_75=1.8
.ic q_43_75=0
.ic qb_43_75=1.8
.ic q_44_75=0
.ic qb_44_75=1.8
.ic q_45_75=0
.ic qb_45_75=1.8
.ic q_46_75=0
.ic qb_46_75=1.8
.ic q_47_75=0
.ic qb_47_75=1.8
.ic q_48_75=0
.ic qb_48_75=1.8
.ic q_49_75=0
.ic qb_49_75=1.8
.ic q_50_75=0
.ic qb_50_75=1.8
.ic q_51_75=0
.ic qb_51_75=1.8
.ic q_52_75=0
.ic qb_52_75=1.8
.ic q_53_75=0
.ic qb_53_75=1.8
.ic q_54_75=0
.ic qb_54_75=1.8
.ic q_55_75=0
.ic qb_55_75=1.8
.ic q_56_75=0
.ic qb_56_75=1.8
.ic q_57_75=0
.ic qb_57_75=1.8
.ic q_58_75=0
.ic qb_58_75=1.8
.ic q_59_75=0
.ic qb_59_75=1.8
.ic q_60_75=0
.ic qb_60_75=1.8
.ic q_61_75=0
.ic qb_61_75=1.8
.ic q_62_75=0
.ic qb_62_75=1.8
.ic q_63_75=0
.ic qb_63_75=1.8
.ic q_64_75=0
.ic qb_64_75=1.8
.ic q_65_75=0
.ic qb_65_75=1.8
.ic q_66_75=0
.ic qb_66_75=1.8
.ic q_67_75=0
.ic qb_67_75=1.8
.ic q_68_75=0
.ic qb_68_75=1.8
.ic q_69_75=0
.ic qb_69_75=1.8
.ic q_70_75=0
.ic qb_70_75=1.8
.ic q_71_75=0
.ic qb_71_75=1.8
.ic q_72_75=0
.ic qb_72_75=1.8
.ic q_73_75=0
.ic qb_73_75=1.8
.ic q_74_75=0
.ic qb_74_75=1.8
.ic q_75_75=0
.ic qb_75_75=1.8
.ic q_76_75=0
.ic qb_76_75=1.8
.ic q_77_75=0
.ic qb_77_75=1.8
.ic q_78_75=0
.ic qb_78_75=1.8
.ic q_79_75=0
.ic qb_79_75=1.8
.ic q_80_75=0
.ic qb_80_75=1.8
.ic q_81_75=0
.ic qb_81_75=1.8
.ic q_82_75=0
.ic qb_82_75=1.8
.ic q_83_75=0
.ic qb_83_75=1.8
.ic q_84_75=0
.ic qb_84_75=1.8
.ic q_85_75=0
.ic qb_85_75=1.8
.ic q_86_75=0
.ic qb_86_75=1.8
.ic q_87_75=0
.ic qb_87_75=1.8
.ic q_88_75=0
.ic qb_88_75=1.8
.ic q_89_75=0
.ic qb_89_75=1.8
.ic q_90_75=0
.ic qb_90_75=1.8
.ic q_91_75=0
.ic qb_91_75=1.8
.ic q_92_75=0
.ic qb_92_75=1.8
.ic q_93_75=0
.ic qb_93_75=1.8
.ic q_94_75=0
.ic qb_94_75=1.8
.ic q_95_75=0
.ic qb_95_75=1.8
.ic q_96_75=0
.ic qb_96_75=1.8
.ic q_97_75=0
.ic qb_97_75=1.8
.ic q_98_75=0
.ic qb_98_75=1.8
.ic q_99_75=0
.ic qb_99_75=1.8
.ic q_0_76=0
.ic qb_0_76=1.8
.ic q_1_76=0
.ic qb_1_76=1.8
.ic q_2_76=0
.ic qb_2_76=1.8
.ic q_3_76=0
.ic qb_3_76=1.8
.ic q_4_76=0
.ic qb_4_76=1.8
.ic q_5_76=0
.ic qb_5_76=1.8
.ic q_6_76=0
.ic qb_6_76=1.8
.ic q_7_76=0
.ic qb_7_76=1.8
.ic q_8_76=0
.ic qb_8_76=1.8
.ic q_9_76=0
.ic qb_9_76=1.8
.ic q_10_76=0
.ic qb_10_76=1.8
.ic q_11_76=0
.ic qb_11_76=1.8
.ic q_12_76=0
.ic qb_12_76=1.8
.ic q_13_76=0
.ic qb_13_76=1.8
.ic q_14_76=0
.ic qb_14_76=1.8
.ic q_15_76=0
.ic qb_15_76=1.8
.ic q_16_76=0
.ic qb_16_76=1.8
.ic q_17_76=0
.ic qb_17_76=1.8
.ic q_18_76=0
.ic qb_18_76=1.8
.ic q_19_76=0
.ic qb_19_76=1.8
.ic q_20_76=0
.ic qb_20_76=1.8
.ic q_21_76=0
.ic qb_21_76=1.8
.ic q_22_76=0
.ic qb_22_76=1.8
.ic q_23_76=0
.ic qb_23_76=1.8
.ic q_24_76=0
.ic qb_24_76=1.8
.ic q_25_76=0
.ic qb_25_76=1.8
.ic q_26_76=0
.ic qb_26_76=1.8
.ic q_27_76=0
.ic qb_27_76=1.8
.ic q_28_76=0
.ic qb_28_76=1.8
.ic q_29_76=0
.ic qb_29_76=1.8
.ic q_30_76=0
.ic qb_30_76=1.8
.ic q_31_76=0
.ic qb_31_76=1.8
.ic q_32_76=0
.ic qb_32_76=1.8
.ic q_33_76=0
.ic qb_33_76=1.8
.ic q_34_76=0
.ic qb_34_76=1.8
.ic q_35_76=0
.ic qb_35_76=1.8
.ic q_36_76=0
.ic qb_36_76=1.8
.ic q_37_76=0
.ic qb_37_76=1.8
.ic q_38_76=0
.ic qb_38_76=1.8
.ic q_39_76=0
.ic qb_39_76=1.8
.ic q_40_76=0
.ic qb_40_76=1.8
.ic q_41_76=0
.ic qb_41_76=1.8
.ic q_42_76=0
.ic qb_42_76=1.8
.ic q_43_76=0
.ic qb_43_76=1.8
.ic q_44_76=0
.ic qb_44_76=1.8
.ic q_45_76=0
.ic qb_45_76=1.8
.ic q_46_76=0
.ic qb_46_76=1.8
.ic q_47_76=0
.ic qb_47_76=1.8
.ic q_48_76=0
.ic qb_48_76=1.8
.ic q_49_76=0
.ic qb_49_76=1.8
.ic q_50_76=0
.ic qb_50_76=1.8
.ic q_51_76=0
.ic qb_51_76=1.8
.ic q_52_76=0
.ic qb_52_76=1.8
.ic q_53_76=0
.ic qb_53_76=1.8
.ic q_54_76=0
.ic qb_54_76=1.8
.ic q_55_76=0
.ic qb_55_76=1.8
.ic q_56_76=0
.ic qb_56_76=1.8
.ic q_57_76=0
.ic qb_57_76=1.8
.ic q_58_76=0
.ic qb_58_76=1.8
.ic q_59_76=0
.ic qb_59_76=1.8
.ic q_60_76=0
.ic qb_60_76=1.8
.ic q_61_76=0
.ic qb_61_76=1.8
.ic q_62_76=0
.ic qb_62_76=1.8
.ic q_63_76=0
.ic qb_63_76=1.8
.ic q_64_76=0
.ic qb_64_76=1.8
.ic q_65_76=0
.ic qb_65_76=1.8
.ic q_66_76=0
.ic qb_66_76=1.8
.ic q_67_76=0
.ic qb_67_76=1.8
.ic q_68_76=0
.ic qb_68_76=1.8
.ic q_69_76=0
.ic qb_69_76=1.8
.ic q_70_76=0
.ic qb_70_76=1.8
.ic q_71_76=0
.ic qb_71_76=1.8
.ic q_72_76=0
.ic qb_72_76=1.8
.ic q_73_76=0
.ic qb_73_76=1.8
.ic q_74_76=0
.ic qb_74_76=1.8
.ic q_75_76=0
.ic qb_75_76=1.8
.ic q_76_76=0
.ic qb_76_76=1.8
.ic q_77_76=0
.ic qb_77_76=1.8
.ic q_78_76=0
.ic qb_78_76=1.8
.ic q_79_76=0
.ic qb_79_76=1.8
.ic q_80_76=0
.ic qb_80_76=1.8
.ic q_81_76=0
.ic qb_81_76=1.8
.ic q_82_76=0
.ic qb_82_76=1.8
.ic q_83_76=0
.ic qb_83_76=1.8
.ic q_84_76=0
.ic qb_84_76=1.8
.ic q_85_76=0
.ic qb_85_76=1.8
.ic q_86_76=0
.ic qb_86_76=1.8
.ic q_87_76=0
.ic qb_87_76=1.8
.ic q_88_76=0
.ic qb_88_76=1.8
.ic q_89_76=0
.ic qb_89_76=1.8
.ic q_90_76=0
.ic qb_90_76=1.8
.ic q_91_76=0
.ic qb_91_76=1.8
.ic q_92_76=0
.ic qb_92_76=1.8
.ic q_93_76=0
.ic qb_93_76=1.8
.ic q_94_76=0
.ic qb_94_76=1.8
.ic q_95_76=0
.ic qb_95_76=1.8
.ic q_96_76=0
.ic qb_96_76=1.8
.ic q_97_76=0
.ic qb_97_76=1.8
.ic q_98_76=0
.ic qb_98_76=1.8
.ic q_99_76=0
.ic qb_99_76=1.8
.ic q_0_77=0
.ic qb_0_77=1.8
.ic q_1_77=0
.ic qb_1_77=1.8
.ic q_2_77=0
.ic qb_2_77=1.8
.ic q_3_77=0
.ic qb_3_77=1.8
.ic q_4_77=0
.ic qb_4_77=1.8
.ic q_5_77=0
.ic qb_5_77=1.8
.ic q_6_77=0
.ic qb_6_77=1.8
.ic q_7_77=0
.ic qb_7_77=1.8
.ic q_8_77=0
.ic qb_8_77=1.8
.ic q_9_77=0
.ic qb_9_77=1.8
.ic q_10_77=0
.ic qb_10_77=1.8
.ic q_11_77=0
.ic qb_11_77=1.8
.ic q_12_77=0
.ic qb_12_77=1.8
.ic q_13_77=0
.ic qb_13_77=1.8
.ic q_14_77=0
.ic qb_14_77=1.8
.ic q_15_77=0
.ic qb_15_77=1.8
.ic q_16_77=0
.ic qb_16_77=1.8
.ic q_17_77=0
.ic qb_17_77=1.8
.ic q_18_77=0
.ic qb_18_77=1.8
.ic q_19_77=0
.ic qb_19_77=1.8
.ic q_20_77=0
.ic qb_20_77=1.8
.ic q_21_77=0
.ic qb_21_77=1.8
.ic q_22_77=0
.ic qb_22_77=1.8
.ic q_23_77=0
.ic qb_23_77=1.8
.ic q_24_77=0
.ic qb_24_77=1.8
.ic q_25_77=0
.ic qb_25_77=1.8
.ic q_26_77=0
.ic qb_26_77=1.8
.ic q_27_77=0
.ic qb_27_77=1.8
.ic q_28_77=0
.ic qb_28_77=1.8
.ic q_29_77=0
.ic qb_29_77=1.8
.ic q_30_77=0
.ic qb_30_77=1.8
.ic q_31_77=0
.ic qb_31_77=1.8
.ic q_32_77=0
.ic qb_32_77=1.8
.ic q_33_77=0
.ic qb_33_77=1.8
.ic q_34_77=0
.ic qb_34_77=1.8
.ic q_35_77=0
.ic qb_35_77=1.8
.ic q_36_77=0
.ic qb_36_77=1.8
.ic q_37_77=0
.ic qb_37_77=1.8
.ic q_38_77=0
.ic qb_38_77=1.8
.ic q_39_77=0
.ic qb_39_77=1.8
.ic q_40_77=0
.ic qb_40_77=1.8
.ic q_41_77=0
.ic qb_41_77=1.8
.ic q_42_77=0
.ic qb_42_77=1.8
.ic q_43_77=0
.ic qb_43_77=1.8
.ic q_44_77=0
.ic qb_44_77=1.8
.ic q_45_77=0
.ic qb_45_77=1.8
.ic q_46_77=0
.ic qb_46_77=1.8
.ic q_47_77=0
.ic qb_47_77=1.8
.ic q_48_77=0
.ic qb_48_77=1.8
.ic q_49_77=0
.ic qb_49_77=1.8
.ic q_50_77=0
.ic qb_50_77=1.8
.ic q_51_77=0
.ic qb_51_77=1.8
.ic q_52_77=0
.ic qb_52_77=1.8
.ic q_53_77=0
.ic qb_53_77=1.8
.ic q_54_77=0
.ic qb_54_77=1.8
.ic q_55_77=0
.ic qb_55_77=1.8
.ic q_56_77=0
.ic qb_56_77=1.8
.ic q_57_77=0
.ic qb_57_77=1.8
.ic q_58_77=0
.ic qb_58_77=1.8
.ic q_59_77=0
.ic qb_59_77=1.8
.ic q_60_77=0
.ic qb_60_77=1.8
.ic q_61_77=0
.ic qb_61_77=1.8
.ic q_62_77=0
.ic qb_62_77=1.8
.ic q_63_77=0
.ic qb_63_77=1.8
.ic q_64_77=0
.ic qb_64_77=1.8
.ic q_65_77=0
.ic qb_65_77=1.8
.ic q_66_77=0
.ic qb_66_77=1.8
.ic q_67_77=0
.ic qb_67_77=1.8
.ic q_68_77=0
.ic qb_68_77=1.8
.ic q_69_77=0
.ic qb_69_77=1.8
.ic q_70_77=0
.ic qb_70_77=1.8
.ic q_71_77=0
.ic qb_71_77=1.8
.ic q_72_77=0
.ic qb_72_77=1.8
.ic q_73_77=0
.ic qb_73_77=1.8
.ic q_74_77=0
.ic qb_74_77=1.8
.ic q_75_77=0
.ic qb_75_77=1.8
.ic q_76_77=0
.ic qb_76_77=1.8
.ic q_77_77=0
.ic qb_77_77=1.8
.ic q_78_77=0
.ic qb_78_77=1.8
.ic q_79_77=0
.ic qb_79_77=1.8
.ic q_80_77=0
.ic qb_80_77=1.8
.ic q_81_77=0
.ic qb_81_77=1.8
.ic q_82_77=0
.ic qb_82_77=1.8
.ic q_83_77=0
.ic qb_83_77=1.8
.ic q_84_77=0
.ic qb_84_77=1.8
.ic q_85_77=0
.ic qb_85_77=1.8
.ic q_86_77=0
.ic qb_86_77=1.8
.ic q_87_77=0
.ic qb_87_77=1.8
.ic q_88_77=0
.ic qb_88_77=1.8
.ic q_89_77=0
.ic qb_89_77=1.8
.ic q_90_77=0
.ic qb_90_77=1.8
.ic q_91_77=0
.ic qb_91_77=1.8
.ic q_92_77=0
.ic qb_92_77=1.8
.ic q_93_77=0
.ic qb_93_77=1.8
.ic q_94_77=0
.ic qb_94_77=1.8
.ic q_95_77=0
.ic qb_95_77=1.8
.ic q_96_77=0
.ic qb_96_77=1.8
.ic q_97_77=0
.ic qb_97_77=1.8
.ic q_98_77=0
.ic qb_98_77=1.8
.ic q_99_77=0
.ic qb_99_77=1.8
.ic q_0_78=0
.ic qb_0_78=1.8
.ic q_1_78=0
.ic qb_1_78=1.8
.ic q_2_78=0
.ic qb_2_78=1.8
.ic q_3_78=0
.ic qb_3_78=1.8
.ic q_4_78=0
.ic qb_4_78=1.8
.ic q_5_78=0
.ic qb_5_78=1.8
.ic q_6_78=0
.ic qb_6_78=1.8
.ic q_7_78=0
.ic qb_7_78=1.8
.ic q_8_78=0
.ic qb_8_78=1.8
.ic q_9_78=0
.ic qb_9_78=1.8
.ic q_10_78=0
.ic qb_10_78=1.8
.ic q_11_78=0
.ic qb_11_78=1.8
.ic q_12_78=0
.ic qb_12_78=1.8
.ic q_13_78=0
.ic qb_13_78=1.8
.ic q_14_78=0
.ic qb_14_78=1.8
.ic q_15_78=0
.ic qb_15_78=1.8
.ic q_16_78=0
.ic qb_16_78=1.8
.ic q_17_78=0
.ic qb_17_78=1.8
.ic q_18_78=0
.ic qb_18_78=1.8
.ic q_19_78=0
.ic qb_19_78=1.8
.ic q_20_78=0
.ic qb_20_78=1.8
.ic q_21_78=0
.ic qb_21_78=1.8
.ic q_22_78=0
.ic qb_22_78=1.8
.ic q_23_78=0
.ic qb_23_78=1.8
.ic q_24_78=0
.ic qb_24_78=1.8
.ic q_25_78=0
.ic qb_25_78=1.8
.ic q_26_78=0
.ic qb_26_78=1.8
.ic q_27_78=0
.ic qb_27_78=1.8
.ic q_28_78=0
.ic qb_28_78=1.8
.ic q_29_78=0
.ic qb_29_78=1.8
.ic q_30_78=0
.ic qb_30_78=1.8
.ic q_31_78=0
.ic qb_31_78=1.8
.ic q_32_78=0
.ic qb_32_78=1.8
.ic q_33_78=0
.ic qb_33_78=1.8
.ic q_34_78=0
.ic qb_34_78=1.8
.ic q_35_78=0
.ic qb_35_78=1.8
.ic q_36_78=0
.ic qb_36_78=1.8
.ic q_37_78=0
.ic qb_37_78=1.8
.ic q_38_78=0
.ic qb_38_78=1.8
.ic q_39_78=0
.ic qb_39_78=1.8
.ic q_40_78=0
.ic qb_40_78=1.8
.ic q_41_78=0
.ic qb_41_78=1.8
.ic q_42_78=0
.ic qb_42_78=1.8
.ic q_43_78=0
.ic qb_43_78=1.8
.ic q_44_78=0
.ic qb_44_78=1.8
.ic q_45_78=0
.ic qb_45_78=1.8
.ic q_46_78=0
.ic qb_46_78=1.8
.ic q_47_78=0
.ic qb_47_78=1.8
.ic q_48_78=0
.ic qb_48_78=1.8
.ic q_49_78=0
.ic qb_49_78=1.8
.ic q_50_78=0
.ic qb_50_78=1.8
.ic q_51_78=0
.ic qb_51_78=1.8
.ic q_52_78=0
.ic qb_52_78=1.8
.ic q_53_78=0
.ic qb_53_78=1.8
.ic q_54_78=0
.ic qb_54_78=1.8
.ic q_55_78=0
.ic qb_55_78=1.8
.ic q_56_78=0
.ic qb_56_78=1.8
.ic q_57_78=0
.ic qb_57_78=1.8
.ic q_58_78=0
.ic qb_58_78=1.8
.ic q_59_78=0
.ic qb_59_78=1.8
.ic q_60_78=0
.ic qb_60_78=1.8
.ic q_61_78=0
.ic qb_61_78=1.8
.ic q_62_78=0
.ic qb_62_78=1.8
.ic q_63_78=0
.ic qb_63_78=1.8
.ic q_64_78=0
.ic qb_64_78=1.8
.ic q_65_78=0
.ic qb_65_78=1.8
.ic q_66_78=0
.ic qb_66_78=1.8
.ic q_67_78=0
.ic qb_67_78=1.8
.ic q_68_78=0
.ic qb_68_78=1.8
.ic q_69_78=0
.ic qb_69_78=1.8
.ic q_70_78=0
.ic qb_70_78=1.8
.ic q_71_78=0
.ic qb_71_78=1.8
.ic q_72_78=0
.ic qb_72_78=1.8
.ic q_73_78=0
.ic qb_73_78=1.8
.ic q_74_78=0
.ic qb_74_78=1.8
.ic q_75_78=0
.ic qb_75_78=1.8
.ic q_76_78=0
.ic qb_76_78=1.8
.ic q_77_78=0
.ic qb_77_78=1.8
.ic q_78_78=0
.ic qb_78_78=1.8
.ic q_79_78=0
.ic qb_79_78=1.8
.ic q_80_78=0
.ic qb_80_78=1.8
.ic q_81_78=0
.ic qb_81_78=1.8
.ic q_82_78=0
.ic qb_82_78=1.8
.ic q_83_78=0
.ic qb_83_78=1.8
.ic q_84_78=0
.ic qb_84_78=1.8
.ic q_85_78=0
.ic qb_85_78=1.8
.ic q_86_78=0
.ic qb_86_78=1.8
.ic q_87_78=0
.ic qb_87_78=1.8
.ic q_88_78=0
.ic qb_88_78=1.8
.ic q_89_78=0
.ic qb_89_78=1.8
.ic q_90_78=0
.ic qb_90_78=1.8
.ic q_91_78=0
.ic qb_91_78=1.8
.ic q_92_78=0
.ic qb_92_78=1.8
.ic q_93_78=0
.ic qb_93_78=1.8
.ic q_94_78=0
.ic qb_94_78=1.8
.ic q_95_78=0
.ic qb_95_78=1.8
.ic q_96_78=0
.ic qb_96_78=1.8
.ic q_97_78=0
.ic qb_97_78=1.8
.ic q_98_78=0
.ic qb_98_78=1.8
.ic q_99_78=0
.ic qb_99_78=1.8
.ic q_0_79=0
.ic qb_0_79=1.8
.ic q_1_79=0
.ic qb_1_79=1.8
.ic q_2_79=0
.ic qb_2_79=1.8
.ic q_3_79=0
.ic qb_3_79=1.8
.ic q_4_79=0
.ic qb_4_79=1.8
.ic q_5_79=0
.ic qb_5_79=1.8
.ic q_6_79=0
.ic qb_6_79=1.8
.ic q_7_79=0
.ic qb_7_79=1.8
.ic q_8_79=0
.ic qb_8_79=1.8
.ic q_9_79=0
.ic qb_9_79=1.8
.ic q_10_79=0
.ic qb_10_79=1.8
.ic q_11_79=0
.ic qb_11_79=1.8
.ic q_12_79=0
.ic qb_12_79=1.8
.ic q_13_79=0
.ic qb_13_79=1.8
.ic q_14_79=0
.ic qb_14_79=1.8
.ic q_15_79=0
.ic qb_15_79=1.8
.ic q_16_79=0
.ic qb_16_79=1.8
.ic q_17_79=0
.ic qb_17_79=1.8
.ic q_18_79=0
.ic qb_18_79=1.8
.ic q_19_79=0
.ic qb_19_79=1.8
.ic q_20_79=0
.ic qb_20_79=1.8
.ic q_21_79=0
.ic qb_21_79=1.8
.ic q_22_79=0
.ic qb_22_79=1.8
.ic q_23_79=0
.ic qb_23_79=1.8
.ic q_24_79=0
.ic qb_24_79=1.8
.ic q_25_79=0
.ic qb_25_79=1.8
.ic q_26_79=0
.ic qb_26_79=1.8
.ic q_27_79=0
.ic qb_27_79=1.8
.ic q_28_79=0
.ic qb_28_79=1.8
.ic q_29_79=0
.ic qb_29_79=1.8
.ic q_30_79=0
.ic qb_30_79=1.8
.ic q_31_79=0
.ic qb_31_79=1.8
.ic q_32_79=0
.ic qb_32_79=1.8
.ic q_33_79=0
.ic qb_33_79=1.8
.ic q_34_79=0
.ic qb_34_79=1.8
.ic q_35_79=0
.ic qb_35_79=1.8
.ic q_36_79=0
.ic qb_36_79=1.8
.ic q_37_79=0
.ic qb_37_79=1.8
.ic q_38_79=0
.ic qb_38_79=1.8
.ic q_39_79=0
.ic qb_39_79=1.8
.ic q_40_79=0
.ic qb_40_79=1.8
.ic q_41_79=0
.ic qb_41_79=1.8
.ic q_42_79=0
.ic qb_42_79=1.8
.ic q_43_79=0
.ic qb_43_79=1.8
.ic q_44_79=0
.ic qb_44_79=1.8
.ic q_45_79=0
.ic qb_45_79=1.8
.ic q_46_79=0
.ic qb_46_79=1.8
.ic q_47_79=0
.ic qb_47_79=1.8
.ic q_48_79=0
.ic qb_48_79=1.8
.ic q_49_79=0
.ic qb_49_79=1.8
.ic q_50_79=0
.ic qb_50_79=1.8
.ic q_51_79=0
.ic qb_51_79=1.8
.ic q_52_79=0
.ic qb_52_79=1.8
.ic q_53_79=0
.ic qb_53_79=1.8
.ic q_54_79=0
.ic qb_54_79=1.8
.ic q_55_79=0
.ic qb_55_79=1.8
.ic q_56_79=0
.ic qb_56_79=1.8
.ic q_57_79=0
.ic qb_57_79=1.8
.ic q_58_79=0
.ic qb_58_79=1.8
.ic q_59_79=0
.ic qb_59_79=1.8
.ic q_60_79=0
.ic qb_60_79=1.8
.ic q_61_79=0
.ic qb_61_79=1.8
.ic q_62_79=0
.ic qb_62_79=1.8
.ic q_63_79=0
.ic qb_63_79=1.8
.ic q_64_79=0
.ic qb_64_79=1.8
.ic q_65_79=0
.ic qb_65_79=1.8
.ic q_66_79=0
.ic qb_66_79=1.8
.ic q_67_79=0
.ic qb_67_79=1.8
.ic q_68_79=0
.ic qb_68_79=1.8
.ic q_69_79=0
.ic qb_69_79=1.8
.ic q_70_79=0
.ic qb_70_79=1.8
.ic q_71_79=0
.ic qb_71_79=1.8
.ic q_72_79=0
.ic qb_72_79=1.8
.ic q_73_79=0
.ic qb_73_79=1.8
.ic q_74_79=0
.ic qb_74_79=1.8
.ic q_75_79=0
.ic qb_75_79=1.8
.ic q_76_79=0
.ic qb_76_79=1.8
.ic q_77_79=0
.ic qb_77_79=1.8
.ic q_78_79=0
.ic qb_78_79=1.8
.ic q_79_79=0
.ic qb_79_79=1.8
.ic q_80_79=0
.ic qb_80_79=1.8
.ic q_81_79=0
.ic qb_81_79=1.8
.ic q_82_79=0
.ic qb_82_79=1.8
.ic q_83_79=0
.ic qb_83_79=1.8
.ic q_84_79=0
.ic qb_84_79=1.8
.ic q_85_79=0
.ic qb_85_79=1.8
.ic q_86_79=0
.ic qb_86_79=1.8
.ic q_87_79=0
.ic qb_87_79=1.8
.ic q_88_79=0
.ic qb_88_79=1.8
.ic q_89_79=0
.ic qb_89_79=1.8
.ic q_90_79=0
.ic qb_90_79=1.8
.ic q_91_79=0
.ic qb_91_79=1.8
.ic q_92_79=0
.ic qb_92_79=1.8
.ic q_93_79=0
.ic qb_93_79=1.8
.ic q_94_79=0
.ic qb_94_79=1.8
.ic q_95_79=0
.ic qb_95_79=1.8
.ic q_96_79=0
.ic qb_96_79=1.8
.ic q_97_79=0
.ic qb_97_79=1.8
.ic q_98_79=0
.ic qb_98_79=1.8
.ic q_99_79=0
.ic qb_99_79=1.8
.ic q_0_80=0
.ic qb_0_80=1.8
.ic q_1_80=0
.ic qb_1_80=1.8
.ic q_2_80=0
.ic qb_2_80=1.8
.ic q_3_80=0
.ic qb_3_80=1.8
.ic q_4_80=0
.ic qb_4_80=1.8
.ic q_5_80=0
.ic qb_5_80=1.8
.ic q_6_80=0
.ic qb_6_80=1.8
.ic q_7_80=0
.ic qb_7_80=1.8
.ic q_8_80=0
.ic qb_8_80=1.8
.ic q_9_80=0
.ic qb_9_80=1.8
.ic q_10_80=0
.ic qb_10_80=1.8
.ic q_11_80=0
.ic qb_11_80=1.8
.ic q_12_80=0
.ic qb_12_80=1.8
.ic q_13_80=0
.ic qb_13_80=1.8
.ic q_14_80=0
.ic qb_14_80=1.8
.ic q_15_80=0
.ic qb_15_80=1.8
.ic q_16_80=0
.ic qb_16_80=1.8
.ic q_17_80=0
.ic qb_17_80=1.8
.ic q_18_80=0
.ic qb_18_80=1.8
.ic q_19_80=0
.ic qb_19_80=1.8
.ic q_20_80=0
.ic qb_20_80=1.8
.ic q_21_80=0
.ic qb_21_80=1.8
.ic q_22_80=0
.ic qb_22_80=1.8
.ic q_23_80=0
.ic qb_23_80=1.8
.ic q_24_80=0
.ic qb_24_80=1.8
.ic q_25_80=0
.ic qb_25_80=1.8
.ic q_26_80=0
.ic qb_26_80=1.8
.ic q_27_80=0
.ic qb_27_80=1.8
.ic q_28_80=0
.ic qb_28_80=1.8
.ic q_29_80=0
.ic qb_29_80=1.8
.ic q_30_80=0
.ic qb_30_80=1.8
.ic q_31_80=0
.ic qb_31_80=1.8
.ic q_32_80=0
.ic qb_32_80=1.8
.ic q_33_80=0
.ic qb_33_80=1.8
.ic q_34_80=0
.ic qb_34_80=1.8
.ic q_35_80=0
.ic qb_35_80=1.8
.ic q_36_80=0
.ic qb_36_80=1.8
.ic q_37_80=0
.ic qb_37_80=1.8
.ic q_38_80=0
.ic qb_38_80=1.8
.ic q_39_80=0
.ic qb_39_80=1.8
.ic q_40_80=0
.ic qb_40_80=1.8
.ic q_41_80=0
.ic qb_41_80=1.8
.ic q_42_80=0
.ic qb_42_80=1.8
.ic q_43_80=0
.ic qb_43_80=1.8
.ic q_44_80=0
.ic qb_44_80=1.8
.ic q_45_80=0
.ic qb_45_80=1.8
.ic q_46_80=0
.ic qb_46_80=1.8
.ic q_47_80=0
.ic qb_47_80=1.8
.ic q_48_80=0
.ic qb_48_80=1.8
.ic q_49_80=0
.ic qb_49_80=1.8
.ic q_50_80=0
.ic qb_50_80=1.8
.ic q_51_80=0
.ic qb_51_80=1.8
.ic q_52_80=0
.ic qb_52_80=1.8
.ic q_53_80=0
.ic qb_53_80=1.8
.ic q_54_80=0
.ic qb_54_80=1.8
.ic q_55_80=0
.ic qb_55_80=1.8
.ic q_56_80=0
.ic qb_56_80=1.8
.ic q_57_80=0
.ic qb_57_80=1.8
.ic q_58_80=0
.ic qb_58_80=1.8
.ic q_59_80=0
.ic qb_59_80=1.8
.ic q_60_80=0
.ic qb_60_80=1.8
.ic q_61_80=0
.ic qb_61_80=1.8
.ic q_62_80=0
.ic qb_62_80=1.8
.ic q_63_80=0
.ic qb_63_80=1.8
.ic q_64_80=0
.ic qb_64_80=1.8
.ic q_65_80=0
.ic qb_65_80=1.8
.ic q_66_80=0
.ic qb_66_80=1.8
.ic q_67_80=0
.ic qb_67_80=1.8
.ic q_68_80=0
.ic qb_68_80=1.8
.ic q_69_80=0
.ic qb_69_80=1.8
.ic q_70_80=0
.ic qb_70_80=1.8
.ic q_71_80=0
.ic qb_71_80=1.8
.ic q_72_80=0
.ic qb_72_80=1.8
.ic q_73_80=0
.ic qb_73_80=1.8
.ic q_74_80=0
.ic qb_74_80=1.8
.ic q_75_80=0
.ic qb_75_80=1.8
.ic q_76_80=0
.ic qb_76_80=1.8
.ic q_77_80=0
.ic qb_77_80=1.8
.ic q_78_80=0
.ic qb_78_80=1.8
.ic q_79_80=0
.ic qb_79_80=1.8
.ic q_80_80=0
.ic qb_80_80=1.8
.ic q_81_80=0
.ic qb_81_80=1.8
.ic q_82_80=0
.ic qb_82_80=1.8
.ic q_83_80=0
.ic qb_83_80=1.8
.ic q_84_80=0
.ic qb_84_80=1.8
.ic q_85_80=0
.ic qb_85_80=1.8
.ic q_86_80=0
.ic qb_86_80=1.8
.ic q_87_80=0
.ic qb_87_80=1.8
.ic q_88_80=0
.ic qb_88_80=1.8
.ic q_89_80=0
.ic qb_89_80=1.8
.ic q_90_80=0
.ic qb_90_80=1.8
.ic q_91_80=0
.ic qb_91_80=1.8
.ic q_92_80=0
.ic qb_92_80=1.8
.ic q_93_80=0
.ic qb_93_80=1.8
.ic q_94_80=0
.ic qb_94_80=1.8
.ic q_95_80=0
.ic qb_95_80=1.8
.ic q_96_80=0
.ic qb_96_80=1.8
.ic q_97_80=0
.ic qb_97_80=1.8
.ic q_98_80=0
.ic qb_98_80=1.8
.ic q_99_80=0
.ic qb_99_80=1.8
.ic q_0_81=0
.ic qb_0_81=1.8
.ic q_1_81=0
.ic qb_1_81=1.8
.ic q_2_81=0
.ic qb_2_81=1.8
.ic q_3_81=0
.ic qb_3_81=1.8
.ic q_4_81=0
.ic qb_4_81=1.8
.ic q_5_81=0
.ic qb_5_81=1.8
.ic q_6_81=0
.ic qb_6_81=1.8
.ic q_7_81=0
.ic qb_7_81=1.8
.ic q_8_81=0
.ic qb_8_81=1.8
.ic q_9_81=0
.ic qb_9_81=1.8
.ic q_10_81=0
.ic qb_10_81=1.8
.ic q_11_81=0
.ic qb_11_81=1.8
.ic q_12_81=0
.ic qb_12_81=1.8
.ic q_13_81=0
.ic qb_13_81=1.8
.ic q_14_81=0
.ic qb_14_81=1.8
.ic q_15_81=0
.ic qb_15_81=1.8
.ic q_16_81=0
.ic qb_16_81=1.8
.ic q_17_81=0
.ic qb_17_81=1.8
.ic q_18_81=0
.ic qb_18_81=1.8
.ic q_19_81=0
.ic qb_19_81=1.8
.ic q_20_81=0
.ic qb_20_81=1.8
.ic q_21_81=0
.ic qb_21_81=1.8
.ic q_22_81=0
.ic qb_22_81=1.8
.ic q_23_81=0
.ic qb_23_81=1.8
.ic q_24_81=0
.ic qb_24_81=1.8
.ic q_25_81=0
.ic qb_25_81=1.8
.ic q_26_81=0
.ic qb_26_81=1.8
.ic q_27_81=0
.ic qb_27_81=1.8
.ic q_28_81=0
.ic qb_28_81=1.8
.ic q_29_81=0
.ic qb_29_81=1.8
.ic q_30_81=0
.ic qb_30_81=1.8
.ic q_31_81=0
.ic qb_31_81=1.8
.ic q_32_81=0
.ic qb_32_81=1.8
.ic q_33_81=0
.ic qb_33_81=1.8
.ic q_34_81=0
.ic qb_34_81=1.8
.ic q_35_81=0
.ic qb_35_81=1.8
.ic q_36_81=0
.ic qb_36_81=1.8
.ic q_37_81=0
.ic qb_37_81=1.8
.ic q_38_81=0
.ic qb_38_81=1.8
.ic q_39_81=0
.ic qb_39_81=1.8
.ic q_40_81=0
.ic qb_40_81=1.8
.ic q_41_81=0
.ic qb_41_81=1.8
.ic q_42_81=0
.ic qb_42_81=1.8
.ic q_43_81=0
.ic qb_43_81=1.8
.ic q_44_81=0
.ic qb_44_81=1.8
.ic q_45_81=0
.ic qb_45_81=1.8
.ic q_46_81=0
.ic qb_46_81=1.8
.ic q_47_81=0
.ic qb_47_81=1.8
.ic q_48_81=0
.ic qb_48_81=1.8
.ic q_49_81=0
.ic qb_49_81=1.8
.ic q_50_81=0
.ic qb_50_81=1.8
.ic q_51_81=0
.ic qb_51_81=1.8
.ic q_52_81=0
.ic qb_52_81=1.8
.ic q_53_81=0
.ic qb_53_81=1.8
.ic q_54_81=0
.ic qb_54_81=1.8
.ic q_55_81=0
.ic qb_55_81=1.8
.ic q_56_81=0
.ic qb_56_81=1.8
.ic q_57_81=0
.ic qb_57_81=1.8
.ic q_58_81=0
.ic qb_58_81=1.8
.ic q_59_81=0
.ic qb_59_81=1.8
.ic q_60_81=0
.ic qb_60_81=1.8
.ic q_61_81=0
.ic qb_61_81=1.8
.ic q_62_81=0
.ic qb_62_81=1.8
.ic q_63_81=0
.ic qb_63_81=1.8
.ic q_64_81=0
.ic qb_64_81=1.8
.ic q_65_81=0
.ic qb_65_81=1.8
.ic q_66_81=0
.ic qb_66_81=1.8
.ic q_67_81=0
.ic qb_67_81=1.8
.ic q_68_81=0
.ic qb_68_81=1.8
.ic q_69_81=0
.ic qb_69_81=1.8
.ic q_70_81=0
.ic qb_70_81=1.8
.ic q_71_81=0
.ic qb_71_81=1.8
.ic q_72_81=0
.ic qb_72_81=1.8
.ic q_73_81=0
.ic qb_73_81=1.8
.ic q_74_81=0
.ic qb_74_81=1.8
.ic q_75_81=0
.ic qb_75_81=1.8
.ic q_76_81=0
.ic qb_76_81=1.8
.ic q_77_81=0
.ic qb_77_81=1.8
.ic q_78_81=0
.ic qb_78_81=1.8
.ic q_79_81=0
.ic qb_79_81=1.8
.ic q_80_81=0
.ic qb_80_81=1.8
.ic q_81_81=0
.ic qb_81_81=1.8
.ic q_82_81=0
.ic qb_82_81=1.8
.ic q_83_81=0
.ic qb_83_81=1.8
.ic q_84_81=0
.ic qb_84_81=1.8
.ic q_85_81=0
.ic qb_85_81=1.8
.ic q_86_81=0
.ic qb_86_81=1.8
.ic q_87_81=0
.ic qb_87_81=1.8
.ic q_88_81=0
.ic qb_88_81=1.8
.ic q_89_81=0
.ic qb_89_81=1.8
.ic q_90_81=0
.ic qb_90_81=1.8
.ic q_91_81=0
.ic qb_91_81=1.8
.ic q_92_81=0
.ic qb_92_81=1.8
.ic q_93_81=0
.ic qb_93_81=1.8
.ic q_94_81=0
.ic qb_94_81=1.8
.ic q_95_81=0
.ic qb_95_81=1.8
.ic q_96_81=0
.ic qb_96_81=1.8
.ic q_97_81=0
.ic qb_97_81=1.8
.ic q_98_81=0
.ic qb_98_81=1.8
.ic q_99_81=0
.ic qb_99_81=1.8
.ic q_0_82=0
.ic qb_0_82=1.8
.ic q_1_82=0
.ic qb_1_82=1.8
.ic q_2_82=0
.ic qb_2_82=1.8
.ic q_3_82=0
.ic qb_3_82=1.8
.ic q_4_82=0
.ic qb_4_82=1.8
.ic q_5_82=0
.ic qb_5_82=1.8
.ic q_6_82=0
.ic qb_6_82=1.8
.ic q_7_82=0
.ic qb_7_82=1.8
.ic q_8_82=0
.ic qb_8_82=1.8
.ic q_9_82=0
.ic qb_9_82=1.8
.ic q_10_82=0
.ic qb_10_82=1.8
.ic q_11_82=0
.ic qb_11_82=1.8
.ic q_12_82=0
.ic qb_12_82=1.8
.ic q_13_82=0
.ic qb_13_82=1.8
.ic q_14_82=0
.ic qb_14_82=1.8
.ic q_15_82=0
.ic qb_15_82=1.8
.ic q_16_82=0
.ic qb_16_82=1.8
.ic q_17_82=0
.ic qb_17_82=1.8
.ic q_18_82=0
.ic qb_18_82=1.8
.ic q_19_82=0
.ic qb_19_82=1.8
.ic q_20_82=0
.ic qb_20_82=1.8
.ic q_21_82=0
.ic qb_21_82=1.8
.ic q_22_82=0
.ic qb_22_82=1.8
.ic q_23_82=0
.ic qb_23_82=1.8
.ic q_24_82=0
.ic qb_24_82=1.8
.ic q_25_82=0
.ic qb_25_82=1.8
.ic q_26_82=0
.ic qb_26_82=1.8
.ic q_27_82=0
.ic qb_27_82=1.8
.ic q_28_82=0
.ic qb_28_82=1.8
.ic q_29_82=0
.ic qb_29_82=1.8
.ic q_30_82=0
.ic qb_30_82=1.8
.ic q_31_82=0
.ic qb_31_82=1.8
.ic q_32_82=0
.ic qb_32_82=1.8
.ic q_33_82=0
.ic qb_33_82=1.8
.ic q_34_82=0
.ic qb_34_82=1.8
.ic q_35_82=0
.ic qb_35_82=1.8
.ic q_36_82=0
.ic qb_36_82=1.8
.ic q_37_82=0
.ic qb_37_82=1.8
.ic q_38_82=0
.ic qb_38_82=1.8
.ic q_39_82=0
.ic qb_39_82=1.8
.ic q_40_82=0
.ic qb_40_82=1.8
.ic q_41_82=0
.ic qb_41_82=1.8
.ic q_42_82=0
.ic qb_42_82=1.8
.ic q_43_82=0
.ic qb_43_82=1.8
.ic q_44_82=0
.ic qb_44_82=1.8
.ic q_45_82=0
.ic qb_45_82=1.8
.ic q_46_82=0
.ic qb_46_82=1.8
.ic q_47_82=0
.ic qb_47_82=1.8
.ic q_48_82=0
.ic qb_48_82=1.8
.ic q_49_82=0
.ic qb_49_82=1.8
.ic q_50_82=0
.ic qb_50_82=1.8
.ic q_51_82=0
.ic qb_51_82=1.8
.ic q_52_82=0
.ic qb_52_82=1.8
.ic q_53_82=0
.ic qb_53_82=1.8
.ic q_54_82=0
.ic qb_54_82=1.8
.ic q_55_82=0
.ic qb_55_82=1.8
.ic q_56_82=0
.ic qb_56_82=1.8
.ic q_57_82=0
.ic qb_57_82=1.8
.ic q_58_82=0
.ic qb_58_82=1.8
.ic q_59_82=0
.ic qb_59_82=1.8
.ic q_60_82=0
.ic qb_60_82=1.8
.ic q_61_82=0
.ic qb_61_82=1.8
.ic q_62_82=0
.ic qb_62_82=1.8
.ic q_63_82=0
.ic qb_63_82=1.8
.ic q_64_82=0
.ic qb_64_82=1.8
.ic q_65_82=0
.ic qb_65_82=1.8
.ic q_66_82=0
.ic qb_66_82=1.8
.ic q_67_82=0
.ic qb_67_82=1.8
.ic q_68_82=0
.ic qb_68_82=1.8
.ic q_69_82=0
.ic qb_69_82=1.8
.ic q_70_82=0
.ic qb_70_82=1.8
.ic q_71_82=0
.ic qb_71_82=1.8
.ic q_72_82=0
.ic qb_72_82=1.8
.ic q_73_82=0
.ic qb_73_82=1.8
.ic q_74_82=0
.ic qb_74_82=1.8
.ic q_75_82=0
.ic qb_75_82=1.8
.ic q_76_82=0
.ic qb_76_82=1.8
.ic q_77_82=0
.ic qb_77_82=1.8
.ic q_78_82=0
.ic qb_78_82=1.8
.ic q_79_82=0
.ic qb_79_82=1.8
.ic q_80_82=0
.ic qb_80_82=1.8
.ic q_81_82=0
.ic qb_81_82=1.8
.ic q_82_82=0
.ic qb_82_82=1.8
.ic q_83_82=0
.ic qb_83_82=1.8
.ic q_84_82=0
.ic qb_84_82=1.8
.ic q_85_82=0
.ic qb_85_82=1.8
.ic q_86_82=0
.ic qb_86_82=1.8
.ic q_87_82=0
.ic qb_87_82=1.8
.ic q_88_82=0
.ic qb_88_82=1.8
.ic q_89_82=0
.ic qb_89_82=1.8
.ic q_90_82=0
.ic qb_90_82=1.8
.ic q_91_82=0
.ic qb_91_82=1.8
.ic q_92_82=0
.ic qb_92_82=1.8
.ic q_93_82=0
.ic qb_93_82=1.8
.ic q_94_82=0
.ic qb_94_82=1.8
.ic q_95_82=0
.ic qb_95_82=1.8
.ic q_96_82=0
.ic qb_96_82=1.8
.ic q_97_82=0
.ic qb_97_82=1.8
.ic q_98_82=0
.ic qb_98_82=1.8
.ic q_99_82=0
.ic qb_99_82=1.8
.ic q_0_83=0
.ic qb_0_83=1.8
.ic q_1_83=0
.ic qb_1_83=1.8
.ic q_2_83=0
.ic qb_2_83=1.8
.ic q_3_83=0
.ic qb_3_83=1.8
.ic q_4_83=0
.ic qb_4_83=1.8
.ic q_5_83=0
.ic qb_5_83=1.8
.ic q_6_83=0
.ic qb_6_83=1.8
.ic q_7_83=0
.ic qb_7_83=1.8
.ic q_8_83=0
.ic qb_8_83=1.8
.ic q_9_83=0
.ic qb_9_83=1.8
.ic q_10_83=0
.ic qb_10_83=1.8
.ic q_11_83=0
.ic qb_11_83=1.8
.ic q_12_83=0
.ic qb_12_83=1.8
.ic q_13_83=0
.ic qb_13_83=1.8
.ic q_14_83=0
.ic qb_14_83=1.8
.ic q_15_83=0
.ic qb_15_83=1.8
.ic q_16_83=0
.ic qb_16_83=1.8
.ic q_17_83=0
.ic qb_17_83=1.8
.ic q_18_83=0
.ic qb_18_83=1.8
.ic q_19_83=0
.ic qb_19_83=1.8
.ic q_20_83=0
.ic qb_20_83=1.8
.ic q_21_83=0
.ic qb_21_83=1.8
.ic q_22_83=0
.ic qb_22_83=1.8
.ic q_23_83=0
.ic qb_23_83=1.8
.ic q_24_83=0
.ic qb_24_83=1.8
.ic q_25_83=0
.ic qb_25_83=1.8
.ic q_26_83=0
.ic qb_26_83=1.8
.ic q_27_83=0
.ic qb_27_83=1.8
.ic q_28_83=0
.ic qb_28_83=1.8
.ic q_29_83=0
.ic qb_29_83=1.8
.ic q_30_83=0
.ic qb_30_83=1.8
.ic q_31_83=0
.ic qb_31_83=1.8
.ic q_32_83=0
.ic qb_32_83=1.8
.ic q_33_83=0
.ic qb_33_83=1.8
.ic q_34_83=0
.ic qb_34_83=1.8
.ic q_35_83=0
.ic qb_35_83=1.8
.ic q_36_83=0
.ic qb_36_83=1.8
.ic q_37_83=0
.ic qb_37_83=1.8
.ic q_38_83=0
.ic qb_38_83=1.8
.ic q_39_83=0
.ic qb_39_83=1.8
.ic q_40_83=0
.ic qb_40_83=1.8
.ic q_41_83=0
.ic qb_41_83=1.8
.ic q_42_83=0
.ic qb_42_83=1.8
.ic q_43_83=0
.ic qb_43_83=1.8
.ic q_44_83=0
.ic qb_44_83=1.8
.ic q_45_83=0
.ic qb_45_83=1.8
.ic q_46_83=0
.ic qb_46_83=1.8
.ic q_47_83=0
.ic qb_47_83=1.8
.ic q_48_83=0
.ic qb_48_83=1.8
.ic q_49_83=0
.ic qb_49_83=1.8
.ic q_50_83=0
.ic qb_50_83=1.8
.ic q_51_83=0
.ic qb_51_83=1.8
.ic q_52_83=0
.ic qb_52_83=1.8
.ic q_53_83=0
.ic qb_53_83=1.8
.ic q_54_83=0
.ic qb_54_83=1.8
.ic q_55_83=0
.ic qb_55_83=1.8
.ic q_56_83=0
.ic qb_56_83=1.8
.ic q_57_83=0
.ic qb_57_83=1.8
.ic q_58_83=0
.ic qb_58_83=1.8
.ic q_59_83=0
.ic qb_59_83=1.8
.ic q_60_83=0
.ic qb_60_83=1.8
.ic q_61_83=0
.ic qb_61_83=1.8
.ic q_62_83=0
.ic qb_62_83=1.8
.ic q_63_83=0
.ic qb_63_83=1.8
.ic q_64_83=0
.ic qb_64_83=1.8
.ic q_65_83=0
.ic qb_65_83=1.8
.ic q_66_83=0
.ic qb_66_83=1.8
.ic q_67_83=0
.ic qb_67_83=1.8
.ic q_68_83=0
.ic qb_68_83=1.8
.ic q_69_83=0
.ic qb_69_83=1.8
.ic q_70_83=0
.ic qb_70_83=1.8
.ic q_71_83=0
.ic qb_71_83=1.8
.ic q_72_83=0
.ic qb_72_83=1.8
.ic q_73_83=0
.ic qb_73_83=1.8
.ic q_74_83=0
.ic qb_74_83=1.8
.ic q_75_83=0
.ic qb_75_83=1.8
.ic q_76_83=0
.ic qb_76_83=1.8
.ic q_77_83=0
.ic qb_77_83=1.8
.ic q_78_83=0
.ic qb_78_83=1.8
.ic q_79_83=0
.ic qb_79_83=1.8
.ic q_80_83=0
.ic qb_80_83=1.8
.ic q_81_83=0
.ic qb_81_83=1.8
.ic q_82_83=0
.ic qb_82_83=1.8
.ic q_83_83=0
.ic qb_83_83=1.8
.ic q_84_83=0
.ic qb_84_83=1.8
.ic q_85_83=0
.ic qb_85_83=1.8
.ic q_86_83=0
.ic qb_86_83=1.8
.ic q_87_83=0
.ic qb_87_83=1.8
.ic q_88_83=0
.ic qb_88_83=1.8
.ic q_89_83=0
.ic qb_89_83=1.8
.ic q_90_83=0
.ic qb_90_83=1.8
.ic q_91_83=0
.ic qb_91_83=1.8
.ic q_92_83=0
.ic qb_92_83=1.8
.ic q_93_83=0
.ic qb_93_83=1.8
.ic q_94_83=0
.ic qb_94_83=1.8
.ic q_95_83=0
.ic qb_95_83=1.8
.ic q_96_83=0
.ic qb_96_83=1.8
.ic q_97_83=0
.ic qb_97_83=1.8
.ic q_98_83=0
.ic qb_98_83=1.8
.ic q_99_83=0
.ic qb_99_83=1.8
.ic q_0_84=0
.ic qb_0_84=1.8
.ic q_1_84=0
.ic qb_1_84=1.8
.ic q_2_84=0
.ic qb_2_84=1.8
.ic q_3_84=0
.ic qb_3_84=1.8
.ic q_4_84=0
.ic qb_4_84=1.8
.ic q_5_84=0
.ic qb_5_84=1.8
.ic q_6_84=0
.ic qb_6_84=1.8
.ic q_7_84=0
.ic qb_7_84=1.8
.ic q_8_84=0
.ic qb_8_84=1.8
.ic q_9_84=0
.ic qb_9_84=1.8
.ic q_10_84=0
.ic qb_10_84=1.8
.ic q_11_84=0
.ic qb_11_84=1.8
.ic q_12_84=0
.ic qb_12_84=1.8
.ic q_13_84=0
.ic qb_13_84=1.8
.ic q_14_84=0
.ic qb_14_84=1.8
.ic q_15_84=0
.ic qb_15_84=1.8
.ic q_16_84=0
.ic qb_16_84=1.8
.ic q_17_84=0
.ic qb_17_84=1.8
.ic q_18_84=0
.ic qb_18_84=1.8
.ic q_19_84=0
.ic qb_19_84=1.8
.ic q_20_84=0
.ic qb_20_84=1.8
.ic q_21_84=0
.ic qb_21_84=1.8
.ic q_22_84=0
.ic qb_22_84=1.8
.ic q_23_84=0
.ic qb_23_84=1.8
.ic q_24_84=0
.ic qb_24_84=1.8
.ic q_25_84=0
.ic qb_25_84=1.8
.ic q_26_84=0
.ic qb_26_84=1.8
.ic q_27_84=0
.ic qb_27_84=1.8
.ic q_28_84=0
.ic qb_28_84=1.8
.ic q_29_84=0
.ic qb_29_84=1.8
.ic q_30_84=0
.ic qb_30_84=1.8
.ic q_31_84=0
.ic qb_31_84=1.8
.ic q_32_84=0
.ic qb_32_84=1.8
.ic q_33_84=0
.ic qb_33_84=1.8
.ic q_34_84=0
.ic qb_34_84=1.8
.ic q_35_84=0
.ic qb_35_84=1.8
.ic q_36_84=0
.ic qb_36_84=1.8
.ic q_37_84=0
.ic qb_37_84=1.8
.ic q_38_84=0
.ic qb_38_84=1.8
.ic q_39_84=0
.ic qb_39_84=1.8
.ic q_40_84=0
.ic qb_40_84=1.8
.ic q_41_84=0
.ic qb_41_84=1.8
.ic q_42_84=0
.ic qb_42_84=1.8
.ic q_43_84=0
.ic qb_43_84=1.8
.ic q_44_84=0
.ic qb_44_84=1.8
.ic q_45_84=0
.ic qb_45_84=1.8
.ic q_46_84=0
.ic qb_46_84=1.8
.ic q_47_84=0
.ic qb_47_84=1.8
.ic q_48_84=0
.ic qb_48_84=1.8
.ic q_49_84=0
.ic qb_49_84=1.8
.ic q_50_84=0
.ic qb_50_84=1.8
.ic q_51_84=0
.ic qb_51_84=1.8
.ic q_52_84=0
.ic qb_52_84=1.8
.ic q_53_84=0
.ic qb_53_84=1.8
.ic q_54_84=0
.ic qb_54_84=1.8
.ic q_55_84=0
.ic qb_55_84=1.8
.ic q_56_84=0
.ic qb_56_84=1.8
.ic q_57_84=0
.ic qb_57_84=1.8
.ic q_58_84=0
.ic qb_58_84=1.8
.ic q_59_84=0
.ic qb_59_84=1.8
.ic q_60_84=0
.ic qb_60_84=1.8
.ic q_61_84=0
.ic qb_61_84=1.8
.ic q_62_84=0
.ic qb_62_84=1.8
.ic q_63_84=0
.ic qb_63_84=1.8
.ic q_64_84=0
.ic qb_64_84=1.8
.ic q_65_84=0
.ic qb_65_84=1.8
.ic q_66_84=0
.ic qb_66_84=1.8
.ic q_67_84=0
.ic qb_67_84=1.8
.ic q_68_84=0
.ic qb_68_84=1.8
.ic q_69_84=0
.ic qb_69_84=1.8
.ic q_70_84=0
.ic qb_70_84=1.8
.ic q_71_84=0
.ic qb_71_84=1.8
.ic q_72_84=0
.ic qb_72_84=1.8
.ic q_73_84=0
.ic qb_73_84=1.8
.ic q_74_84=0
.ic qb_74_84=1.8
.ic q_75_84=0
.ic qb_75_84=1.8
.ic q_76_84=0
.ic qb_76_84=1.8
.ic q_77_84=0
.ic qb_77_84=1.8
.ic q_78_84=0
.ic qb_78_84=1.8
.ic q_79_84=0
.ic qb_79_84=1.8
.ic q_80_84=0
.ic qb_80_84=1.8
.ic q_81_84=0
.ic qb_81_84=1.8
.ic q_82_84=0
.ic qb_82_84=1.8
.ic q_83_84=0
.ic qb_83_84=1.8
.ic q_84_84=0
.ic qb_84_84=1.8
.ic q_85_84=0
.ic qb_85_84=1.8
.ic q_86_84=0
.ic qb_86_84=1.8
.ic q_87_84=0
.ic qb_87_84=1.8
.ic q_88_84=0
.ic qb_88_84=1.8
.ic q_89_84=0
.ic qb_89_84=1.8
.ic q_90_84=0
.ic qb_90_84=1.8
.ic q_91_84=0
.ic qb_91_84=1.8
.ic q_92_84=0
.ic qb_92_84=1.8
.ic q_93_84=0
.ic qb_93_84=1.8
.ic q_94_84=0
.ic qb_94_84=1.8
.ic q_95_84=0
.ic qb_95_84=1.8
.ic q_96_84=0
.ic qb_96_84=1.8
.ic q_97_84=0
.ic qb_97_84=1.8
.ic q_98_84=0
.ic qb_98_84=1.8
.ic q_99_84=0
.ic qb_99_84=1.8
.ic q_0_85=0
.ic qb_0_85=1.8
.ic q_1_85=0
.ic qb_1_85=1.8
.ic q_2_85=0
.ic qb_2_85=1.8
.ic q_3_85=0
.ic qb_3_85=1.8
.ic q_4_85=0
.ic qb_4_85=1.8
.ic q_5_85=0
.ic qb_5_85=1.8
.ic q_6_85=0
.ic qb_6_85=1.8
.ic q_7_85=0
.ic qb_7_85=1.8
.ic q_8_85=0
.ic qb_8_85=1.8
.ic q_9_85=0
.ic qb_9_85=1.8
.ic q_10_85=0
.ic qb_10_85=1.8
.ic q_11_85=0
.ic qb_11_85=1.8
.ic q_12_85=0
.ic qb_12_85=1.8
.ic q_13_85=0
.ic qb_13_85=1.8
.ic q_14_85=0
.ic qb_14_85=1.8
.ic q_15_85=0
.ic qb_15_85=1.8
.ic q_16_85=0
.ic qb_16_85=1.8
.ic q_17_85=0
.ic qb_17_85=1.8
.ic q_18_85=0
.ic qb_18_85=1.8
.ic q_19_85=0
.ic qb_19_85=1.8
.ic q_20_85=0
.ic qb_20_85=1.8
.ic q_21_85=0
.ic qb_21_85=1.8
.ic q_22_85=0
.ic qb_22_85=1.8
.ic q_23_85=0
.ic qb_23_85=1.8
.ic q_24_85=0
.ic qb_24_85=1.8
.ic q_25_85=0
.ic qb_25_85=1.8
.ic q_26_85=0
.ic qb_26_85=1.8
.ic q_27_85=0
.ic qb_27_85=1.8
.ic q_28_85=0
.ic qb_28_85=1.8
.ic q_29_85=0
.ic qb_29_85=1.8
.ic q_30_85=0
.ic qb_30_85=1.8
.ic q_31_85=0
.ic qb_31_85=1.8
.ic q_32_85=0
.ic qb_32_85=1.8
.ic q_33_85=0
.ic qb_33_85=1.8
.ic q_34_85=0
.ic qb_34_85=1.8
.ic q_35_85=0
.ic qb_35_85=1.8
.ic q_36_85=0
.ic qb_36_85=1.8
.ic q_37_85=0
.ic qb_37_85=1.8
.ic q_38_85=0
.ic qb_38_85=1.8
.ic q_39_85=0
.ic qb_39_85=1.8
.ic q_40_85=0
.ic qb_40_85=1.8
.ic q_41_85=0
.ic qb_41_85=1.8
.ic q_42_85=0
.ic qb_42_85=1.8
.ic q_43_85=0
.ic qb_43_85=1.8
.ic q_44_85=0
.ic qb_44_85=1.8
.ic q_45_85=0
.ic qb_45_85=1.8
.ic q_46_85=0
.ic qb_46_85=1.8
.ic q_47_85=0
.ic qb_47_85=1.8
.ic q_48_85=0
.ic qb_48_85=1.8
.ic q_49_85=0
.ic qb_49_85=1.8
.ic q_50_85=0
.ic qb_50_85=1.8
.ic q_51_85=0
.ic qb_51_85=1.8
.ic q_52_85=0
.ic qb_52_85=1.8
.ic q_53_85=0
.ic qb_53_85=1.8
.ic q_54_85=0
.ic qb_54_85=1.8
.ic q_55_85=0
.ic qb_55_85=1.8
.ic q_56_85=0
.ic qb_56_85=1.8
.ic q_57_85=0
.ic qb_57_85=1.8
.ic q_58_85=0
.ic qb_58_85=1.8
.ic q_59_85=0
.ic qb_59_85=1.8
.ic q_60_85=0
.ic qb_60_85=1.8
.ic q_61_85=0
.ic qb_61_85=1.8
.ic q_62_85=0
.ic qb_62_85=1.8
.ic q_63_85=0
.ic qb_63_85=1.8
.ic q_64_85=0
.ic qb_64_85=1.8
.ic q_65_85=0
.ic qb_65_85=1.8
.ic q_66_85=0
.ic qb_66_85=1.8
.ic q_67_85=0
.ic qb_67_85=1.8
.ic q_68_85=0
.ic qb_68_85=1.8
.ic q_69_85=0
.ic qb_69_85=1.8
.ic q_70_85=0
.ic qb_70_85=1.8
.ic q_71_85=0
.ic qb_71_85=1.8
.ic q_72_85=0
.ic qb_72_85=1.8
.ic q_73_85=0
.ic qb_73_85=1.8
.ic q_74_85=0
.ic qb_74_85=1.8
.ic q_75_85=0
.ic qb_75_85=1.8
.ic q_76_85=0
.ic qb_76_85=1.8
.ic q_77_85=0
.ic qb_77_85=1.8
.ic q_78_85=0
.ic qb_78_85=1.8
.ic q_79_85=0
.ic qb_79_85=1.8
.ic q_80_85=0
.ic qb_80_85=1.8
.ic q_81_85=0
.ic qb_81_85=1.8
.ic q_82_85=0
.ic qb_82_85=1.8
.ic q_83_85=0
.ic qb_83_85=1.8
.ic q_84_85=0
.ic qb_84_85=1.8
.ic q_85_85=0
.ic qb_85_85=1.8
.ic q_86_85=0
.ic qb_86_85=1.8
.ic q_87_85=0
.ic qb_87_85=1.8
.ic q_88_85=0
.ic qb_88_85=1.8
.ic q_89_85=0
.ic qb_89_85=1.8
.ic q_90_85=0
.ic qb_90_85=1.8
.ic q_91_85=0
.ic qb_91_85=1.8
.ic q_92_85=0
.ic qb_92_85=1.8
.ic q_93_85=0
.ic qb_93_85=1.8
.ic q_94_85=0
.ic qb_94_85=1.8
.ic q_95_85=0
.ic qb_95_85=1.8
.ic q_96_85=0
.ic qb_96_85=1.8
.ic q_97_85=0
.ic qb_97_85=1.8
.ic q_98_85=0
.ic qb_98_85=1.8
.ic q_99_85=0
.ic qb_99_85=1.8
.ic q_0_86=0
.ic qb_0_86=1.8
.ic q_1_86=0
.ic qb_1_86=1.8
.ic q_2_86=0
.ic qb_2_86=1.8
.ic q_3_86=0
.ic qb_3_86=1.8
.ic q_4_86=0
.ic qb_4_86=1.8
.ic q_5_86=0
.ic qb_5_86=1.8
.ic q_6_86=0
.ic qb_6_86=1.8
.ic q_7_86=0
.ic qb_7_86=1.8
.ic q_8_86=0
.ic qb_8_86=1.8
.ic q_9_86=0
.ic qb_9_86=1.8
.ic q_10_86=0
.ic qb_10_86=1.8
.ic q_11_86=0
.ic qb_11_86=1.8
.ic q_12_86=0
.ic qb_12_86=1.8
.ic q_13_86=0
.ic qb_13_86=1.8
.ic q_14_86=0
.ic qb_14_86=1.8
.ic q_15_86=0
.ic qb_15_86=1.8
.ic q_16_86=0
.ic qb_16_86=1.8
.ic q_17_86=0
.ic qb_17_86=1.8
.ic q_18_86=0
.ic qb_18_86=1.8
.ic q_19_86=0
.ic qb_19_86=1.8
.ic q_20_86=0
.ic qb_20_86=1.8
.ic q_21_86=0
.ic qb_21_86=1.8
.ic q_22_86=0
.ic qb_22_86=1.8
.ic q_23_86=0
.ic qb_23_86=1.8
.ic q_24_86=0
.ic qb_24_86=1.8
.ic q_25_86=0
.ic qb_25_86=1.8
.ic q_26_86=0
.ic qb_26_86=1.8
.ic q_27_86=0
.ic qb_27_86=1.8
.ic q_28_86=0
.ic qb_28_86=1.8
.ic q_29_86=0
.ic qb_29_86=1.8
.ic q_30_86=0
.ic qb_30_86=1.8
.ic q_31_86=0
.ic qb_31_86=1.8
.ic q_32_86=0
.ic qb_32_86=1.8
.ic q_33_86=0
.ic qb_33_86=1.8
.ic q_34_86=0
.ic qb_34_86=1.8
.ic q_35_86=0
.ic qb_35_86=1.8
.ic q_36_86=0
.ic qb_36_86=1.8
.ic q_37_86=0
.ic qb_37_86=1.8
.ic q_38_86=0
.ic qb_38_86=1.8
.ic q_39_86=0
.ic qb_39_86=1.8
.ic q_40_86=0
.ic qb_40_86=1.8
.ic q_41_86=0
.ic qb_41_86=1.8
.ic q_42_86=0
.ic qb_42_86=1.8
.ic q_43_86=0
.ic qb_43_86=1.8
.ic q_44_86=0
.ic qb_44_86=1.8
.ic q_45_86=0
.ic qb_45_86=1.8
.ic q_46_86=0
.ic qb_46_86=1.8
.ic q_47_86=0
.ic qb_47_86=1.8
.ic q_48_86=0
.ic qb_48_86=1.8
.ic q_49_86=0
.ic qb_49_86=1.8
.ic q_50_86=0
.ic qb_50_86=1.8
.ic q_51_86=0
.ic qb_51_86=1.8
.ic q_52_86=0
.ic qb_52_86=1.8
.ic q_53_86=0
.ic qb_53_86=1.8
.ic q_54_86=0
.ic qb_54_86=1.8
.ic q_55_86=0
.ic qb_55_86=1.8
.ic q_56_86=0
.ic qb_56_86=1.8
.ic q_57_86=0
.ic qb_57_86=1.8
.ic q_58_86=0
.ic qb_58_86=1.8
.ic q_59_86=0
.ic qb_59_86=1.8
.ic q_60_86=0
.ic qb_60_86=1.8
.ic q_61_86=0
.ic qb_61_86=1.8
.ic q_62_86=0
.ic qb_62_86=1.8
.ic q_63_86=0
.ic qb_63_86=1.8
.ic q_64_86=0
.ic qb_64_86=1.8
.ic q_65_86=0
.ic qb_65_86=1.8
.ic q_66_86=0
.ic qb_66_86=1.8
.ic q_67_86=0
.ic qb_67_86=1.8
.ic q_68_86=0
.ic qb_68_86=1.8
.ic q_69_86=0
.ic qb_69_86=1.8
.ic q_70_86=0
.ic qb_70_86=1.8
.ic q_71_86=0
.ic qb_71_86=1.8
.ic q_72_86=0
.ic qb_72_86=1.8
.ic q_73_86=0
.ic qb_73_86=1.8
.ic q_74_86=0
.ic qb_74_86=1.8
.ic q_75_86=0
.ic qb_75_86=1.8
.ic q_76_86=0
.ic qb_76_86=1.8
.ic q_77_86=0
.ic qb_77_86=1.8
.ic q_78_86=0
.ic qb_78_86=1.8
.ic q_79_86=0
.ic qb_79_86=1.8
.ic q_80_86=0
.ic qb_80_86=1.8
.ic q_81_86=0
.ic qb_81_86=1.8
.ic q_82_86=0
.ic qb_82_86=1.8
.ic q_83_86=0
.ic qb_83_86=1.8
.ic q_84_86=0
.ic qb_84_86=1.8
.ic q_85_86=0
.ic qb_85_86=1.8
.ic q_86_86=0
.ic qb_86_86=1.8
.ic q_87_86=0
.ic qb_87_86=1.8
.ic q_88_86=0
.ic qb_88_86=1.8
.ic q_89_86=0
.ic qb_89_86=1.8
.ic q_90_86=0
.ic qb_90_86=1.8
.ic q_91_86=0
.ic qb_91_86=1.8
.ic q_92_86=0
.ic qb_92_86=1.8
.ic q_93_86=0
.ic qb_93_86=1.8
.ic q_94_86=0
.ic qb_94_86=1.8
.ic q_95_86=0
.ic qb_95_86=1.8
.ic q_96_86=0
.ic qb_96_86=1.8
.ic q_97_86=0
.ic qb_97_86=1.8
.ic q_98_86=0
.ic qb_98_86=1.8
.ic q_99_86=0
.ic qb_99_86=1.8
.ic q_0_87=0
.ic qb_0_87=1.8
.ic q_1_87=0
.ic qb_1_87=1.8
.ic q_2_87=0
.ic qb_2_87=1.8
.ic q_3_87=0
.ic qb_3_87=1.8
.ic q_4_87=0
.ic qb_4_87=1.8
.ic q_5_87=0
.ic qb_5_87=1.8
.ic q_6_87=0
.ic qb_6_87=1.8
.ic q_7_87=0
.ic qb_7_87=1.8
.ic q_8_87=0
.ic qb_8_87=1.8
.ic q_9_87=0
.ic qb_9_87=1.8
.ic q_10_87=0
.ic qb_10_87=1.8
.ic q_11_87=0
.ic qb_11_87=1.8
.ic q_12_87=0
.ic qb_12_87=1.8
.ic q_13_87=0
.ic qb_13_87=1.8
.ic q_14_87=0
.ic qb_14_87=1.8
.ic q_15_87=0
.ic qb_15_87=1.8
.ic q_16_87=0
.ic qb_16_87=1.8
.ic q_17_87=0
.ic qb_17_87=1.8
.ic q_18_87=0
.ic qb_18_87=1.8
.ic q_19_87=0
.ic qb_19_87=1.8
.ic q_20_87=0
.ic qb_20_87=1.8
.ic q_21_87=0
.ic qb_21_87=1.8
.ic q_22_87=0
.ic qb_22_87=1.8
.ic q_23_87=0
.ic qb_23_87=1.8
.ic q_24_87=0
.ic qb_24_87=1.8
.ic q_25_87=0
.ic qb_25_87=1.8
.ic q_26_87=0
.ic qb_26_87=1.8
.ic q_27_87=0
.ic qb_27_87=1.8
.ic q_28_87=0
.ic qb_28_87=1.8
.ic q_29_87=0
.ic qb_29_87=1.8
.ic q_30_87=0
.ic qb_30_87=1.8
.ic q_31_87=0
.ic qb_31_87=1.8
.ic q_32_87=0
.ic qb_32_87=1.8
.ic q_33_87=0
.ic qb_33_87=1.8
.ic q_34_87=0
.ic qb_34_87=1.8
.ic q_35_87=0
.ic qb_35_87=1.8
.ic q_36_87=0
.ic qb_36_87=1.8
.ic q_37_87=0
.ic qb_37_87=1.8
.ic q_38_87=0
.ic qb_38_87=1.8
.ic q_39_87=0
.ic qb_39_87=1.8
.ic q_40_87=0
.ic qb_40_87=1.8
.ic q_41_87=0
.ic qb_41_87=1.8
.ic q_42_87=0
.ic qb_42_87=1.8
.ic q_43_87=0
.ic qb_43_87=1.8
.ic q_44_87=0
.ic qb_44_87=1.8
.ic q_45_87=0
.ic qb_45_87=1.8
.ic q_46_87=0
.ic qb_46_87=1.8
.ic q_47_87=0
.ic qb_47_87=1.8
.ic q_48_87=0
.ic qb_48_87=1.8
.ic q_49_87=0
.ic qb_49_87=1.8
.ic q_50_87=0
.ic qb_50_87=1.8
.ic q_51_87=0
.ic qb_51_87=1.8
.ic q_52_87=0
.ic qb_52_87=1.8
.ic q_53_87=0
.ic qb_53_87=1.8
.ic q_54_87=0
.ic qb_54_87=1.8
.ic q_55_87=0
.ic qb_55_87=1.8
.ic q_56_87=0
.ic qb_56_87=1.8
.ic q_57_87=0
.ic qb_57_87=1.8
.ic q_58_87=0
.ic qb_58_87=1.8
.ic q_59_87=0
.ic qb_59_87=1.8
.ic q_60_87=0
.ic qb_60_87=1.8
.ic q_61_87=0
.ic qb_61_87=1.8
.ic q_62_87=0
.ic qb_62_87=1.8
.ic q_63_87=0
.ic qb_63_87=1.8
.ic q_64_87=0
.ic qb_64_87=1.8
.ic q_65_87=0
.ic qb_65_87=1.8
.ic q_66_87=0
.ic qb_66_87=1.8
.ic q_67_87=0
.ic qb_67_87=1.8
.ic q_68_87=0
.ic qb_68_87=1.8
.ic q_69_87=0
.ic qb_69_87=1.8
.ic q_70_87=0
.ic qb_70_87=1.8
.ic q_71_87=0
.ic qb_71_87=1.8
.ic q_72_87=0
.ic qb_72_87=1.8
.ic q_73_87=0
.ic qb_73_87=1.8
.ic q_74_87=0
.ic qb_74_87=1.8
.ic q_75_87=0
.ic qb_75_87=1.8
.ic q_76_87=0
.ic qb_76_87=1.8
.ic q_77_87=0
.ic qb_77_87=1.8
.ic q_78_87=0
.ic qb_78_87=1.8
.ic q_79_87=0
.ic qb_79_87=1.8
.ic q_80_87=0
.ic qb_80_87=1.8
.ic q_81_87=0
.ic qb_81_87=1.8
.ic q_82_87=0
.ic qb_82_87=1.8
.ic q_83_87=0
.ic qb_83_87=1.8
.ic q_84_87=0
.ic qb_84_87=1.8
.ic q_85_87=0
.ic qb_85_87=1.8
.ic q_86_87=0
.ic qb_86_87=1.8
.ic q_87_87=0
.ic qb_87_87=1.8
.ic q_88_87=0
.ic qb_88_87=1.8
.ic q_89_87=0
.ic qb_89_87=1.8
.ic q_90_87=0
.ic qb_90_87=1.8
.ic q_91_87=0
.ic qb_91_87=1.8
.ic q_92_87=0
.ic qb_92_87=1.8
.ic q_93_87=0
.ic qb_93_87=1.8
.ic q_94_87=0
.ic qb_94_87=1.8
.ic q_95_87=0
.ic qb_95_87=1.8
.ic q_96_87=0
.ic qb_96_87=1.8
.ic q_97_87=0
.ic qb_97_87=1.8
.ic q_98_87=0
.ic qb_98_87=1.8
.ic q_99_87=0
.ic qb_99_87=1.8
.ic q_0_88=0
.ic qb_0_88=1.8
.ic q_1_88=0
.ic qb_1_88=1.8
.ic q_2_88=0
.ic qb_2_88=1.8
.ic q_3_88=0
.ic qb_3_88=1.8
.ic q_4_88=0
.ic qb_4_88=1.8
.ic q_5_88=0
.ic qb_5_88=1.8
.ic q_6_88=0
.ic qb_6_88=1.8
.ic q_7_88=0
.ic qb_7_88=1.8
.ic q_8_88=0
.ic qb_8_88=1.8
.ic q_9_88=0
.ic qb_9_88=1.8
.ic q_10_88=0
.ic qb_10_88=1.8
.ic q_11_88=0
.ic qb_11_88=1.8
.ic q_12_88=0
.ic qb_12_88=1.8
.ic q_13_88=0
.ic qb_13_88=1.8
.ic q_14_88=0
.ic qb_14_88=1.8
.ic q_15_88=0
.ic qb_15_88=1.8
.ic q_16_88=0
.ic qb_16_88=1.8
.ic q_17_88=0
.ic qb_17_88=1.8
.ic q_18_88=0
.ic qb_18_88=1.8
.ic q_19_88=0
.ic qb_19_88=1.8
.ic q_20_88=0
.ic qb_20_88=1.8
.ic q_21_88=0
.ic qb_21_88=1.8
.ic q_22_88=0
.ic qb_22_88=1.8
.ic q_23_88=0
.ic qb_23_88=1.8
.ic q_24_88=0
.ic qb_24_88=1.8
.ic q_25_88=0
.ic qb_25_88=1.8
.ic q_26_88=0
.ic qb_26_88=1.8
.ic q_27_88=0
.ic qb_27_88=1.8
.ic q_28_88=0
.ic qb_28_88=1.8
.ic q_29_88=0
.ic qb_29_88=1.8
.ic q_30_88=0
.ic qb_30_88=1.8
.ic q_31_88=0
.ic qb_31_88=1.8
.ic q_32_88=0
.ic qb_32_88=1.8
.ic q_33_88=0
.ic qb_33_88=1.8
.ic q_34_88=0
.ic qb_34_88=1.8
.ic q_35_88=0
.ic qb_35_88=1.8
.ic q_36_88=0
.ic qb_36_88=1.8
.ic q_37_88=0
.ic qb_37_88=1.8
.ic q_38_88=0
.ic qb_38_88=1.8
.ic q_39_88=0
.ic qb_39_88=1.8
.ic q_40_88=0
.ic qb_40_88=1.8
.ic q_41_88=0
.ic qb_41_88=1.8
.ic q_42_88=0
.ic qb_42_88=1.8
.ic q_43_88=0
.ic qb_43_88=1.8
.ic q_44_88=0
.ic qb_44_88=1.8
.ic q_45_88=0
.ic qb_45_88=1.8
.ic q_46_88=0
.ic qb_46_88=1.8
.ic q_47_88=0
.ic qb_47_88=1.8
.ic q_48_88=0
.ic qb_48_88=1.8
.ic q_49_88=0
.ic qb_49_88=1.8
.ic q_50_88=0
.ic qb_50_88=1.8
.ic q_51_88=0
.ic qb_51_88=1.8
.ic q_52_88=0
.ic qb_52_88=1.8
.ic q_53_88=0
.ic qb_53_88=1.8
.ic q_54_88=0
.ic qb_54_88=1.8
.ic q_55_88=0
.ic qb_55_88=1.8
.ic q_56_88=0
.ic qb_56_88=1.8
.ic q_57_88=0
.ic qb_57_88=1.8
.ic q_58_88=0
.ic qb_58_88=1.8
.ic q_59_88=0
.ic qb_59_88=1.8
.ic q_60_88=0
.ic qb_60_88=1.8
.ic q_61_88=0
.ic qb_61_88=1.8
.ic q_62_88=0
.ic qb_62_88=1.8
.ic q_63_88=0
.ic qb_63_88=1.8
.ic q_64_88=0
.ic qb_64_88=1.8
.ic q_65_88=0
.ic qb_65_88=1.8
.ic q_66_88=0
.ic qb_66_88=1.8
.ic q_67_88=0
.ic qb_67_88=1.8
.ic q_68_88=0
.ic qb_68_88=1.8
.ic q_69_88=0
.ic qb_69_88=1.8
.ic q_70_88=0
.ic qb_70_88=1.8
.ic q_71_88=0
.ic qb_71_88=1.8
.ic q_72_88=0
.ic qb_72_88=1.8
.ic q_73_88=0
.ic qb_73_88=1.8
.ic q_74_88=0
.ic qb_74_88=1.8
.ic q_75_88=0
.ic qb_75_88=1.8
.ic q_76_88=0
.ic qb_76_88=1.8
.ic q_77_88=0
.ic qb_77_88=1.8
.ic q_78_88=0
.ic qb_78_88=1.8
.ic q_79_88=0
.ic qb_79_88=1.8
.ic q_80_88=0
.ic qb_80_88=1.8
.ic q_81_88=0
.ic qb_81_88=1.8
.ic q_82_88=0
.ic qb_82_88=1.8
.ic q_83_88=0
.ic qb_83_88=1.8
.ic q_84_88=0
.ic qb_84_88=1.8
.ic q_85_88=0
.ic qb_85_88=1.8
.ic q_86_88=0
.ic qb_86_88=1.8
.ic q_87_88=0
.ic qb_87_88=1.8
.ic q_88_88=0
.ic qb_88_88=1.8
.ic q_89_88=0
.ic qb_89_88=1.8
.ic q_90_88=0
.ic qb_90_88=1.8
.ic q_91_88=0
.ic qb_91_88=1.8
.ic q_92_88=0
.ic qb_92_88=1.8
.ic q_93_88=0
.ic qb_93_88=1.8
.ic q_94_88=0
.ic qb_94_88=1.8
.ic q_95_88=0
.ic qb_95_88=1.8
.ic q_96_88=0
.ic qb_96_88=1.8
.ic q_97_88=0
.ic qb_97_88=1.8
.ic q_98_88=0
.ic qb_98_88=1.8
.ic q_99_88=0
.ic qb_99_88=1.8
.ic q_0_89=0
.ic qb_0_89=1.8
.ic q_1_89=0
.ic qb_1_89=1.8
.ic q_2_89=0
.ic qb_2_89=1.8
.ic q_3_89=0
.ic qb_3_89=1.8
.ic q_4_89=0
.ic qb_4_89=1.8
.ic q_5_89=0
.ic qb_5_89=1.8
.ic q_6_89=0
.ic qb_6_89=1.8
.ic q_7_89=0
.ic qb_7_89=1.8
.ic q_8_89=0
.ic qb_8_89=1.8
.ic q_9_89=0
.ic qb_9_89=1.8
.ic q_10_89=0
.ic qb_10_89=1.8
.ic q_11_89=0
.ic qb_11_89=1.8
.ic q_12_89=0
.ic qb_12_89=1.8
.ic q_13_89=0
.ic qb_13_89=1.8
.ic q_14_89=0
.ic qb_14_89=1.8
.ic q_15_89=0
.ic qb_15_89=1.8
.ic q_16_89=0
.ic qb_16_89=1.8
.ic q_17_89=0
.ic qb_17_89=1.8
.ic q_18_89=0
.ic qb_18_89=1.8
.ic q_19_89=0
.ic qb_19_89=1.8
.ic q_20_89=0
.ic qb_20_89=1.8
.ic q_21_89=0
.ic qb_21_89=1.8
.ic q_22_89=0
.ic qb_22_89=1.8
.ic q_23_89=0
.ic qb_23_89=1.8
.ic q_24_89=0
.ic qb_24_89=1.8
.ic q_25_89=0
.ic qb_25_89=1.8
.ic q_26_89=0
.ic qb_26_89=1.8
.ic q_27_89=0
.ic qb_27_89=1.8
.ic q_28_89=0
.ic qb_28_89=1.8
.ic q_29_89=0
.ic qb_29_89=1.8
.ic q_30_89=0
.ic qb_30_89=1.8
.ic q_31_89=0
.ic qb_31_89=1.8
.ic q_32_89=0
.ic qb_32_89=1.8
.ic q_33_89=0
.ic qb_33_89=1.8
.ic q_34_89=0
.ic qb_34_89=1.8
.ic q_35_89=0
.ic qb_35_89=1.8
.ic q_36_89=0
.ic qb_36_89=1.8
.ic q_37_89=0
.ic qb_37_89=1.8
.ic q_38_89=0
.ic qb_38_89=1.8
.ic q_39_89=0
.ic qb_39_89=1.8
.ic q_40_89=0
.ic qb_40_89=1.8
.ic q_41_89=0
.ic qb_41_89=1.8
.ic q_42_89=0
.ic qb_42_89=1.8
.ic q_43_89=0
.ic qb_43_89=1.8
.ic q_44_89=0
.ic qb_44_89=1.8
.ic q_45_89=0
.ic qb_45_89=1.8
.ic q_46_89=0
.ic qb_46_89=1.8
.ic q_47_89=0
.ic qb_47_89=1.8
.ic q_48_89=0
.ic qb_48_89=1.8
.ic q_49_89=0
.ic qb_49_89=1.8
.ic q_50_89=0
.ic qb_50_89=1.8
.ic q_51_89=0
.ic qb_51_89=1.8
.ic q_52_89=0
.ic qb_52_89=1.8
.ic q_53_89=0
.ic qb_53_89=1.8
.ic q_54_89=0
.ic qb_54_89=1.8
.ic q_55_89=0
.ic qb_55_89=1.8
.ic q_56_89=0
.ic qb_56_89=1.8
.ic q_57_89=0
.ic qb_57_89=1.8
.ic q_58_89=0
.ic qb_58_89=1.8
.ic q_59_89=0
.ic qb_59_89=1.8
.ic q_60_89=0
.ic qb_60_89=1.8
.ic q_61_89=0
.ic qb_61_89=1.8
.ic q_62_89=0
.ic qb_62_89=1.8
.ic q_63_89=0
.ic qb_63_89=1.8
.ic q_64_89=0
.ic qb_64_89=1.8
.ic q_65_89=0
.ic qb_65_89=1.8
.ic q_66_89=0
.ic qb_66_89=1.8
.ic q_67_89=0
.ic qb_67_89=1.8
.ic q_68_89=0
.ic qb_68_89=1.8
.ic q_69_89=0
.ic qb_69_89=1.8
.ic q_70_89=0
.ic qb_70_89=1.8
.ic q_71_89=0
.ic qb_71_89=1.8
.ic q_72_89=0
.ic qb_72_89=1.8
.ic q_73_89=0
.ic qb_73_89=1.8
.ic q_74_89=0
.ic qb_74_89=1.8
.ic q_75_89=0
.ic qb_75_89=1.8
.ic q_76_89=0
.ic qb_76_89=1.8
.ic q_77_89=0
.ic qb_77_89=1.8
.ic q_78_89=0
.ic qb_78_89=1.8
.ic q_79_89=0
.ic qb_79_89=1.8
.ic q_80_89=0
.ic qb_80_89=1.8
.ic q_81_89=0
.ic qb_81_89=1.8
.ic q_82_89=0
.ic qb_82_89=1.8
.ic q_83_89=0
.ic qb_83_89=1.8
.ic q_84_89=0
.ic qb_84_89=1.8
.ic q_85_89=0
.ic qb_85_89=1.8
.ic q_86_89=0
.ic qb_86_89=1.8
.ic q_87_89=0
.ic qb_87_89=1.8
.ic q_88_89=0
.ic qb_88_89=1.8
.ic q_89_89=0
.ic qb_89_89=1.8
.ic q_90_89=0
.ic qb_90_89=1.8
.ic q_91_89=0
.ic qb_91_89=1.8
.ic q_92_89=0
.ic qb_92_89=1.8
.ic q_93_89=0
.ic qb_93_89=1.8
.ic q_94_89=0
.ic qb_94_89=1.8
.ic q_95_89=0
.ic qb_95_89=1.8
.ic q_96_89=0
.ic qb_96_89=1.8
.ic q_97_89=0
.ic qb_97_89=1.8
.ic q_98_89=0
.ic qb_98_89=1.8
.ic q_99_89=0
.ic qb_99_89=1.8
.ic q_0_90=0
.ic qb_0_90=1.8
.ic q_1_90=0
.ic qb_1_90=1.8
.ic q_2_90=0
.ic qb_2_90=1.8
.ic q_3_90=0
.ic qb_3_90=1.8
.ic q_4_90=0
.ic qb_4_90=1.8
.ic q_5_90=0
.ic qb_5_90=1.8
.ic q_6_90=0
.ic qb_6_90=1.8
.ic q_7_90=0
.ic qb_7_90=1.8
.ic q_8_90=0
.ic qb_8_90=1.8
.ic q_9_90=0
.ic qb_9_90=1.8
.ic q_10_90=0
.ic qb_10_90=1.8
.ic q_11_90=0
.ic qb_11_90=1.8
.ic q_12_90=0
.ic qb_12_90=1.8
.ic q_13_90=0
.ic qb_13_90=1.8
.ic q_14_90=0
.ic qb_14_90=1.8
.ic q_15_90=0
.ic qb_15_90=1.8
.ic q_16_90=0
.ic qb_16_90=1.8
.ic q_17_90=0
.ic qb_17_90=1.8
.ic q_18_90=0
.ic qb_18_90=1.8
.ic q_19_90=0
.ic qb_19_90=1.8
.ic q_20_90=0
.ic qb_20_90=1.8
.ic q_21_90=0
.ic qb_21_90=1.8
.ic q_22_90=0
.ic qb_22_90=1.8
.ic q_23_90=0
.ic qb_23_90=1.8
.ic q_24_90=0
.ic qb_24_90=1.8
.ic q_25_90=0
.ic qb_25_90=1.8
.ic q_26_90=0
.ic qb_26_90=1.8
.ic q_27_90=0
.ic qb_27_90=1.8
.ic q_28_90=0
.ic qb_28_90=1.8
.ic q_29_90=0
.ic qb_29_90=1.8
.ic q_30_90=0
.ic qb_30_90=1.8
.ic q_31_90=0
.ic qb_31_90=1.8
.ic q_32_90=0
.ic qb_32_90=1.8
.ic q_33_90=0
.ic qb_33_90=1.8
.ic q_34_90=0
.ic qb_34_90=1.8
.ic q_35_90=0
.ic qb_35_90=1.8
.ic q_36_90=0
.ic qb_36_90=1.8
.ic q_37_90=0
.ic qb_37_90=1.8
.ic q_38_90=0
.ic qb_38_90=1.8
.ic q_39_90=0
.ic qb_39_90=1.8
.ic q_40_90=0
.ic qb_40_90=1.8
.ic q_41_90=0
.ic qb_41_90=1.8
.ic q_42_90=0
.ic qb_42_90=1.8
.ic q_43_90=0
.ic qb_43_90=1.8
.ic q_44_90=0
.ic qb_44_90=1.8
.ic q_45_90=0
.ic qb_45_90=1.8
.ic q_46_90=0
.ic qb_46_90=1.8
.ic q_47_90=0
.ic qb_47_90=1.8
.ic q_48_90=0
.ic qb_48_90=1.8
.ic q_49_90=0
.ic qb_49_90=1.8
.ic q_50_90=0
.ic qb_50_90=1.8
.ic q_51_90=0
.ic qb_51_90=1.8
.ic q_52_90=0
.ic qb_52_90=1.8
.ic q_53_90=0
.ic qb_53_90=1.8
.ic q_54_90=0
.ic qb_54_90=1.8
.ic q_55_90=0
.ic qb_55_90=1.8
.ic q_56_90=0
.ic qb_56_90=1.8
.ic q_57_90=0
.ic qb_57_90=1.8
.ic q_58_90=0
.ic qb_58_90=1.8
.ic q_59_90=0
.ic qb_59_90=1.8
.ic q_60_90=0
.ic qb_60_90=1.8
.ic q_61_90=0
.ic qb_61_90=1.8
.ic q_62_90=0
.ic qb_62_90=1.8
.ic q_63_90=0
.ic qb_63_90=1.8
.ic q_64_90=0
.ic qb_64_90=1.8
.ic q_65_90=0
.ic qb_65_90=1.8
.ic q_66_90=0
.ic qb_66_90=1.8
.ic q_67_90=0
.ic qb_67_90=1.8
.ic q_68_90=0
.ic qb_68_90=1.8
.ic q_69_90=0
.ic qb_69_90=1.8
.ic q_70_90=0
.ic qb_70_90=1.8
.ic q_71_90=0
.ic qb_71_90=1.8
.ic q_72_90=0
.ic qb_72_90=1.8
.ic q_73_90=0
.ic qb_73_90=1.8
.ic q_74_90=0
.ic qb_74_90=1.8
.ic q_75_90=0
.ic qb_75_90=1.8
.ic q_76_90=0
.ic qb_76_90=1.8
.ic q_77_90=0
.ic qb_77_90=1.8
.ic q_78_90=0
.ic qb_78_90=1.8
.ic q_79_90=0
.ic qb_79_90=1.8
.ic q_80_90=0
.ic qb_80_90=1.8
.ic q_81_90=0
.ic qb_81_90=1.8
.ic q_82_90=0
.ic qb_82_90=1.8
.ic q_83_90=0
.ic qb_83_90=1.8
.ic q_84_90=0
.ic qb_84_90=1.8
.ic q_85_90=0
.ic qb_85_90=1.8
.ic q_86_90=0
.ic qb_86_90=1.8
.ic q_87_90=0
.ic qb_87_90=1.8
.ic q_88_90=0
.ic qb_88_90=1.8
.ic q_89_90=0
.ic qb_89_90=1.8
.ic q_90_90=0
.ic qb_90_90=1.8
.ic q_91_90=0
.ic qb_91_90=1.8
.ic q_92_90=0
.ic qb_92_90=1.8
.ic q_93_90=0
.ic qb_93_90=1.8
.ic q_94_90=0
.ic qb_94_90=1.8
.ic q_95_90=0
.ic qb_95_90=1.8
.ic q_96_90=0
.ic qb_96_90=1.8
.ic q_97_90=0
.ic qb_97_90=1.8
.ic q_98_90=0
.ic qb_98_90=1.8
.ic q_99_90=0
.ic qb_99_90=1.8
.ic q_0_91=0
.ic qb_0_91=1.8
.ic q_1_91=0
.ic qb_1_91=1.8
.ic q_2_91=0
.ic qb_2_91=1.8
.ic q_3_91=0
.ic qb_3_91=1.8
.ic q_4_91=0
.ic qb_4_91=1.8
.ic q_5_91=0
.ic qb_5_91=1.8
.ic q_6_91=0
.ic qb_6_91=1.8
.ic q_7_91=0
.ic qb_7_91=1.8
.ic q_8_91=0
.ic qb_8_91=1.8
.ic q_9_91=0
.ic qb_9_91=1.8
.ic q_10_91=0
.ic qb_10_91=1.8
.ic q_11_91=0
.ic qb_11_91=1.8
.ic q_12_91=0
.ic qb_12_91=1.8
.ic q_13_91=0
.ic qb_13_91=1.8
.ic q_14_91=0
.ic qb_14_91=1.8
.ic q_15_91=0
.ic qb_15_91=1.8
.ic q_16_91=0
.ic qb_16_91=1.8
.ic q_17_91=0
.ic qb_17_91=1.8
.ic q_18_91=0
.ic qb_18_91=1.8
.ic q_19_91=0
.ic qb_19_91=1.8
.ic q_20_91=0
.ic qb_20_91=1.8
.ic q_21_91=0
.ic qb_21_91=1.8
.ic q_22_91=0
.ic qb_22_91=1.8
.ic q_23_91=0
.ic qb_23_91=1.8
.ic q_24_91=0
.ic qb_24_91=1.8
.ic q_25_91=0
.ic qb_25_91=1.8
.ic q_26_91=0
.ic qb_26_91=1.8
.ic q_27_91=0
.ic qb_27_91=1.8
.ic q_28_91=0
.ic qb_28_91=1.8
.ic q_29_91=0
.ic qb_29_91=1.8
.ic q_30_91=0
.ic qb_30_91=1.8
.ic q_31_91=0
.ic qb_31_91=1.8
.ic q_32_91=0
.ic qb_32_91=1.8
.ic q_33_91=0
.ic qb_33_91=1.8
.ic q_34_91=0
.ic qb_34_91=1.8
.ic q_35_91=0
.ic qb_35_91=1.8
.ic q_36_91=0
.ic qb_36_91=1.8
.ic q_37_91=0
.ic qb_37_91=1.8
.ic q_38_91=0
.ic qb_38_91=1.8
.ic q_39_91=0
.ic qb_39_91=1.8
.ic q_40_91=0
.ic qb_40_91=1.8
.ic q_41_91=0
.ic qb_41_91=1.8
.ic q_42_91=0
.ic qb_42_91=1.8
.ic q_43_91=0
.ic qb_43_91=1.8
.ic q_44_91=0
.ic qb_44_91=1.8
.ic q_45_91=0
.ic qb_45_91=1.8
.ic q_46_91=0
.ic qb_46_91=1.8
.ic q_47_91=0
.ic qb_47_91=1.8
.ic q_48_91=0
.ic qb_48_91=1.8
.ic q_49_91=0
.ic qb_49_91=1.8
.ic q_50_91=0
.ic qb_50_91=1.8
.ic q_51_91=0
.ic qb_51_91=1.8
.ic q_52_91=0
.ic qb_52_91=1.8
.ic q_53_91=0
.ic qb_53_91=1.8
.ic q_54_91=0
.ic qb_54_91=1.8
.ic q_55_91=0
.ic qb_55_91=1.8
.ic q_56_91=0
.ic qb_56_91=1.8
.ic q_57_91=0
.ic qb_57_91=1.8
.ic q_58_91=0
.ic qb_58_91=1.8
.ic q_59_91=0
.ic qb_59_91=1.8
.ic q_60_91=0
.ic qb_60_91=1.8
.ic q_61_91=0
.ic qb_61_91=1.8
.ic q_62_91=0
.ic qb_62_91=1.8
.ic q_63_91=0
.ic qb_63_91=1.8
.ic q_64_91=0
.ic qb_64_91=1.8
.ic q_65_91=0
.ic qb_65_91=1.8
.ic q_66_91=0
.ic qb_66_91=1.8
.ic q_67_91=0
.ic qb_67_91=1.8
.ic q_68_91=0
.ic qb_68_91=1.8
.ic q_69_91=0
.ic qb_69_91=1.8
.ic q_70_91=0
.ic qb_70_91=1.8
.ic q_71_91=0
.ic qb_71_91=1.8
.ic q_72_91=0
.ic qb_72_91=1.8
.ic q_73_91=0
.ic qb_73_91=1.8
.ic q_74_91=0
.ic qb_74_91=1.8
.ic q_75_91=0
.ic qb_75_91=1.8
.ic q_76_91=0
.ic qb_76_91=1.8
.ic q_77_91=0
.ic qb_77_91=1.8
.ic q_78_91=0
.ic qb_78_91=1.8
.ic q_79_91=0
.ic qb_79_91=1.8
.ic q_80_91=0
.ic qb_80_91=1.8
.ic q_81_91=0
.ic qb_81_91=1.8
.ic q_82_91=0
.ic qb_82_91=1.8
.ic q_83_91=0
.ic qb_83_91=1.8
.ic q_84_91=0
.ic qb_84_91=1.8
.ic q_85_91=0
.ic qb_85_91=1.8
.ic q_86_91=0
.ic qb_86_91=1.8
.ic q_87_91=0
.ic qb_87_91=1.8
.ic q_88_91=0
.ic qb_88_91=1.8
.ic q_89_91=0
.ic qb_89_91=1.8
.ic q_90_91=0
.ic qb_90_91=1.8
.ic q_91_91=0
.ic qb_91_91=1.8
.ic q_92_91=0
.ic qb_92_91=1.8
.ic q_93_91=0
.ic qb_93_91=1.8
.ic q_94_91=0
.ic qb_94_91=1.8
.ic q_95_91=0
.ic qb_95_91=1.8
.ic q_96_91=0
.ic qb_96_91=1.8
.ic q_97_91=0
.ic qb_97_91=1.8
.ic q_98_91=0
.ic qb_98_91=1.8
.ic q_99_91=0
.ic qb_99_91=1.8
.ic q_0_92=0
.ic qb_0_92=1.8
.ic q_1_92=0
.ic qb_1_92=1.8
.ic q_2_92=0
.ic qb_2_92=1.8
.ic q_3_92=0
.ic qb_3_92=1.8
.ic q_4_92=0
.ic qb_4_92=1.8
.ic q_5_92=0
.ic qb_5_92=1.8
.ic q_6_92=0
.ic qb_6_92=1.8
.ic q_7_92=0
.ic qb_7_92=1.8
.ic q_8_92=0
.ic qb_8_92=1.8
.ic q_9_92=0
.ic qb_9_92=1.8
.ic q_10_92=0
.ic qb_10_92=1.8
.ic q_11_92=0
.ic qb_11_92=1.8
.ic q_12_92=0
.ic qb_12_92=1.8
.ic q_13_92=0
.ic qb_13_92=1.8
.ic q_14_92=0
.ic qb_14_92=1.8
.ic q_15_92=0
.ic qb_15_92=1.8
.ic q_16_92=0
.ic qb_16_92=1.8
.ic q_17_92=0
.ic qb_17_92=1.8
.ic q_18_92=0
.ic qb_18_92=1.8
.ic q_19_92=0
.ic qb_19_92=1.8
.ic q_20_92=0
.ic qb_20_92=1.8
.ic q_21_92=0
.ic qb_21_92=1.8
.ic q_22_92=0
.ic qb_22_92=1.8
.ic q_23_92=0
.ic qb_23_92=1.8
.ic q_24_92=0
.ic qb_24_92=1.8
.ic q_25_92=0
.ic qb_25_92=1.8
.ic q_26_92=0
.ic qb_26_92=1.8
.ic q_27_92=0
.ic qb_27_92=1.8
.ic q_28_92=0
.ic qb_28_92=1.8
.ic q_29_92=0
.ic qb_29_92=1.8
.ic q_30_92=0
.ic qb_30_92=1.8
.ic q_31_92=0
.ic qb_31_92=1.8
.ic q_32_92=0
.ic qb_32_92=1.8
.ic q_33_92=0
.ic qb_33_92=1.8
.ic q_34_92=0
.ic qb_34_92=1.8
.ic q_35_92=0
.ic qb_35_92=1.8
.ic q_36_92=0
.ic qb_36_92=1.8
.ic q_37_92=0
.ic qb_37_92=1.8
.ic q_38_92=0
.ic qb_38_92=1.8
.ic q_39_92=0
.ic qb_39_92=1.8
.ic q_40_92=0
.ic qb_40_92=1.8
.ic q_41_92=0
.ic qb_41_92=1.8
.ic q_42_92=0
.ic qb_42_92=1.8
.ic q_43_92=0
.ic qb_43_92=1.8
.ic q_44_92=0
.ic qb_44_92=1.8
.ic q_45_92=0
.ic qb_45_92=1.8
.ic q_46_92=0
.ic qb_46_92=1.8
.ic q_47_92=0
.ic qb_47_92=1.8
.ic q_48_92=0
.ic qb_48_92=1.8
.ic q_49_92=0
.ic qb_49_92=1.8
.ic q_50_92=0
.ic qb_50_92=1.8
.ic q_51_92=0
.ic qb_51_92=1.8
.ic q_52_92=0
.ic qb_52_92=1.8
.ic q_53_92=0
.ic qb_53_92=1.8
.ic q_54_92=0
.ic qb_54_92=1.8
.ic q_55_92=0
.ic qb_55_92=1.8
.ic q_56_92=0
.ic qb_56_92=1.8
.ic q_57_92=0
.ic qb_57_92=1.8
.ic q_58_92=0
.ic qb_58_92=1.8
.ic q_59_92=0
.ic qb_59_92=1.8
.ic q_60_92=0
.ic qb_60_92=1.8
.ic q_61_92=0
.ic qb_61_92=1.8
.ic q_62_92=0
.ic qb_62_92=1.8
.ic q_63_92=0
.ic qb_63_92=1.8
.ic q_64_92=0
.ic qb_64_92=1.8
.ic q_65_92=0
.ic qb_65_92=1.8
.ic q_66_92=0
.ic qb_66_92=1.8
.ic q_67_92=0
.ic qb_67_92=1.8
.ic q_68_92=0
.ic qb_68_92=1.8
.ic q_69_92=0
.ic qb_69_92=1.8
.ic q_70_92=0
.ic qb_70_92=1.8
.ic q_71_92=0
.ic qb_71_92=1.8
.ic q_72_92=0
.ic qb_72_92=1.8
.ic q_73_92=0
.ic qb_73_92=1.8
.ic q_74_92=0
.ic qb_74_92=1.8
.ic q_75_92=0
.ic qb_75_92=1.8
.ic q_76_92=0
.ic qb_76_92=1.8
.ic q_77_92=0
.ic qb_77_92=1.8
.ic q_78_92=0
.ic qb_78_92=1.8
.ic q_79_92=0
.ic qb_79_92=1.8
.ic q_80_92=0
.ic qb_80_92=1.8
.ic q_81_92=0
.ic qb_81_92=1.8
.ic q_82_92=0
.ic qb_82_92=1.8
.ic q_83_92=0
.ic qb_83_92=1.8
.ic q_84_92=0
.ic qb_84_92=1.8
.ic q_85_92=0
.ic qb_85_92=1.8
.ic q_86_92=0
.ic qb_86_92=1.8
.ic q_87_92=0
.ic qb_87_92=1.8
.ic q_88_92=0
.ic qb_88_92=1.8
.ic q_89_92=0
.ic qb_89_92=1.8
.ic q_90_92=0
.ic qb_90_92=1.8
.ic q_91_92=0
.ic qb_91_92=1.8
.ic q_92_92=0
.ic qb_92_92=1.8
.ic q_93_92=0
.ic qb_93_92=1.8
.ic q_94_92=0
.ic qb_94_92=1.8
.ic q_95_92=0
.ic qb_95_92=1.8
.ic q_96_92=0
.ic qb_96_92=1.8
.ic q_97_92=0
.ic qb_97_92=1.8
.ic q_98_92=0
.ic qb_98_92=1.8
.ic q_99_92=0
.ic qb_99_92=1.8
.ic q_0_93=0
.ic qb_0_93=1.8
.ic q_1_93=0
.ic qb_1_93=1.8
.ic q_2_93=0
.ic qb_2_93=1.8
.ic q_3_93=0
.ic qb_3_93=1.8
.ic q_4_93=0
.ic qb_4_93=1.8
.ic q_5_93=0
.ic qb_5_93=1.8
.ic q_6_93=0
.ic qb_6_93=1.8
.ic q_7_93=0
.ic qb_7_93=1.8
.ic q_8_93=0
.ic qb_8_93=1.8
.ic q_9_93=0
.ic qb_9_93=1.8
.ic q_10_93=0
.ic qb_10_93=1.8
.ic q_11_93=0
.ic qb_11_93=1.8
.ic q_12_93=0
.ic qb_12_93=1.8
.ic q_13_93=0
.ic qb_13_93=1.8
.ic q_14_93=0
.ic qb_14_93=1.8
.ic q_15_93=0
.ic qb_15_93=1.8
.ic q_16_93=0
.ic qb_16_93=1.8
.ic q_17_93=0
.ic qb_17_93=1.8
.ic q_18_93=0
.ic qb_18_93=1.8
.ic q_19_93=0
.ic qb_19_93=1.8
.ic q_20_93=0
.ic qb_20_93=1.8
.ic q_21_93=0
.ic qb_21_93=1.8
.ic q_22_93=0
.ic qb_22_93=1.8
.ic q_23_93=0
.ic qb_23_93=1.8
.ic q_24_93=0
.ic qb_24_93=1.8
.ic q_25_93=0
.ic qb_25_93=1.8
.ic q_26_93=0
.ic qb_26_93=1.8
.ic q_27_93=0
.ic qb_27_93=1.8
.ic q_28_93=0
.ic qb_28_93=1.8
.ic q_29_93=0
.ic qb_29_93=1.8
.ic q_30_93=0
.ic qb_30_93=1.8
.ic q_31_93=0
.ic qb_31_93=1.8
.ic q_32_93=0
.ic qb_32_93=1.8
.ic q_33_93=0
.ic qb_33_93=1.8
.ic q_34_93=0
.ic qb_34_93=1.8
.ic q_35_93=0
.ic qb_35_93=1.8
.ic q_36_93=0
.ic qb_36_93=1.8
.ic q_37_93=0
.ic qb_37_93=1.8
.ic q_38_93=0
.ic qb_38_93=1.8
.ic q_39_93=0
.ic qb_39_93=1.8
.ic q_40_93=0
.ic qb_40_93=1.8
.ic q_41_93=0
.ic qb_41_93=1.8
.ic q_42_93=0
.ic qb_42_93=1.8
.ic q_43_93=0
.ic qb_43_93=1.8
.ic q_44_93=0
.ic qb_44_93=1.8
.ic q_45_93=0
.ic qb_45_93=1.8
.ic q_46_93=0
.ic qb_46_93=1.8
.ic q_47_93=0
.ic qb_47_93=1.8
.ic q_48_93=0
.ic qb_48_93=1.8
.ic q_49_93=0
.ic qb_49_93=1.8
.ic q_50_93=0
.ic qb_50_93=1.8
.ic q_51_93=0
.ic qb_51_93=1.8
.ic q_52_93=0
.ic qb_52_93=1.8
.ic q_53_93=0
.ic qb_53_93=1.8
.ic q_54_93=0
.ic qb_54_93=1.8
.ic q_55_93=0
.ic qb_55_93=1.8
.ic q_56_93=0
.ic qb_56_93=1.8
.ic q_57_93=0
.ic qb_57_93=1.8
.ic q_58_93=0
.ic qb_58_93=1.8
.ic q_59_93=0
.ic qb_59_93=1.8
.ic q_60_93=0
.ic qb_60_93=1.8
.ic q_61_93=0
.ic qb_61_93=1.8
.ic q_62_93=0
.ic qb_62_93=1.8
.ic q_63_93=0
.ic qb_63_93=1.8
.ic q_64_93=0
.ic qb_64_93=1.8
.ic q_65_93=0
.ic qb_65_93=1.8
.ic q_66_93=0
.ic qb_66_93=1.8
.ic q_67_93=0
.ic qb_67_93=1.8
.ic q_68_93=0
.ic qb_68_93=1.8
.ic q_69_93=0
.ic qb_69_93=1.8
.ic q_70_93=0
.ic qb_70_93=1.8
.ic q_71_93=0
.ic qb_71_93=1.8
.ic q_72_93=0
.ic qb_72_93=1.8
.ic q_73_93=0
.ic qb_73_93=1.8
.ic q_74_93=0
.ic qb_74_93=1.8
.ic q_75_93=0
.ic qb_75_93=1.8
.ic q_76_93=0
.ic qb_76_93=1.8
.ic q_77_93=0
.ic qb_77_93=1.8
.ic q_78_93=0
.ic qb_78_93=1.8
.ic q_79_93=0
.ic qb_79_93=1.8
.ic q_80_93=0
.ic qb_80_93=1.8
.ic q_81_93=0
.ic qb_81_93=1.8
.ic q_82_93=0
.ic qb_82_93=1.8
.ic q_83_93=0
.ic qb_83_93=1.8
.ic q_84_93=0
.ic qb_84_93=1.8
.ic q_85_93=0
.ic qb_85_93=1.8
.ic q_86_93=0
.ic qb_86_93=1.8
.ic q_87_93=0
.ic qb_87_93=1.8
.ic q_88_93=0
.ic qb_88_93=1.8
.ic q_89_93=0
.ic qb_89_93=1.8
.ic q_90_93=0
.ic qb_90_93=1.8
.ic q_91_93=0
.ic qb_91_93=1.8
.ic q_92_93=0
.ic qb_92_93=1.8
.ic q_93_93=0
.ic qb_93_93=1.8
.ic q_94_93=0
.ic qb_94_93=1.8
.ic q_95_93=0
.ic qb_95_93=1.8
.ic q_96_93=0
.ic qb_96_93=1.8
.ic q_97_93=0
.ic qb_97_93=1.8
.ic q_98_93=0
.ic qb_98_93=1.8
.ic q_99_93=0
.ic qb_99_93=1.8
.ic q_0_94=0
.ic qb_0_94=1.8
.ic q_1_94=0
.ic qb_1_94=1.8
.ic q_2_94=0
.ic qb_2_94=1.8
.ic q_3_94=0
.ic qb_3_94=1.8
.ic q_4_94=0
.ic qb_4_94=1.8
.ic q_5_94=0
.ic qb_5_94=1.8
.ic q_6_94=0
.ic qb_6_94=1.8
.ic q_7_94=0
.ic qb_7_94=1.8
.ic q_8_94=0
.ic qb_8_94=1.8
.ic q_9_94=0
.ic qb_9_94=1.8
.ic q_10_94=0
.ic qb_10_94=1.8
.ic q_11_94=0
.ic qb_11_94=1.8
.ic q_12_94=0
.ic qb_12_94=1.8
.ic q_13_94=0
.ic qb_13_94=1.8
.ic q_14_94=0
.ic qb_14_94=1.8
.ic q_15_94=0
.ic qb_15_94=1.8
.ic q_16_94=0
.ic qb_16_94=1.8
.ic q_17_94=0
.ic qb_17_94=1.8
.ic q_18_94=0
.ic qb_18_94=1.8
.ic q_19_94=0
.ic qb_19_94=1.8
.ic q_20_94=0
.ic qb_20_94=1.8
.ic q_21_94=0
.ic qb_21_94=1.8
.ic q_22_94=0
.ic qb_22_94=1.8
.ic q_23_94=0
.ic qb_23_94=1.8
.ic q_24_94=0
.ic qb_24_94=1.8
.ic q_25_94=0
.ic qb_25_94=1.8
.ic q_26_94=0
.ic qb_26_94=1.8
.ic q_27_94=0
.ic qb_27_94=1.8
.ic q_28_94=0
.ic qb_28_94=1.8
.ic q_29_94=0
.ic qb_29_94=1.8
.ic q_30_94=0
.ic qb_30_94=1.8
.ic q_31_94=0
.ic qb_31_94=1.8
.ic q_32_94=0
.ic qb_32_94=1.8
.ic q_33_94=0
.ic qb_33_94=1.8
.ic q_34_94=0
.ic qb_34_94=1.8
.ic q_35_94=0
.ic qb_35_94=1.8
.ic q_36_94=0
.ic qb_36_94=1.8
.ic q_37_94=0
.ic qb_37_94=1.8
.ic q_38_94=0
.ic qb_38_94=1.8
.ic q_39_94=0
.ic qb_39_94=1.8
.ic q_40_94=0
.ic qb_40_94=1.8
.ic q_41_94=0
.ic qb_41_94=1.8
.ic q_42_94=0
.ic qb_42_94=1.8
.ic q_43_94=0
.ic qb_43_94=1.8
.ic q_44_94=0
.ic qb_44_94=1.8
.ic q_45_94=0
.ic qb_45_94=1.8
.ic q_46_94=0
.ic qb_46_94=1.8
.ic q_47_94=0
.ic qb_47_94=1.8
.ic q_48_94=0
.ic qb_48_94=1.8
.ic q_49_94=0
.ic qb_49_94=1.8
.ic q_50_94=0
.ic qb_50_94=1.8
.ic q_51_94=0
.ic qb_51_94=1.8
.ic q_52_94=0
.ic qb_52_94=1.8
.ic q_53_94=0
.ic qb_53_94=1.8
.ic q_54_94=0
.ic qb_54_94=1.8
.ic q_55_94=0
.ic qb_55_94=1.8
.ic q_56_94=0
.ic qb_56_94=1.8
.ic q_57_94=0
.ic qb_57_94=1.8
.ic q_58_94=0
.ic qb_58_94=1.8
.ic q_59_94=0
.ic qb_59_94=1.8
.ic q_60_94=0
.ic qb_60_94=1.8
.ic q_61_94=0
.ic qb_61_94=1.8
.ic q_62_94=0
.ic qb_62_94=1.8
.ic q_63_94=0
.ic qb_63_94=1.8
.ic q_64_94=0
.ic qb_64_94=1.8
.ic q_65_94=0
.ic qb_65_94=1.8
.ic q_66_94=0
.ic qb_66_94=1.8
.ic q_67_94=0
.ic qb_67_94=1.8
.ic q_68_94=0
.ic qb_68_94=1.8
.ic q_69_94=0
.ic qb_69_94=1.8
.ic q_70_94=0
.ic qb_70_94=1.8
.ic q_71_94=0
.ic qb_71_94=1.8
.ic q_72_94=0
.ic qb_72_94=1.8
.ic q_73_94=0
.ic qb_73_94=1.8
.ic q_74_94=0
.ic qb_74_94=1.8
.ic q_75_94=0
.ic qb_75_94=1.8
.ic q_76_94=0
.ic qb_76_94=1.8
.ic q_77_94=0
.ic qb_77_94=1.8
.ic q_78_94=0
.ic qb_78_94=1.8
.ic q_79_94=0
.ic qb_79_94=1.8
.ic q_80_94=0
.ic qb_80_94=1.8
.ic q_81_94=0
.ic qb_81_94=1.8
.ic q_82_94=0
.ic qb_82_94=1.8
.ic q_83_94=0
.ic qb_83_94=1.8
.ic q_84_94=0
.ic qb_84_94=1.8
.ic q_85_94=0
.ic qb_85_94=1.8
.ic q_86_94=0
.ic qb_86_94=1.8
.ic q_87_94=0
.ic qb_87_94=1.8
.ic q_88_94=0
.ic qb_88_94=1.8
.ic q_89_94=0
.ic qb_89_94=1.8
.ic q_90_94=0
.ic qb_90_94=1.8
.ic q_91_94=0
.ic qb_91_94=1.8
.ic q_92_94=0
.ic qb_92_94=1.8
.ic q_93_94=0
.ic qb_93_94=1.8
.ic q_94_94=0
.ic qb_94_94=1.8
.ic q_95_94=0
.ic qb_95_94=1.8
.ic q_96_94=0
.ic qb_96_94=1.8
.ic q_97_94=0
.ic qb_97_94=1.8
.ic q_98_94=0
.ic qb_98_94=1.8
.ic q_99_94=0
.ic qb_99_94=1.8
.ic q_0_95=0
.ic qb_0_95=1.8
.ic q_1_95=0
.ic qb_1_95=1.8
.ic q_2_95=0
.ic qb_2_95=1.8
.ic q_3_95=0
.ic qb_3_95=1.8
.ic q_4_95=0
.ic qb_4_95=1.8
.ic q_5_95=0
.ic qb_5_95=1.8
.ic q_6_95=0
.ic qb_6_95=1.8
.ic q_7_95=0
.ic qb_7_95=1.8
.ic q_8_95=0
.ic qb_8_95=1.8
.ic q_9_95=0
.ic qb_9_95=1.8
.ic q_10_95=0
.ic qb_10_95=1.8
.ic q_11_95=0
.ic qb_11_95=1.8
.ic q_12_95=0
.ic qb_12_95=1.8
.ic q_13_95=0
.ic qb_13_95=1.8
.ic q_14_95=0
.ic qb_14_95=1.8
.ic q_15_95=0
.ic qb_15_95=1.8
.ic q_16_95=0
.ic qb_16_95=1.8
.ic q_17_95=0
.ic qb_17_95=1.8
.ic q_18_95=0
.ic qb_18_95=1.8
.ic q_19_95=0
.ic qb_19_95=1.8
.ic q_20_95=0
.ic qb_20_95=1.8
.ic q_21_95=0
.ic qb_21_95=1.8
.ic q_22_95=0
.ic qb_22_95=1.8
.ic q_23_95=0
.ic qb_23_95=1.8
.ic q_24_95=0
.ic qb_24_95=1.8
.ic q_25_95=0
.ic qb_25_95=1.8
.ic q_26_95=0
.ic qb_26_95=1.8
.ic q_27_95=0
.ic qb_27_95=1.8
.ic q_28_95=0
.ic qb_28_95=1.8
.ic q_29_95=0
.ic qb_29_95=1.8
.ic q_30_95=0
.ic qb_30_95=1.8
.ic q_31_95=0
.ic qb_31_95=1.8
.ic q_32_95=0
.ic qb_32_95=1.8
.ic q_33_95=0
.ic qb_33_95=1.8
.ic q_34_95=0
.ic qb_34_95=1.8
.ic q_35_95=0
.ic qb_35_95=1.8
.ic q_36_95=0
.ic qb_36_95=1.8
.ic q_37_95=0
.ic qb_37_95=1.8
.ic q_38_95=0
.ic qb_38_95=1.8
.ic q_39_95=0
.ic qb_39_95=1.8
.ic q_40_95=0
.ic qb_40_95=1.8
.ic q_41_95=0
.ic qb_41_95=1.8
.ic q_42_95=0
.ic qb_42_95=1.8
.ic q_43_95=0
.ic qb_43_95=1.8
.ic q_44_95=0
.ic qb_44_95=1.8
.ic q_45_95=0
.ic qb_45_95=1.8
.ic q_46_95=0
.ic qb_46_95=1.8
.ic q_47_95=0
.ic qb_47_95=1.8
.ic q_48_95=0
.ic qb_48_95=1.8
.ic q_49_95=0
.ic qb_49_95=1.8
.ic q_50_95=0
.ic qb_50_95=1.8
.ic q_51_95=0
.ic qb_51_95=1.8
.ic q_52_95=0
.ic qb_52_95=1.8
.ic q_53_95=0
.ic qb_53_95=1.8
.ic q_54_95=0
.ic qb_54_95=1.8
.ic q_55_95=0
.ic qb_55_95=1.8
.ic q_56_95=0
.ic qb_56_95=1.8
.ic q_57_95=0
.ic qb_57_95=1.8
.ic q_58_95=0
.ic qb_58_95=1.8
.ic q_59_95=0
.ic qb_59_95=1.8
.ic q_60_95=0
.ic qb_60_95=1.8
.ic q_61_95=0
.ic qb_61_95=1.8
.ic q_62_95=0
.ic qb_62_95=1.8
.ic q_63_95=0
.ic qb_63_95=1.8
.ic q_64_95=0
.ic qb_64_95=1.8
.ic q_65_95=0
.ic qb_65_95=1.8
.ic q_66_95=0
.ic qb_66_95=1.8
.ic q_67_95=0
.ic qb_67_95=1.8
.ic q_68_95=0
.ic qb_68_95=1.8
.ic q_69_95=0
.ic qb_69_95=1.8
.ic q_70_95=0
.ic qb_70_95=1.8
.ic q_71_95=0
.ic qb_71_95=1.8
.ic q_72_95=0
.ic qb_72_95=1.8
.ic q_73_95=0
.ic qb_73_95=1.8
.ic q_74_95=0
.ic qb_74_95=1.8
.ic q_75_95=0
.ic qb_75_95=1.8
.ic q_76_95=0
.ic qb_76_95=1.8
.ic q_77_95=0
.ic qb_77_95=1.8
.ic q_78_95=0
.ic qb_78_95=1.8
.ic q_79_95=0
.ic qb_79_95=1.8
.ic q_80_95=0
.ic qb_80_95=1.8
.ic q_81_95=0
.ic qb_81_95=1.8
.ic q_82_95=0
.ic qb_82_95=1.8
.ic q_83_95=0
.ic qb_83_95=1.8
.ic q_84_95=0
.ic qb_84_95=1.8
.ic q_85_95=0
.ic qb_85_95=1.8
.ic q_86_95=0
.ic qb_86_95=1.8
.ic q_87_95=0
.ic qb_87_95=1.8
.ic q_88_95=0
.ic qb_88_95=1.8
.ic q_89_95=0
.ic qb_89_95=1.8
.ic q_90_95=0
.ic qb_90_95=1.8
.ic q_91_95=0
.ic qb_91_95=1.8
.ic q_92_95=0
.ic qb_92_95=1.8
.ic q_93_95=0
.ic qb_93_95=1.8
.ic q_94_95=0
.ic qb_94_95=1.8
.ic q_95_95=0
.ic qb_95_95=1.8
.ic q_96_95=0
.ic qb_96_95=1.8
.ic q_97_95=0
.ic qb_97_95=1.8
.ic q_98_95=0
.ic qb_98_95=1.8
.ic q_99_95=0
.ic qb_99_95=1.8
.ic q_0_96=0
.ic qb_0_96=1.8
.ic q_1_96=0
.ic qb_1_96=1.8
.ic q_2_96=0
.ic qb_2_96=1.8
.ic q_3_96=0
.ic qb_3_96=1.8
.ic q_4_96=0
.ic qb_4_96=1.8
.ic q_5_96=0
.ic qb_5_96=1.8
.ic q_6_96=0
.ic qb_6_96=1.8
.ic q_7_96=0
.ic qb_7_96=1.8
.ic q_8_96=0
.ic qb_8_96=1.8
.ic q_9_96=0
.ic qb_9_96=1.8
.ic q_10_96=0
.ic qb_10_96=1.8
.ic q_11_96=0
.ic qb_11_96=1.8
.ic q_12_96=0
.ic qb_12_96=1.8
.ic q_13_96=0
.ic qb_13_96=1.8
.ic q_14_96=0
.ic qb_14_96=1.8
.ic q_15_96=0
.ic qb_15_96=1.8
.ic q_16_96=0
.ic qb_16_96=1.8
.ic q_17_96=0
.ic qb_17_96=1.8
.ic q_18_96=0
.ic qb_18_96=1.8
.ic q_19_96=0
.ic qb_19_96=1.8
.ic q_20_96=0
.ic qb_20_96=1.8
.ic q_21_96=0
.ic qb_21_96=1.8
.ic q_22_96=0
.ic qb_22_96=1.8
.ic q_23_96=0
.ic qb_23_96=1.8
.ic q_24_96=0
.ic qb_24_96=1.8
.ic q_25_96=0
.ic qb_25_96=1.8
.ic q_26_96=0
.ic qb_26_96=1.8
.ic q_27_96=0
.ic qb_27_96=1.8
.ic q_28_96=0
.ic qb_28_96=1.8
.ic q_29_96=0
.ic qb_29_96=1.8
.ic q_30_96=0
.ic qb_30_96=1.8
.ic q_31_96=0
.ic qb_31_96=1.8
.ic q_32_96=0
.ic qb_32_96=1.8
.ic q_33_96=0
.ic qb_33_96=1.8
.ic q_34_96=0
.ic qb_34_96=1.8
.ic q_35_96=0
.ic qb_35_96=1.8
.ic q_36_96=0
.ic qb_36_96=1.8
.ic q_37_96=0
.ic qb_37_96=1.8
.ic q_38_96=0
.ic qb_38_96=1.8
.ic q_39_96=0
.ic qb_39_96=1.8
.ic q_40_96=0
.ic qb_40_96=1.8
.ic q_41_96=0
.ic qb_41_96=1.8
.ic q_42_96=0
.ic qb_42_96=1.8
.ic q_43_96=0
.ic qb_43_96=1.8
.ic q_44_96=0
.ic qb_44_96=1.8
.ic q_45_96=0
.ic qb_45_96=1.8
.ic q_46_96=0
.ic qb_46_96=1.8
.ic q_47_96=0
.ic qb_47_96=1.8
.ic q_48_96=0
.ic qb_48_96=1.8
.ic q_49_96=0
.ic qb_49_96=1.8
.ic q_50_96=0
.ic qb_50_96=1.8
.ic q_51_96=0
.ic qb_51_96=1.8
.ic q_52_96=0
.ic qb_52_96=1.8
.ic q_53_96=0
.ic qb_53_96=1.8
.ic q_54_96=0
.ic qb_54_96=1.8
.ic q_55_96=0
.ic qb_55_96=1.8
.ic q_56_96=0
.ic qb_56_96=1.8
.ic q_57_96=0
.ic qb_57_96=1.8
.ic q_58_96=0
.ic qb_58_96=1.8
.ic q_59_96=0
.ic qb_59_96=1.8
.ic q_60_96=0
.ic qb_60_96=1.8
.ic q_61_96=0
.ic qb_61_96=1.8
.ic q_62_96=0
.ic qb_62_96=1.8
.ic q_63_96=0
.ic qb_63_96=1.8
.ic q_64_96=0
.ic qb_64_96=1.8
.ic q_65_96=0
.ic qb_65_96=1.8
.ic q_66_96=0
.ic qb_66_96=1.8
.ic q_67_96=0
.ic qb_67_96=1.8
.ic q_68_96=0
.ic qb_68_96=1.8
.ic q_69_96=0
.ic qb_69_96=1.8
.ic q_70_96=0
.ic qb_70_96=1.8
.ic q_71_96=0
.ic qb_71_96=1.8
.ic q_72_96=0
.ic qb_72_96=1.8
.ic q_73_96=0
.ic qb_73_96=1.8
.ic q_74_96=0
.ic qb_74_96=1.8
.ic q_75_96=0
.ic qb_75_96=1.8
.ic q_76_96=0
.ic qb_76_96=1.8
.ic q_77_96=0
.ic qb_77_96=1.8
.ic q_78_96=0
.ic qb_78_96=1.8
.ic q_79_96=0
.ic qb_79_96=1.8
.ic q_80_96=0
.ic qb_80_96=1.8
.ic q_81_96=0
.ic qb_81_96=1.8
.ic q_82_96=0
.ic qb_82_96=1.8
.ic q_83_96=0
.ic qb_83_96=1.8
.ic q_84_96=0
.ic qb_84_96=1.8
.ic q_85_96=0
.ic qb_85_96=1.8
.ic q_86_96=0
.ic qb_86_96=1.8
.ic q_87_96=0
.ic qb_87_96=1.8
.ic q_88_96=0
.ic qb_88_96=1.8
.ic q_89_96=0
.ic qb_89_96=1.8
.ic q_90_96=0
.ic qb_90_96=1.8
.ic q_91_96=0
.ic qb_91_96=1.8
.ic q_92_96=0
.ic qb_92_96=1.8
.ic q_93_96=0
.ic qb_93_96=1.8
.ic q_94_96=0
.ic qb_94_96=1.8
.ic q_95_96=0
.ic qb_95_96=1.8
.ic q_96_96=0
.ic qb_96_96=1.8
.ic q_97_96=0
.ic qb_97_96=1.8
.ic q_98_96=0
.ic qb_98_96=1.8
.ic q_99_96=0
.ic qb_99_96=1.8
.ic q_0_97=0
.ic qb_0_97=1.8
.ic q_1_97=0
.ic qb_1_97=1.8
.ic q_2_97=0
.ic qb_2_97=1.8
.ic q_3_97=0
.ic qb_3_97=1.8
.ic q_4_97=0
.ic qb_4_97=1.8
.ic q_5_97=0
.ic qb_5_97=1.8
.ic q_6_97=0
.ic qb_6_97=1.8
.ic q_7_97=0
.ic qb_7_97=1.8
.ic q_8_97=0
.ic qb_8_97=1.8
.ic q_9_97=0
.ic qb_9_97=1.8
.ic q_10_97=0
.ic qb_10_97=1.8
.ic q_11_97=0
.ic qb_11_97=1.8
.ic q_12_97=0
.ic qb_12_97=1.8
.ic q_13_97=0
.ic qb_13_97=1.8
.ic q_14_97=0
.ic qb_14_97=1.8
.ic q_15_97=0
.ic qb_15_97=1.8
.ic q_16_97=0
.ic qb_16_97=1.8
.ic q_17_97=0
.ic qb_17_97=1.8
.ic q_18_97=0
.ic qb_18_97=1.8
.ic q_19_97=0
.ic qb_19_97=1.8
.ic q_20_97=0
.ic qb_20_97=1.8
.ic q_21_97=0
.ic qb_21_97=1.8
.ic q_22_97=0
.ic qb_22_97=1.8
.ic q_23_97=0
.ic qb_23_97=1.8
.ic q_24_97=0
.ic qb_24_97=1.8
.ic q_25_97=0
.ic qb_25_97=1.8
.ic q_26_97=0
.ic qb_26_97=1.8
.ic q_27_97=0
.ic qb_27_97=1.8
.ic q_28_97=0
.ic qb_28_97=1.8
.ic q_29_97=0
.ic qb_29_97=1.8
.ic q_30_97=0
.ic qb_30_97=1.8
.ic q_31_97=0
.ic qb_31_97=1.8
.ic q_32_97=0
.ic qb_32_97=1.8
.ic q_33_97=0
.ic qb_33_97=1.8
.ic q_34_97=0
.ic qb_34_97=1.8
.ic q_35_97=0
.ic qb_35_97=1.8
.ic q_36_97=0
.ic qb_36_97=1.8
.ic q_37_97=0
.ic qb_37_97=1.8
.ic q_38_97=0
.ic qb_38_97=1.8
.ic q_39_97=0
.ic qb_39_97=1.8
.ic q_40_97=0
.ic qb_40_97=1.8
.ic q_41_97=0
.ic qb_41_97=1.8
.ic q_42_97=0
.ic qb_42_97=1.8
.ic q_43_97=0
.ic qb_43_97=1.8
.ic q_44_97=0
.ic qb_44_97=1.8
.ic q_45_97=0
.ic qb_45_97=1.8
.ic q_46_97=0
.ic qb_46_97=1.8
.ic q_47_97=0
.ic qb_47_97=1.8
.ic q_48_97=0
.ic qb_48_97=1.8
.ic q_49_97=0
.ic qb_49_97=1.8
.ic q_50_97=0
.ic qb_50_97=1.8
.ic q_51_97=0
.ic qb_51_97=1.8
.ic q_52_97=0
.ic qb_52_97=1.8
.ic q_53_97=0
.ic qb_53_97=1.8
.ic q_54_97=0
.ic qb_54_97=1.8
.ic q_55_97=0
.ic qb_55_97=1.8
.ic q_56_97=0
.ic qb_56_97=1.8
.ic q_57_97=0
.ic qb_57_97=1.8
.ic q_58_97=0
.ic qb_58_97=1.8
.ic q_59_97=0
.ic qb_59_97=1.8
.ic q_60_97=0
.ic qb_60_97=1.8
.ic q_61_97=0
.ic qb_61_97=1.8
.ic q_62_97=0
.ic qb_62_97=1.8
.ic q_63_97=0
.ic qb_63_97=1.8
.ic q_64_97=0
.ic qb_64_97=1.8
.ic q_65_97=0
.ic qb_65_97=1.8
.ic q_66_97=0
.ic qb_66_97=1.8
.ic q_67_97=0
.ic qb_67_97=1.8
.ic q_68_97=0
.ic qb_68_97=1.8
.ic q_69_97=0
.ic qb_69_97=1.8
.ic q_70_97=0
.ic qb_70_97=1.8
.ic q_71_97=0
.ic qb_71_97=1.8
.ic q_72_97=0
.ic qb_72_97=1.8
.ic q_73_97=0
.ic qb_73_97=1.8
.ic q_74_97=0
.ic qb_74_97=1.8
.ic q_75_97=0
.ic qb_75_97=1.8
.ic q_76_97=0
.ic qb_76_97=1.8
.ic q_77_97=0
.ic qb_77_97=1.8
.ic q_78_97=0
.ic qb_78_97=1.8
.ic q_79_97=0
.ic qb_79_97=1.8
.ic q_80_97=0
.ic qb_80_97=1.8
.ic q_81_97=0
.ic qb_81_97=1.8
.ic q_82_97=0
.ic qb_82_97=1.8
.ic q_83_97=0
.ic qb_83_97=1.8
.ic q_84_97=0
.ic qb_84_97=1.8
.ic q_85_97=0
.ic qb_85_97=1.8
.ic q_86_97=0
.ic qb_86_97=1.8
.ic q_87_97=0
.ic qb_87_97=1.8
.ic q_88_97=0
.ic qb_88_97=1.8
.ic q_89_97=0
.ic qb_89_97=1.8
.ic q_90_97=0
.ic qb_90_97=1.8
.ic q_91_97=0
.ic qb_91_97=1.8
.ic q_92_97=0
.ic qb_92_97=1.8
.ic q_93_97=0
.ic qb_93_97=1.8
.ic q_94_97=0
.ic qb_94_97=1.8
.ic q_95_97=0
.ic qb_95_97=1.8
.ic q_96_97=0
.ic qb_96_97=1.8
.ic q_97_97=0
.ic qb_97_97=1.8
.ic q_98_97=0
.ic qb_98_97=1.8
.ic q_99_97=0
.ic qb_99_97=1.8
.ic q_0_98=0
.ic qb_0_98=1.8
.ic q_1_98=0
.ic qb_1_98=1.8
.ic q_2_98=0
.ic qb_2_98=1.8
.ic q_3_98=0
.ic qb_3_98=1.8
.ic q_4_98=0
.ic qb_4_98=1.8
.ic q_5_98=0
.ic qb_5_98=1.8
.ic q_6_98=0
.ic qb_6_98=1.8
.ic q_7_98=0
.ic qb_7_98=1.8
.ic q_8_98=0
.ic qb_8_98=1.8
.ic q_9_98=0
.ic qb_9_98=1.8
.ic q_10_98=0
.ic qb_10_98=1.8
.ic q_11_98=0
.ic qb_11_98=1.8
.ic q_12_98=0
.ic qb_12_98=1.8
.ic q_13_98=0
.ic qb_13_98=1.8
.ic q_14_98=0
.ic qb_14_98=1.8
.ic q_15_98=0
.ic qb_15_98=1.8
.ic q_16_98=0
.ic qb_16_98=1.8
.ic q_17_98=0
.ic qb_17_98=1.8
.ic q_18_98=0
.ic qb_18_98=1.8
.ic q_19_98=0
.ic qb_19_98=1.8
.ic q_20_98=0
.ic qb_20_98=1.8
.ic q_21_98=0
.ic qb_21_98=1.8
.ic q_22_98=0
.ic qb_22_98=1.8
.ic q_23_98=0
.ic qb_23_98=1.8
.ic q_24_98=0
.ic qb_24_98=1.8
.ic q_25_98=0
.ic qb_25_98=1.8
.ic q_26_98=0
.ic qb_26_98=1.8
.ic q_27_98=0
.ic qb_27_98=1.8
.ic q_28_98=0
.ic qb_28_98=1.8
.ic q_29_98=0
.ic qb_29_98=1.8
.ic q_30_98=0
.ic qb_30_98=1.8
.ic q_31_98=0
.ic qb_31_98=1.8
.ic q_32_98=0
.ic qb_32_98=1.8
.ic q_33_98=0
.ic qb_33_98=1.8
.ic q_34_98=0
.ic qb_34_98=1.8
.ic q_35_98=0
.ic qb_35_98=1.8
.ic q_36_98=0
.ic qb_36_98=1.8
.ic q_37_98=0
.ic qb_37_98=1.8
.ic q_38_98=0
.ic qb_38_98=1.8
.ic q_39_98=0
.ic qb_39_98=1.8
.ic q_40_98=0
.ic qb_40_98=1.8
.ic q_41_98=0
.ic qb_41_98=1.8
.ic q_42_98=0
.ic qb_42_98=1.8
.ic q_43_98=0
.ic qb_43_98=1.8
.ic q_44_98=0
.ic qb_44_98=1.8
.ic q_45_98=0
.ic qb_45_98=1.8
.ic q_46_98=0
.ic qb_46_98=1.8
.ic q_47_98=0
.ic qb_47_98=1.8
.ic q_48_98=0
.ic qb_48_98=1.8
.ic q_49_98=0
.ic qb_49_98=1.8
.ic q_50_98=0
.ic qb_50_98=1.8
.ic q_51_98=0
.ic qb_51_98=1.8
.ic q_52_98=0
.ic qb_52_98=1.8
.ic q_53_98=0
.ic qb_53_98=1.8
.ic q_54_98=0
.ic qb_54_98=1.8
.ic q_55_98=0
.ic qb_55_98=1.8
.ic q_56_98=0
.ic qb_56_98=1.8
.ic q_57_98=0
.ic qb_57_98=1.8
.ic q_58_98=0
.ic qb_58_98=1.8
.ic q_59_98=0
.ic qb_59_98=1.8
.ic q_60_98=0
.ic qb_60_98=1.8
.ic q_61_98=0
.ic qb_61_98=1.8
.ic q_62_98=0
.ic qb_62_98=1.8
.ic q_63_98=0
.ic qb_63_98=1.8
.ic q_64_98=0
.ic qb_64_98=1.8
.ic q_65_98=0
.ic qb_65_98=1.8
.ic q_66_98=0
.ic qb_66_98=1.8
.ic q_67_98=0
.ic qb_67_98=1.8
.ic q_68_98=0
.ic qb_68_98=1.8
.ic q_69_98=0
.ic qb_69_98=1.8
.ic q_70_98=0
.ic qb_70_98=1.8
.ic q_71_98=0
.ic qb_71_98=1.8
.ic q_72_98=0
.ic qb_72_98=1.8
.ic q_73_98=0
.ic qb_73_98=1.8
.ic q_74_98=0
.ic qb_74_98=1.8
.ic q_75_98=0
.ic qb_75_98=1.8
.ic q_76_98=0
.ic qb_76_98=1.8
.ic q_77_98=0
.ic qb_77_98=1.8
.ic q_78_98=0
.ic qb_78_98=1.8
.ic q_79_98=0
.ic qb_79_98=1.8
.ic q_80_98=0
.ic qb_80_98=1.8
.ic q_81_98=0
.ic qb_81_98=1.8
.ic q_82_98=0
.ic qb_82_98=1.8
.ic q_83_98=0
.ic qb_83_98=1.8
.ic q_84_98=0
.ic qb_84_98=1.8
.ic q_85_98=0
.ic qb_85_98=1.8
.ic q_86_98=0
.ic qb_86_98=1.8
.ic q_87_98=0
.ic qb_87_98=1.8
.ic q_88_98=0
.ic qb_88_98=1.8
.ic q_89_98=0
.ic qb_89_98=1.8
.ic q_90_98=0
.ic qb_90_98=1.8
.ic q_91_98=0
.ic qb_91_98=1.8
.ic q_92_98=0
.ic qb_92_98=1.8
.ic q_93_98=0
.ic qb_93_98=1.8
.ic q_94_98=0
.ic qb_94_98=1.8
.ic q_95_98=0
.ic qb_95_98=1.8
.ic q_96_98=0
.ic qb_96_98=1.8
.ic q_97_98=0
.ic qb_97_98=1.8
.ic q_98_98=0
.ic qb_98_98=1.8
.ic q_99_98=0
.ic qb_99_98=1.8
.ic q_0_99=0
.ic qb_0_99=1.8
.ic q_1_99=0
.ic qb_1_99=1.8
.ic q_2_99=0
.ic qb_2_99=1.8
.ic q_3_99=0
.ic qb_3_99=1.8
.ic q_4_99=0
.ic qb_4_99=1.8
.ic q_5_99=0
.ic qb_5_99=1.8
.ic q_6_99=0
.ic qb_6_99=1.8
.ic q_7_99=0
.ic qb_7_99=1.8
.ic q_8_99=0
.ic qb_8_99=1.8
.ic q_9_99=0
.ic qb_9_99=1.8
.ic q_10_99=0
.ic qb_10_99=1.8
.ic q_11_99=0
.ic qb_11_99=1.8
.ic q_12_99=0
.ic qb_12_99=1.8
.ic q_13_99=0
.ic qb_13_99=1.8
.ic q_14_99=0
.ic qb_14_99=1.8
.ic q_15_99=0
.ic qb_15_99=1.8
.ic q_16_99=0
.ic qb_16_99=1.8
.ic q_17_99=0
.ic qb_17_99=1.8
.ic q_18_99=0
.ic qb_18_99=1.8
.ic q_19_99=0
.ic qb_19_99=1.8
.ic q_20_99=0
.ic qb_20_99=1.8
.ic q_21_99=0
.ic qb_21_99=1.8
.ic q_22_99=0
.ic qb_22_99=1.8
.ic q_23_99=0
.ic qb_23_99=1.8
.ic q_24_99=0
.ic qb_24_99=1.8
.ic q_25_99=0
.ic qb_25_99=1.8
.ic q_26_99=0
.ic qb_26_99=1.8
.ic q_27_99=0
.ic qb_27_99=1.8
.ic q_28_99=0
.ic qb_28_99=1.8
.ic q_29_99=0
.ic qb_29_99=1.8
.ic q_30_99=0
.ic qb_30_99=1.8
.ic q_31_99=0
.ic qb_31_99=1.8
.ic q_32_99=0
.ic qb_32_99=1.8
.ic q_33_99=0
.ic qb_33_99=1.8
.ic q_34_99=0
.ic qb_34_99=1.8
.ic q_35_99=0
.ic qb_35_99=1.8
.ic q_36_99=0
.ic qb_36_99=1.8
.ic q_37_99=0
.ic qb_37_99=1.8
.ic q_38_99=0
.ic qb_38_99=1.8
.ic q_39_99=0
.ic qb_39_99=1.8
.ic q_40_99=0
.ic qb_40_99=1.8
.ic q_41_99=0
.ic qb_41_99=1.8
.ic q_42_99=0
.ic qb_42_99=1.8
.ic q_43_99=0
.ic qb_43_99=1.8
.ic q_44_99=0
.ic qb_44_99=1.8
.ic q_45_99=0
.ic qb_45_99=1.8
.ic q_46_99=0
.ic qb_46_99=1.8
.ic q_47_99=0
.ic qb_47_99=1.8
.ic q_48_99=0
.ic qb_48_99=1.8
.ic q_49_99=0
.ic qb_49_99=1.8
.ic q_50_99=0
.ic qb_50_99=1.8
.ic q_51_99=0
.ic qb_51_99=1.8
.ic q_52_99=0
.ic qb_52_99=1.8
.ic q_53_99=0
.ic qb_53_99=1.8
.ic q_54_99=0
.ic qb_54_99=1.8
.ic q_55_99=0
.ic qb_55_99=1.8
.ic q_56_99=0
.ic qb_56_99=1.8
.ic q_57_99=0
.ic qb_57_99=1.8
.ic q_58_99=0
.ic qb_58_99=1.8
.ic q_59_99=0
.ic qb_59_99=1.8
.ic q_60_99=0
.ic qb_60_99=1.8
.ic q_61_99=0
.ic qb_61_99=1.8
.ic q_62_99=0
.ic qb_62_99=1.8
.ic q_63_99=0
.ic qb_63_99=1.8
.ic q_64_99=0
.ic qb_64_99=1.8
.ic q_65_99=0
.ic qb_65_99=1.8
.ic q_66_99=0
.ic qb_66_99=1.8
.ic q_67_99=0
.ic qb_67_99=1.8
.ic q_68_99=0
.ic qb_68_99=1.8
.ic q_69_99=0
.ic qb_69_99=1.8
.ic q_70_99=0
.ic qb_70_99=1.8
.ic q_71_99=0
.ic qb_71_99=1.8
.ic q_72_99=0
.ic qb_72_99=1.8
.ic q_73_99=0
.ic qb_73_99=1.8
.ic q_74_99=0
.ic qb_74_99=1.8
.ic q_75_99=0
.ic qb_75_99=1.8
.ic q_76_99=0
.ic qb_76_99=1.8
.ic q_77_99=0
.ic qb_77_99=1.8
.ic q_78_99=0
.ic qb_78_99=1.8
.ic q_79_99=0
.ic qb_79_99=1.8
.ic q_80_99=0
.ic qb_80_99=1.8
.ic q_81_99=0
.ic qb_81_99=1.8
.ic q_82_99=0
.ic qb_82_99=1.8
.ic q_83_99=0
.ic qb_83_99=1.8
.ic q_84_99=0
.ic qb_84_99=1.8
.ic q_85_99=0
.ic qb_85_99=1.8
.ic q_86_99=0
.ic qb_86_99=1.8
.ic q_87_99=0
.ic qb_87_99=1.8
.ic q_88_99=0
.ic qb_88_99=1.8
.ic q_89_99=0
.ic qb_89_99=1.8
.ic q_90_99=0
.ic qb_90_99=1.8
.ic q_91_99=0
.ic qb_91_99=1.8
.ic q_92_99=0
.ic qb_92_99=1.8
.ic q_93_99=0
.ic qb_93_99=1.8
.ic q_94_99=0
.ic qb_94_99=1.8
.ic q_95_99=0
.ic qb_95_99=1.8
.ic q_96_99=0
.ic qb_96_99=1.8
.ic q_97_99=0
.ic qb_97_99=1.8
.ic q_98_99=0
.ic qb_98_99=1.8
.ic q_99_99=1.8
.ic qb_99_99=0
.param W1=4
.param W5=2
X0_0 q_0_0 qb_0_0 bit_0_0 bitb_0_0 word0_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_0 q_1_0 qb_1_0 bit_1_0 bitb_1_0 word1_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_0 q_2_0 qb_2_0 bit_2_0 bitb_2_0 word2_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_0 q_3_0 qb_3_0 bit_3_0 bitb_3_0 word3_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_0 q_4_0 qb_4_0 bit_4_0 bitb_4_0 word4_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_0 q_5_0 qb_5_0 bit_5_0 bitb_5_0 word5_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_0 q_6_0 qb_6_0 bit_6_0 bitb_6_0 word6_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_0 q_7_0 qb_7_0 bit_7_0 bitb_7_0 word7_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_0 q_8_0 qb_8_0 bit_8_0 bitb_8_0 word8_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_0 q_9_0 qb_9_0 bit_9_0 bitb_9_0 word9_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_0 q_10_0 qb_10_0 bit_10_0 bitb_10_0 word10_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_0 q_11_0 qb_11_0 bit_11_0 bitb_11_0 word11_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_0 q_12_0 qb_12_0 bit_12_0 bitb_12_0 word12_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_0 q_13_0 qb_13_0 bit_13_0 bitb_13_0 word13_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_0 q_14_0 qb_14_0 bit_14_0 bitb_14_0 word14_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_0 q_15_0 qb_15_0 bit_15_0 bitb_15_0 word15_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_0 q_16_0 qb_16_0 bit_16_0 bitb_16_0 word16_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_0 q_17_0 qb_17_0 bit_17_0 bitb_17_0 word17_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_0 q_18_0 qb_18_0 bit_18_0 bitb_18_0 word18_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_0 q_19_0 qb_19_0 bit_19_0 bitb_19_0 word19_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_0 q_20_0 qb_20_0 bit_20_0 bitb_20_0 word20_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_0 q_21_0 qb_21_0 bit_21_0 bitb_21_0 word21_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_0 q_22_0 qb_22_0 bit_22_0 bitb_22_0 word22_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_0 q_23_0 qb_23_0 bit_23_0 bitb_23_0 word23_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_0 q_24_0 qb_24_0 bit_24_0 bitb_24_0 word24_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_0 q_25_0 qb_25_0 bit_25_0 bitb_25_0 word25_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_0 q_26_0 qb_26_0 bit_26_0 bitb_26_0 word26_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_0 q_27_0 qb_27_0 bit_27_0 bitb_27_0 word27_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_0 q_28_0 qb_28_0 bit_28_0 bitb_28_0 word28_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_0 q_29_0 qb_29_0 bit_29_0 bitb_29_0 word29_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_0 q_30_0 qb_30_0 bit_30_0 bitb_30_0 word30_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_0 q_31_0 qb_31_0 bit_31_0 bitb_31_0 word31_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_0 q_32_0 qb_32_0 bit_32_0 bitb_32_0 word32_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_0 q_33_0 qb_33_0 bit_33_0 bitb_33_0 word33_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_0 q_34_0 qb_34_0 bit_34_0 bitb_34_0 word34_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_0 q_35_0 qb_35_0 bit_35_0 bitb_35_0 word35_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_0 q_36_0 qb_36_0 bit_36_0 bitb_36_0 word36_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_0 q_37_0 qb_37_0 bit_37_0 bitb_37_0 word37_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_0 q_38_0 qb_38_0 bit_38_0 bitb_38_0 word38_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_0 q_39_0 qb_39_0 bit_39_0 bitb_39_0 word39_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_0 q_40_0 qb_40_0 bit_40_0 bitb_40_0 word40_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_0 q_41_0 qb_41_0 bit_41_0 bitb_41_0 word41_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_0 q_42_0 qb_42_0 bit_42_0 bitb_42_0 word42_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_0 q_43_0 qb_43_0 bit_43_0 bitb_43_0 word43_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_0 q_44_0 qb_44_0 bit_44_0 bitb_44_0 word44_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_0 q_45_0 qb_45_0 bit_45_0 bitb_45_0 word45_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_0 q_46_0 qb_46_0 bit_46_0 bitb_46_0 word46_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_0 q_47_0 qb_47_0 bit_47_0 bitb_47_0 word47_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_0 q_48_0 qb_48_0 bit_48_0 bitb_48_0 word48_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_0 q_49_0 qb_49_0 bit_49_0 bitb_49_0 word49_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_0 q_50_0 qb_50_0 bit_50_0 bitb_50_0 word50_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_0 q_51_0 qb_51_0 bit_51_0 bitb_51_0 word51_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_0 q_52_0 qb_52_0 bit_52_0 bitb_52_0 word52_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_0 q_53_0 qb_53_0 bit_53_0 bitb_53_0 word53_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_0 q_54_0 qb_54_0 bit_54_0 bitb_54_0 word54_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_0 q_55_0 qb_55_0 bit_55_0 bitb_55_0 word55_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_0 q_56_0 qb_56_0 bit_56_0 bitb_56_0 word56_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_0 q_57_0 qb_57_0 bit_57_0 bitb_57_0 word57_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_0 q_58_0 qb_58_0 bit_58_0 bitb_58_0 word58_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_0 q_59_0 qb_59_0 bit_59_0 bitb_59_0 word59_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_0 q_60_0 qb_60_0 bit_60_0 bitb_60_0 word60_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_0 q_61_0 qb_61_0 bit_61_0 bitb_61_0 word61_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_0 q_62_0 qb_62_0 bit_62_0 bitb_62_0 word62_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_0 q_63_0 qb_63_0 bit_63_0 bitb_63_0 word63_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_0 q_64_0 qb_64_0 bit_64_0 bitb_64_0 word64_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_0 q_65_0 qb_65_0 bit_65_0 bitb_65_0 word65_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_0 q_66_0 qb_66_0 bit_66_0 bitb_66_0 word66_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_0 q_67_0 qb_67_0 bit_67_0 bitb_67_0 word67_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_0 q_68_0 qb_68_0 bit_68_0 bitb_68_0 word68_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_0 q_69_0 qb_69_0 bit_69_0 bitb_69_0 word69_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_0 q_70_0 qb_70_0 bit_70_0 bitb_70_0 word70_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_0 q_71_0 qb_71_0 bit_71_0 bitb_71_0 word71_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_0 q_72_0 qb_72_0 bit_72_0 bitb_72_0 word72_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_0 q_73_0 qb_73_0 bit_73_0 bitb_73_0 word73_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_0 q_74_0 qb_74_0 bit_74_0 bitb_74_0 word74_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_0 q_75_0 qb_75_0 bit_75_0 bitb_75_0 word75_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_0 q_76_0 qb_76_0 bit_76_0 bitb_76_0 word76_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_0 q_77_0 qb_77_0 bit_77_0 bitb_77_0 word77_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_0 q_78_0 qb_78_0 bit_78_0 bitb_78_0 word78_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_0 q_79_0 qb_79_0 bit_79_0 bitb_79_0 word79_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_0 q_80_0 qb_80_0 bit_80_0 bitb_80_0 word80_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_0 q_81_0 qb_81_0 bit_81_0 bitb_81_0 word81_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_0 q_82_0 qb_82_0 bit_82_0 bitb_82_0 word82_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_0 q_83_0 qb_83_0 bit_83_0 bitb_83_0 word83_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_0 q_84_0 qb_84_0 bit_84_0 bitb_84_0 word84_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_0 q_85_0 qb_85_0 bit_85_0 bitb_85_0 word85_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_0 q_86_0 qb_86_0 bit_86_0 bitb_86_0 word86_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_0 q_87_0 qb_87_0 bit_87_0 bitb_87_0 word87_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_0 q_88_0 qb_88_0 bit_88_0 bitb_88_0 word88_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_0 q_89_0 qb_89_0 bit_89_0 bitb_89_0 word89_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_0 q_90_0 qb_90_0 bit_90_0 bitb_90_0 word90_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_0 q_91_0 qb_91_0 bit_91_0 bitb_91_0 word91_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_0 q_92_0 qb_92_0 bit_92_0 bitb_92_0 word92_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_0 q_93_0 qb_93_0 bit_93_0 bitb_93_0 word93_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_0 q_94_0 qb_94_0 bit_94_0 bitb_94_0 word94_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_0 q_95_0 qb_95_0 bit_95_0 bitb_95_0 word95_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_0 q_96_0 qb_96_0 bit_96_0 bitb_96_0 word96_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_0 q_97_0 qb_97_0 bit_97_0 bitb_97_0 word97_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_0 q_98_0 qb_98_0 bit_98_0 bitb_98_0 word98_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_0 q_99_0 qb_99_0 bit_99_0 bitb_99_0 word99_0 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_1 q_0_1 qb_0_1 bit_0_1 bitb_0_1 word0_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_1 q_1_1 qb_1_1 bit_1_1 bitb_1_1 word1_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_1 q_2_1 qb_2_1 bit_2_1 bitb_2_1 word2_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_1 q_3_1 qb_3_1 bit_3_1 bitb_3_1 word3_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_1 q_4_1 qb_4_1 bit_4_1 bitb_4_1 word4_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_1 q_5_1 qb_5_1 bit_5_1 bitb_5_1 word5_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_1 q_6_1 qb_6_1 bit_6_1 bitb_6_1 word6_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_1 q_7_1 qb_7_1 bit_7_1 bitb_7_1 word7_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_1 q_8_1 qb_8_1 bit_8_1 bitb_8_1 word8_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_1 q_9_1 qb_9_1 bit_9_1 bitb_9_1 word9_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_1 q_10_1 qb_10_1 bit_10_1 bitb_10_1 word10_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_1 q_11_1 qb_11_1 bit_11_1 bitb_11_1 word11_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_1 q_12_1 qb_12_1 bit_12_1 bitb_12_1 word12_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_1 q_13_1 qb_13_1 bit_13_1 bitb_13_1 word13_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_1 q_14_1 qb_14_1 bit_14_1 bitb_14_1 word14_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_1 q_15_1 qb_15_1 bit_15_1 bitb_15_1 word15_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_1 q_16_1 qb_16_1 bit_16_1 bitb_16_1 word16_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_1 q_17_1 qb_17_1 bit_17_1 bitb_17_1 word17_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_1 q_18_1 qb_18_1 bit_18_1 bitb_18_1 word18_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_1 q_19_1 qb_19_1 bit_19_1 bitb_19_1 word19_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_1 q_20_1 qb_20_1 bit_20_1 bitb_20_1 word20_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_1 q_21_1 qb_21_1 bit_21_1 bitb_21_1 word21_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_1 q_22_1 qb_22_1 bit_22_1 bitb_22_1 word22_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_1 q_23_1 qb_23_1 bit_23_1 bitb_23_1 word23_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_1 q_24_1 qb_24_1 bit_24_1 bitb_24_1 word24_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_1 q_25_1 qb_25_1 bit_25_1 bitb_25_1 word25_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_1 q_26_1 qb_26_1 bit_26_1 bitb_26_1 word26_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_1 q_27_1 qb_27_1 bit_27_1 bitb_27_1 word27_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_1 q_28_1 qb_28_1 bit_28_1 bitb_28_1 word28_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_1 q_29_1 qb_29_1 bit_29_1 bitb_29_1 word29_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_1 q_30_1 qb_30_1 bit_30_1 bitb_30_1 word30_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_1 q_31_1 qb_31_1 bit_31_1 bitb_31_1 word31_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_1 q_32_1 qb_32_1 bit_32_1 bitb_32_1 word32_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_1 q_33_1 qb_33_1 bit_33_1 bitb_33_1 word33_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_1 q_34_1 qb_34_1 bit_34_1 bitb_34_1 word34_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_1 q_35_1 qb_35_1 bit_35_1 bitb_35_1 word35_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_1 q_36_1 qb_36_1 bit_36_1 bitb_36_1 word36_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_1 q_37_1 qb_37_1 bit_37_1 bitb_37_1 word37_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_1 q_38_1 qb_38_1 bit_38_1 bitb_38_1 word38_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_1 q_39_1 qb_39_1 bit_39_1 bitb_39_1 word39_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_1 q_40_1 qb_40_1 bit_40_1 bitb_40_1 word40_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_1 q_41_1 qb_41_1 bit_41_1 bitb_41_1 word41_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_1 q_42_1 qb_42_1 bit_42_1 bitb_42_1 word42_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_1 q_43_1 qb_43_1 bit_43_1 bitb_43_1 word43_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_1 q_44_1 qb_44_1 bit_44_1 bitb_44_1 word44_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_1 q_45_1 qb_45_1 bit_45_1 bitb_45_1 word45_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_1 q_46_1 qb_46_1 bit_46_1 bitb_46_1 word46_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_1 q_47_1 qb_47_1 bit_47_1 bitb_47_1 word47_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_1 q_48_1 qb_48_1 bit_48_1 bitb_48_1 word48_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_1 q_49_1 qb_49_1 bit_49_1 bitb_49_1 word49_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_1 q_50_1 qb_50_1 bit_50_1 bitb_50_1 word50_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_1 q_51_1 qb_51_1 bit_51_1 bitb_51_1 word51_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_1 q_52_1 qb_52_1 bit_52_1 bitb_52_1 word52_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_1 q_53_1 qb_53_1 bit_53_1 bitb_53_1 word53_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_1 q_54_1 qb_54_1 bit_54_1 bitb_54_1 word54_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_1 q_55_1 qb_55_1 bit_55_1 bitb_55_1 word55_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_1 q_56_1 qb_56_1 bit_56_1 bitb_56_1 word56_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_1 q_57_1 qb_57_1 bit_57_1 bitb_57_1 word57_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_1 q_58_1 qb_58_1 bit_58_1 bitb_58_1 word58_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_1 q_59_1 qb_59_1 bit_59_1 bitb_59_1 word59_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_1 q_60_1 qb_60_1 bit_60_1 bitb_60_1 word60_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_1 q_61_1 qb_61_1 bit_61_1 bitb_61_1 word61_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_1 q_62_1 qb_62_1 bit_62_1 bitb_62_1 word62_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_1 q_63_1 qb_63_1 bit_63_1 bitb_63_1 word63_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_1 q_64_1 qb_64_1 bit_64_1 bitb_64_1 word64_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_1 q_65_1 qb_65_1 bit_65_1 bitb_65_1 word65_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_1 q_66_1 qb_66_1 bit_66_1 bitb_66_1 word66_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_1 q_67_1 qb_67_1 bit_67_1 bitb_67_1 word67_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_1 q_68_1 qb_68_1 bit_68_1 bitb_68_1 word68_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_1 q_69_1 qb_69_1 bit_69_1 bitb_69_1 word69_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_1 q_70_1 qb_70_1 bit_70_1 bitb_70_1 word70_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_1 q_71_1 qb_71_1 bit_71_1 bitb_71_1 word71_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_1 q_72_1 qb_72_1 bit_72_1 bitb_72_1 word72_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_1 q_73_1 qb_73_1 bit_73_1 bitb_73_1 word73_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_1 q_74_1 qb_74_1 bit_74_1 bitb_74_1 word74_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_1 q_75_1 qb_75_1 bit_75_1 bitb_75_1 word75_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_1 q_76_1 qb_76_1 bit_76_1 bitb_76_1 word76_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_1 q_77_1 qb_77_1 bit_77_1 bitb_77_1 word77_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_1 q_78_1 qb_78_1 bit_78_1 bitb_78_1 word78_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_1 q_79_1 qb_79_1 bit_79_1 bitb_79_1 word79_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_1 q_80_1 qb_80_1 bit_80_1 bitb_80_1 word80_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_1 q_81_1 qb_81_1 bit_81_1 bitb_81_1 word81_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_1 q_82_1 qb_82_1 bit_82_1 bitb_82_1 word82_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_1 q_83_1 qb_83_1 bit_83_1 bitb_83_1 word83_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_1 q_84_1 qb_84_1 bit_84_1 bitb_84_1 word84_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_1 q_85_1 qb_85_1 bit_85_1 bitb_85_1 word85_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_1 q_86_1 qb_86_1 bit_86_1 bitb_86_1 word86_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_1 q_87_1 qb_87_1 bit_87_1 bitb_87_1 word87_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_1 q_88_1 qb_88_1 bit_88_1 bitb_88_1 word88_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_1 q_89_1 qb_89_1 bit_89_1 bitb_89_1 word89_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_1 q_90_1 qb_90_1 bit_90_1 bitb_90_1 word90_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_1 q_91_1 qb_91_1 bit_91_1 bitb_91_1 word91_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_1 q_92_1 qb_92_1 bit_92_1 bitb_92_1 word92_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_1 q_93_1 qb_93_1 bit_93_1 bitb_93_1 word93_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_1 q_94_1 qb_94_1 bit_94_1 bitb_94_1 word94_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_1 q_95_1 qb_95_1 bit_95_1 bitb_95_1 word95_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_1 q_96_1 qb_96_1 bit_96_1 bitb_96_1 word96_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_1 q_97_1 qb_97_1 bit_97_1 bitb_97_1 word97_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_1 q_98_1 qb_98_1 bit_98_1 bitb_98_1 word98_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_1 q_99_1 qb_99_1 bit_99_1 bitb_99_1 word99_1 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_2 q_0_2 qb_0_2 bit_0_2 bitb_0_2 word0_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_2 q_1_2 qb_1_2 bit_1_2 bitb_1_2 word1_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_2 q_2_2 qb_2_2 bit_2_2 bitb_2_2 word2_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_2 q_3_2 qb_3_2 bit_3_2 bitb_3_2 word3_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_2 q_4_2 qb_4_2 bit_4_2 bitb_4_2 word4_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_2 q_5_2 qb_5_2 bit_5_2 bitb_5_2 word5_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_2 q_6_2 qb_6_2 bit_6_2 bitb_6_2 word6_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_2 q_7_2 qb_7_2 bit_7_2 bitb_7_2 word7_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_2 q_8_2 qb_8_2 bit_8_2 bitb_8_2 word8_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_2 q_9_2 qb_9_2 bit_9_2 bitb_9_2 word9_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_2 q_10_2 qb_10_2 bit_10_2 bitb_10_2 word10_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_2 q_11_2 qb_11_2 bit_11_2 bitb_11_2 word11_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_2 q_12_2 qb_12_2 bit_12_2 bitb_12_2 word12_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_2 q_13_2 qb_13_2 bit_13_2 bitb_13_2 word13_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_2 q_14_2 qb_14_2 bit_14_2 bitb_14_2 word14_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_2 q_15_2 qb_15_2 bit_15_2 bitb_15_2 word15_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_2 q_16_2 qb_16_2 bit_16_2 bitb_16_2 word16_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_2 q_17_2 qb_17_2 bit_17_2 bitb_17_2 word17_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_2 q_18_2 qb_18_2 bit_18_2 bitb_18_2 word18_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_2 q_19_2 qb_19_2 bit_19_2 bitb_19_2 word19_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_2 q_20_2 qb_20_2 bit_20_2 bitb_20_2 word20_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_2 q_21_2 qb_21_2 bit_21_2 bitb_21_2 word21_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_2 q_22_2 qb_22_2 bit_22_2 bitb_22_2 word22_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_2 q_23_2 qb_23_2 bit_23_2 bitb_23_2 word23_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_2 q_24_2 qb_24_2 bit_24_2 bitb_24_2 word24_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_2 q_25_2 qb_25_2 bit_25_2 bitb_25_2 word25_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_2 q_26_2 qb_26_2 bit_26_2 bitb_26_2 word26_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_2 q_27_2 qb_27_2 bit_27_2 bitb_27_2 word27_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_2 q_28_2 qb_28_2 bit_28_2 bitb_28_2 word28_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_2 q_29_2 qb_29_2 bit_29_2 bitb_29_2 word29_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_2 q_30_2 qb_30_2 bit_30_2 bitb_30_2 word30_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_2 q_31_2 qb_31_2 bit_31_2 bitb_31_2 word31_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_2 q_32_2 qb_32_2 bit_32_2 bitb_32_2 word32_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_2 q_33_2 qb_33_2 bit_33_2 bitb_33_2 word33_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_2 q_34_2 qb_34_2 bit_34_2 bitb_34_2 word34_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_2 q_35_2 qb_35_2 bit_35_2 bitb_35_2 word35_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_2 q_36_2 qb_36_2 bit_36_2 bitb_36_2 word36_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_2 q_37_2 qb_37_2 bit_37_2 bitb_37_2 word37_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_2 q_38_2 qb_38_2 bit_38_2 bitb_38_2 word38_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_2 q_39_2 qb_39_2 bit_39_2 bitb_39_2 word39_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_2 q_40_2 qb_40_2 bit_40_2 bitb_40_2 word40_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_2 q_41_2 qb_41_2 bit_41_2 bitb_41_2 word41_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_2 q_42_2 qb_42_2 bit_42_2 bitb_42_2 word42_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_2 q_43_2 qb_43_2 bit_43_2 bitb_43_2 word43_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_2 q_44_2 qb_44_2 bit_44_2 bitb_44_2 word44_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_2 q_45_2 qb_45_2 bit_45_2 bitb_45_2 word45_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_2 q_46_2 qb_46_2 bit_46_2 bitb_46_2 word46_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_2 q_47_2 qb_47_2 bit_47_2 bitb_47_2 word47_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_2 q_48_2 qb_48_2 bit_48_2 bitb_48_2 word48_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_2 q_49_2 qb_49_2 bit_49_2 bitb_49_2 word49_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_2 q_50_2 qb_50_2 bit_50_2 bitb_50_2 word50_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_2 q_51_2 qb_51_2 bit_51_2 bitb_51_2 word51_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_2 q_52_2 qb_52_2 bit_52_2 bitb_52_2 word52_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_2 q_53_2 qb_53_2 bit_53_2 bitb_53_2 word53_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_2 q_54_2 qb_54_2 bit_54_2 bitb_54_2 word54_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_2 q_55_2 qb_55_2 bit_55_2 bitb_55_2 word55_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_2 q_56_2 qb_56_2 bit_56_2 bitb_56_2 word56_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_2 q_57_2 qb_57_2 bit_57_2 bitb_57_2 word57_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_2 q_58_2 qb_58_2 bit_58_2 bitb_58_2 word58_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_2 q_59_2 qb_59_2 bit_59_2 bitb_59_2 word59_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_2 q_60_2 qb_60_2 bit_60_2 bitb_60_2 word60_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_2 q_61_2 qb_61_2 bit_61_2 bitb_61_2 word61_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_2 q_62_2 qb_62_2 bit_62_2 bitb_62_2 word62_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_2 q_63_2 qb_63_2 bit_63_2 bitb_63_2 word63_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_2 q_64_2 qb_64_2 bit_64_2 bitb_64_2 word64_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_2 q_65_2 qb_65_2 bit_65_2 bitb_65_2 word65_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_2 q_66_2 qb_66_2 bit_66_2 bitb_66_2 word66_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_2 q_67_2 qb_67_2 bit_67_2 bitb_67_2 word67_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_2 q_68_2 qb_68_2 bit_68_2 bitb_68_2 word68_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_2 q_69_2 qb_69_2 bit_69_2 bitb_69_2 word69_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_2 q_70_2 qb_70_2 bit_70_2 bitb_70_2 word70_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_2 q_71_2 qb_71_2 bit_71_2 bitb_71_2 word71_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_2 q_72_2 qb_72_2 bit_72_2 bitb_72_2 word72_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_2 q_73_2 qb_73_2 bit_73_2 bitb_73_2 word73_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_2 q_74_2 qb_74_2 bit_74_2 bitb_74_2 word74_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_2 q_75_2 qb_75_2 bit_75_2 bitb_75_2 word75_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_2 q_76_2 qb_76_2 bit_76_2 bitb_76_2 word76_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_2 q_77_2 qb_77_2 bit_77_2 bitb_77_2 word77_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_2 q_78_2 qb_78_2 bit_78_2 bitb_78_2 word78_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_2 q_79_2 qb_79_2 bit_79_2 bitb_79_2 word79_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_2 q_80_2 qb_80_2 bit_80_2 bitb_80_2 word80_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_2 q_81_2 qb_81_2 bit_81_2 bitb_81_2 word81_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_2 q_82_2 qb_82_2 bit_82_2 bitb_82_2 word82_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_2 q_83_2 qb_83_2 bit_83_2 bitb_83_2 word83_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_2 q_84_2 qb_84_2 bit_84_2 bitb_84_2 word84_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_2 q_85_2 qb_85_2 bit_85_2 bitb_85_2 word85_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_2 q_86_2 qb_86_2 bit_86_2 bitb_86_2 word86_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_2 q_87_2 qb_87_2 bit_87_2 bitb_87_2 word87_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_2 q_88_2 qb_88_2 bit_88_2 bitb_88_2 word88_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_2 q_89_2 qb_89_2 bit_89_2 bitb_89_2 word89_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_2 q_90_2 qb_90_2 bit_90_2 bitb_90_2 word90_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_2 q_91_2 qb_91_2 bit_91_2 bitb_91_2 word91_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_2 q_92_2 qb_92_2 bit_92_2 bitb_92_2 word92_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_2 q_93_2 qb_93_2 bit_93_2 bitb_93_2 word93_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_2 q_94_2 qb_94_2 bit_94_2 bitb_94_2 word94_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_2 q_95_2 qb_95_2 bit_95_2 bitb_95_2 word95_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_2 q_96_2 qb_96_2 bit_96_2 bitb_96_2 word96_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_2 q_97_2 qb_97_2 bit_97_2 bitb_97_2 word97_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_2 q_98_2 qb_98_2 bit_98_2 bitb_98_2 word98_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_2 q_99_2 qb_99_2 bit_99_2 bitb_99_2 word99_2 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_3 q_0_3 qb_0_3 bit_0_3 bitb_0_3 word0_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_3 q_1_3 qb_1_3 bit_1_3 bitb_1_3 word1_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_3 q_2_3 qb_2_3 bit_2_3 bitb_2_3 word2_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_3 q_3_3 qb_3_3 bit_3_3 bitb_3_3 word3_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_3 q_4_3 qb_4_3 bit_4_3 bitb_4_3 word4_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_3 q_5_3 qb_5_3 bit_5_3 bitb_5_3 word5_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_3 q_6_3 qb_6_3 bit_6_3 bitb_6_3 word6_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_3 q_7_3 qb_7_3 bit_7_3 bitb_7_3 word7_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_3 q_8_3 qb_8_3 bit_8_3 bitb_8_3 word8_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_3 q_9_3 qb_9_3 bit_9_3 bitb_9_3 word9_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_3 q_10_3 qb_10_3 bit_10_3 bitb_10_3 word10_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_3 q_11_3 qb_11_3 bit_11_3 bitb_11_3 word11_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_3 q_12_3 qb_12_3 bit_12_3 bitb_12_3 word12_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_3 q_13_3 qb_13_3 bit_13_3 bitb_13_3 word13_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_3 q_14_3 qb_14_3 bit_14_3 bitb_14_3 word14_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_3 q_15_3 qb_15_3 bit_15_3 bitb_15_3 word15_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_3 q_16_3 qb_16_3 bit_16_3 bitb_16_3 word16_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_3 q_17_3 qb_17_3 bit_17_3 bitb_17_3 word17_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_3 q_18_3 qb_18_3 bit_18_3 bitb_18_3 word18_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_3 q_19_3 qb_19_3 bit_19_3 bitb_19_3 word19_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_3 q_20_3 qb_20_3 bit_20_3 bitb_20_3 word20_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_3 q_21_3 qb_21_3 bit_21_3 bitb_21_3 word21_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_3 q_22_3 qb_22_3 bit_22_3 bitb_22_3 word22_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_3 q_23_3 qb_23_3 bit_23_3 bitb_23_3 word23_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_3 q_24_3 qb_24_3 bit_24_3 bitb_24_3 word24_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_3 q_25_3 qb_25_3 bit_25_3 bitb_25_3 word25_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_3 q_26_3 qb_26_3 bit_26_3 bitb_26_3 word26_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_3 q_27_3 qb_27_3 bit_27_3 bitb_27_3 word27_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_3 q_28_3 qb_28_3 bit_28_3 bitb_28_3 word28_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_3 q_29_3 qb_29_3 bit_29_3 bitb_29_3 word29_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_3 q_30_3 qb_30_3 bit_30_3 bitb_30_3 word30_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_3 q_31_3 qb_31_3 bit_31_3 bitb_31_3 word31_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_3 q_32_3 qb_32_3 bit_32_3 bitb_32_3 word32_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_3 q_33_3 qb_33_3 bit_33_3 bitb_33_3 word33_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_3 q_34_3 qb_34_3 bit_34_3 bitb_34_3 word34_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_3 q_35_3 qb_35_3 bit_35_3 bitb_35_3 word35_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_3 q_36_3 qb_36_3 bit_36_3 bitb_36_3 word36_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_3 q_37_3 qb_37_3 bit_37_3 bitb_37_3 word37_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_3 q_38_3 qb_38_3 bit_38_3 bitb_38_3 word38_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_3 q_39_3 qb_39_3 bit_39_3 bitb_39_3 word39_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_3 q_40_3 qb_40_3 bit_40_3 bitb_40_3 word40_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_3 q_41_3 qb_41_3 bit_41_3 bitb_41_3 word41_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_3 q_42_3 qb_42_3 bit_42_3 bitb_42_3 word42_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_3 q_43_3 qb_43_3 bit_43_3 bitb_43_3 word43_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_3 q_44_3 qb_44_3 bit_44_3 bitb_44_3 word44_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_3 q_45_3 qb_45_3 bit_45_3 bitb_45_3 word45_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_3 q_46_3 qb_46_3 bit_46_3 bitb_46_3 word46_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_3 q_47_3 qb_47_3 bit_47_3 bitb_47_3 word47_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_3 q_48_3 qb_48_3 bit_48_3 bitb_48_3 word48_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_3 q_49_3 qb_49_3 bit_49_3 bitb_49_3 word49_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_3 q_50_3 qb_50_3 bit_50_3 bitb_50_3 word50_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_3 q_51_3 qb_51_3 bit_51_3 bitb_51_3 word51_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_3 q_52_3 qb_52_3 bit_52_3 bitb_52_3 word52_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_3 q_53_3 qb_53_3 bit_53_3 bitb_53_3 word53_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_3 q_54_3 qb_54_3 bit_54_3 bitb_54_3 word54_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_3 q_55_3 qb_55_3 bit_55_3 bitb_55_3 word55_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_3 q_56_3 qb_56_3 bit_56_3 bitb_56_3 word56_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_3 q_57_3 qb_57_3 bit_57_3 bitb_57_3 word57_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_3 q_58_3 qb_58_3 bit_58_3 bitb_58_3 word58_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_3 q_59_3 qb_59_3 bit_59_3 bitb_59_3 word59_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_3 q_60_3 qb_60_3 bit_60_3 bitb_60_3 word60_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_3 q_61_3 qb_61_3 bit_61_3 bitb_61_3 word61_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_3 q_62_3 qb_62_3 bit_62_3 bitb_62_3 word62_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_3 q_63_3 qb_63_3 bit_63_3 bitb_63_3 word63_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_3 q_64_3 qb_64_3 bit_64_3 bitb_64_3 word64_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_3 q_65_3 qb_65_3 bit_65_3 bitb_65_3 word65_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_3 q_66_3 qb_66_3 bit_66_3 bitb_66_3 word66_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_3 q_67_3 qb_67_3 bit_67_3 bitb_67_3 word67_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_3 q_68_3 qb_68_3 bit_68_3 bitb_68_3 word68_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_3 q_69_3 qb_69_3 bit_69_3 bitb_69_3 word69_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_3 q_70_3 qb_70_3 bit_70_3 bitb_70_3 word70_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_3 q_71_3 qb_71_3 bit_71_3 bitb_71_3 word71_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_3 q_72_3 qb_72_3 bit_72_3 bitb_72_3 word72_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_3 q_73_3 qb_73_3 bit_73_3 bitb_73_3 word73_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_3 q_74_3 qb_74_3 bit_74_3 bitb_74_3 word74_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_3 q_75_3 qb_75_3 bit_75_3 bitb_75_3 word75_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_3 q_76_3 qb_76_3 bit_76_3 bitb_76_3 word76_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_3 q_77_3 qb_77_3 bit_77_3 bitb_77_3 word77_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_3 q_78_3 qb_78_3 bit_78_3 bitb_78_3 word78_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_3 q_79_3 qb_79_3 bit_79_3 bitb_79_3 word79_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_3 q_80_3 qb_80_3 bit_80_3 bitb_80_3 word80_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_3 q_81_3 qb_81_3 bit_81_3 bitb_81_3 word81_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_3 q_82_3 qb_82_3 bit_82_3 bitb_82_3 word82_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_3 q_83_3 qb_83_3 bit_83_3 bitb_83_3 word83_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_3 q_84_3 qb_84_3 bit_84_3 bitb_84_3 word84_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_3 q_85_3 qb_85_3 bit_85_3 bitb_85_3 word85_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_3 q_86_3 qb_86_3 bit_86_3 bitb_86_3 word86_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_3 q_87_3 qb_87_3 bit_87_3 bitb_87_3 word87_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_3 q_88_3 qb_88_3 bit_88_3 bitb_88_3 word88_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_3 q_89_3 qb_89_3 bit_89_3 bitb_89_3 word89_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_3 q_90_3 qb_90_3 bit_90_3 bitb_90_3 word90_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_3 q_91_3 qb_91_3 bit_91_3 bitb_91_3 word91_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_3 q_92_3 qb_92_3 bit_92_3 bitb_92_3 word92_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_3 q_93_3 qb_93_3 bit_93_3 bitb_93_3 word93_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_3 q_94_3 qb_94_3 bit_94_3 bitb_94_3 word94_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_3 q_95_3 qb_95_3 bit_95_3 bitb_95_3 word95_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_3 q_96_3 qb_96_3 bit_96_3 bitb_96_3 word96_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_3 q_97_3 qb_97_3 bit_97_3 bitb_97_3 word97_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_3 q_98_3 qb_98_3 bit_98_3 bitb_98_3 word98_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_3 q_99_3 qb_99_3 bit_99_3 bitb_99_3 word99_3 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_4 q_0_4 qb_0_4 bit_0_4 bitb_0_4 word0_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_4 q_1_4 qb_1_4 bit_1_4 bitb_1_4 word1_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_4 q_2_4 qb_2_4 bit_2_4 bitb_2_4 word2_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_4 q_3_4 qb_3_4 bit_3_4 bitb_3_4 word3_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_4 q_4_4 qb_4_4 bit_4_4 bitb_4_4 word4_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_4 q_5_4 qb_5_4 bit_5_4 bitb_5_4 word5_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_4 q_6_4 qb_6_4 bit_6_4 bitb_6_4 word6_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_4 q_7_4 qb_7_4 bit_7_4 bitb_7_4 word7_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_4 q_8_4 qb_8_4 bit_8_4 bitb_8_4 word8_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_4 q_9_4 qb_9_4 bit_9_4 bitb_9_4 word9_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_4 q_10_4 qb_10_4 bit_10_4 bitb_10_4 word10_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_4 q_11_4 qb_11_4 bit_11_4 bitb_11_4 word11_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_4 q_12_4 qb_12_4 bit_12_4 bitb_12_4 word12_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_4 q_13_4 qb_13_4 bit_13_4 bitb_13_4 word13_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_4 q_14_4 qb_14_4 bit_14_4 bitb_14_4 word14_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_4 q_15_4 qb_15_4 bit_15_4 bitb_15_4 word15_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_4 q_16_4 qb_16_4 bit_16_4 bitb_16_4 word16_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_4 q_17_4 qb_17_4 bit_17_4 bitb_17_4 word17_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_4 q_18_4 qb_18_4 bit_18_4 bitb_18_4 word18_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_4 q_19_4 qb_19_4 bit_19_4 bitb_19_4 word19_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_4 q_20_4 qb_20_4 bit_20_4 bitb_20_4 word20_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_4 q_21_4 qb_21_4 bit_21_4 bitb_21_4 word21_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_4 q_22_4 qb_22_4 bit_22_4 bitb_22_4 word22_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_4 q_23_4 qb_23_4 bit_23_4 bitb_23_4 word23_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_4 q_24_4 qb_24_4 bit_24_4 bitb_24_4 word24_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_4 q_25_4 qb_25_4 bit_25_4 bitb_25_4 word25_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_4 q_26_4 qb_26_4 bit_26_4 bitb_26_4 word26_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_4 q_27_4 qb_27_4 bit_27_4 bitb_27_4 word27_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_4 q_28_4 qb_28_4 bit_28_4 bitb_28_4 word28_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_4 q_29_4 qb_29_4 bit_29_4 bitb_29_4 word29_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_4 q_30_4 qb_30_4 bit_30_4 bitb_30_4 word30_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_4 q_31_4 qb_31_4 bit_31_4 bitb_31_4 word31_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_4 q_32_4 qb_32_4 bit_32_4 bitb_32_4 word32_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_4 q_33_4 qb_33_4 bit_33_4 bitb_33_4 word33_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_4 q_34_4 qb_34_4 bit_34_4 bitb_34_4 word34_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_4 q_35_4 qb_35_4 bit_35_4 bitb_35_4 word35_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_4 q_36_4 qb_36_4 bit_36_4 bitb_36_4 word36_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_4 q_37_4 qb_37_4 bit_37_4 bitb_37_4 word37_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_4 q_38_4 qb_38_4 bit_38_4 bitb_38_4 word38_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_4 q_39_4 qb_39_4 bit_39_4 bitb_39_4 word39_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_4 q_40_4 qb_40_4 bit_40_4 bitb_40_4 word40_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_4 q_41_4 qb_41_4 bit_41_4 bitb_41_4 word41_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_4 q_42_4 qb_42_4 bit_42_4 bitb_42_4 word42_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_4 q_43_4 qb_43_4 bit_43_4 bitb_43_4 word43_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_4 q_44_4 qb_44_4 bit_44_4 bitb_44_4 word44_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_4 q_45_4 qb_45_4 bit_45_4 bitb_45_4 word45_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_4 q_46_4 qb_46_4 bit_46_4 bitb_46_4 word46_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_4 q_47_4 qb_47_4 bit_47_4 bitb_47_4 word47_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_4 q_48_4 qb_48_4 bit_48_4 bitb_48_4 word48_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_4 q_49_4 qb_49_4 bit_49_4 bitb_49_4 word49_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_4 q_50_4 qb_50_4 bit_50_4 bitb_50_4 word50_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_4 q_51_4 qb_51_4 bit_51_4 bitb_51_4 word51_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_4 q_52_4 qb_52_4 bit_52_4 bitb_52_4 word52_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_4 q_53_4 qb_53_4 bit_53_4 bitb_53_4 word53_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_4 q_54_4 qb_54_4 bit_54_4 bitb_54_4 word54_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_4 q_55_4 qb_55_4 bit_55_4 bitb_55_4 word55_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_4 q_56_4 qb_56_4 bit_56_4 bitb_56_4 word56_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_4 q_57_4 qb_57_4 bit_57_4 bitb_57_4 word57_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_4 q_58_4 qb_58_4 bit_58_4 bitb_58_4 word58_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_4 q_59_4 qb_59_4 bit_59_4 bitb_59_4 word59_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_4 q_60_4 qb_60_4 bit_60_4 bitb_60_4 word60_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_4 q_61_4 qb_61_4 bit_61_4 bitb_61_4 word61_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_4 q_62_4 qb_62_4 bit_62_4 bitb_62_4 word62_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_4 q_63_4 qb_63_4 bit_63_4 bitb_63_4 word63_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_4 q_64_4 qb_64_4 bit_64_4 bitb_64_4 word64_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_4 q_65_4 qb_65_4 bit_65_4 bitb_65_4 word65_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_4 q_66_4 qb_66_4 bit_66_4 bitb_66_4 word66_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_4 q_67_4 qb_67_4 bit_67_4 bitb_67_4 word67_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_4 q_68_4 qb_68_4 bit_68_4 bitb_68_4 word68_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_4 q_69_4 qb_69_4 bit_69_4 bitb_69_4 word69_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_4 q_70_4 qb_70_4 bit_70_4 bitb_70_4 word70_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_4 q_71_4 qb_71_4 bit_71_4 bitb_71_4 word71_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_4 q_72_4 qb_72_4 bit_72_4 bitb_72_4 word72_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_4 q_73_4 qb_73_4 bit_73_4 bitb_73_4 word73_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_4 q_74_4 qb_74_4 bit_74_4 bitb_74_4 word74_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_4 q_75_4 qb_75_4 bit_75_4 bitb_75_4 word75_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_4 q_76_4 qb_76_4 bit_76_4 bitb_76_4 word76_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_4 q_77_4 qb_77_4 bit_77_4 bitb_77_4 word77_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_4 q_78_4 qb_78_4 bit_78_4 bitb_78_4 word78_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_4 q_79_4 qb_79_4 bit_79_4 bitb_79_4 word79_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_4 q_80_4 qb_80_4 bit_80_4 bitb_80_4 word80_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_4 q_81_4 qb_81_4 bit_81_4 bitb_81_4 word81_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_4 q_82_4 qb_82_4 bit_82_4 bitb_82_4 word82_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_4 q_83_4 qb_83_4 bit_83_4 bitb_83_4 word83_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_4 q_84_4 qb_84_4 bit_84_4 bitb_84_4 word84_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_4 q_85_4 qb_85_4 bit_85_4 bitb_85_4 word85_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_4 q_86_4 qb_86_4 bit_86_4 bitb_86_4 word86_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_4 q_87_4 qb_87_4 bit_87_4 bitb_87_4 word87_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_4 q_88_4 qb_88_4 bit_88_4 bitb_88_4 word88_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_4 q_89_4 qb_89_4 bit_89_4 bitb_89_4 word89_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_4 q_90_4 qb_90_4 bit_90_4 bitb_90_4 word90_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_4 q_91_4 qb_91_4 bit_91_4 bitb_91_4 word91_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_4 q_92_4 qb_92_4 bit_92_4 bitb_92_4 word92_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_4 q_93_4 qb_93_4 bit_93_4 bitb_93_4 word93_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_4 q_94_4 qb_94_4 bit_94_4 bitb_94_4 word94_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_4 q_95_4 qb_95_4 bit_95_4 bitb_95_4 word95_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_4 q_96_4 qb_96_4 bit_96_4 bitb_96_4 word96_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_4 q_97_4 qb_97_4 bit_97_4 bitb_97_4 word97_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_4 q_98_4 qb_98_4 bit_98_4 bitb_98_4 word98_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_4 q_99_4 qb_99_4 bit_99_4 bitb_99_4 word99_4 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_5 q_0_5 qb_0_5 bit_0_5 bitb_0_5 word0_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_5 q_1_5 qb_1_5 bit_1_5 bitb_1_5 word1_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_5 q_2_5 qb_2_5 bit_2_5 bitb_2_5 word2_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_5 q_3_5 qb_3_5 bit_3_5 bitb_3_5 word3_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_5 q_4_5 qb_4_5 bit_4_5 bitb_4_5 word4_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_5 q_5_5 qb_5_5 bit_5_5 bitb_5_5 word5_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_5 q_6_5 qb_6_5 bit_6_5 bitb_6_5 word6_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_5 q_7_5 qb_7_5 bit_7_5 bitb_7_5 word7_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_5 q_8_5 qb_8_5 bit_8_5 bitb_8_5 word8_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_5 q_9_5 qb_9_5 bit_9_5 bitb_9_5 word9_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_5 q_10_5 qb_10_5 bit_10_5 bitb_10_5 word10_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_5 q_11_5 qb_11_5 bit_11_5 bitb_11_5 word11_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_5 q_12_5 qb_12_5 bit_12_5 bitb_12_5 word12_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_5 q_13_5 qb_13_5 bit_13_5 bitb_13_5 word13_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_5 q_14_5 qb_14_5 bit_14_5 bitb_14_5 word14_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_5 q_15_5 qb_15_5 bit_15_5 bitb_15_5 word15_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_5 q_16_5 qb_16_5 bit_16_5 bitb_16_5 word16_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_5 q_17_5 qb_17_5 bit_17_5 bitb_17_5 word17_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_5 q_18_5 qb_18_5 bit_18_5 bitb_18_5 word18_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_5 q_19_5 qb_19_5 bit_19_5 bitb_19_5 word19_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_5 q_20_5 qb_20_5 bit_20_5 bitb_20_5 word20_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_5 q_21_5 qb_21_5 bit_21_5 bitb_21_5 word21_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_5 q_22_5 qb_22_5 bit_22_5 bitb_22_5 word22_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_5 q_23_5 qb_23_5 bit_23_5 bitb_23_5 word23_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_5 q_24_5 qb_24_5 bit_24_5 bitb_24_5 word24_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_5 q_25_5 qb_25_5 bit_25_5 bitb_25_5 word25_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_5 q_26_5 qb_26_5 bit_26_5 bitb_26_5 word26_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_5 q_27_5 qb_27_5 bit_27_5 bitb_27_5 word27_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_5 q_28_5 qb_28_5 bit_28_5 bitb_28_5 word28_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_5 q_29_5 qb_29_5 bit_29_5 bitb_29_5 word29_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_5 q_30_5 qb_30_5 bit_30_5 bitb_30_5 word30_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_5 q_31_5 qb_31_5 bit_31_5 bitb_31_5 word31_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_5 q_32_5 qb_32_5 bit_32_5 bitb_32_5 word32_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_5 q_33_5 qb_33_5 bit_33_5 bitb_33_5 word33_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_5 q_34_5 qb_34_5 bit_34_5 bitb_34_5 word34_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_5 q_35_5 qb_35_5 bit_35_5 bitb_35_5 word35_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_5 q_36_5 qb_36_5 bit_36_5 bitb_36_5 word36_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_5 q_37_5 qb_37_5 bit_37_5 bitb_37_5 word37_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_5 q_38_5 qb_38_5 bit_38_5 bitb_38_5 word38_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_5 q_39_5 qb_39_5 bit_39_5 bitb_39_5 word39_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_5 q_40_5 qb_40_5 bit_40_5 bitb_40_5 word40_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_5 q_41_5 qb_41_5 bit_41_5 bitb_41_5 word41_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_5 q_42_5 qb_42_5 bit_42_5 bitb_42_5 word42_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_5 q_43_5 qb_43_5 bit_43_5 bitb_43_5 word43_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_5 q_44_5 qb_44_5 bit_44_5 bitb_44_5 word44_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_5 q_45_5 qb_45_5 bit_45_5 bitb_45_5 word45_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_5 q_46_5 qb_46_5 bit_46_5 bitb_46_5 word46_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_5 q_47_5 qb_47_5 bit_47_5 bitb_47_5 word47_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_5 q_48_5 qb_48_5 bit_48_5 bitb_48_5 word48_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_5 q_49_5 qb_49_5 bit_49_5 bitb_49_5 word49_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_5 q_50_5 qb_50_5 bit_50_5 bitb_50_5 word50_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_5 q_51_5 qb_51_5 bit_51_5 bitb_51_5 word51_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_5 q_52_5 qb_52_5 bit_52_5 bitb_52_5 word52_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_5 q_53_5 qb_53_5 bit_53_5 bitb_53_5 word53_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_5 q_54_5 qb_54_5 bit_54_5 bitb_54_5 word54_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_5 q_55_5 qb_55_5 bit_55_5 bitb_55_5 word55_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_5 q_56_5 qb_56_5 bit_56_5 bitb_56_5 word56_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_5 q_57_5 qb_57_5 bit_57_5 bitb_57_5 word57_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_5 q_58_5 qb_58_5 bit_58_5 bitb_58_5 word58_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_5 q_59_5 qb_59_5 bit_59_5 bitb_59_5 word59_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_5 q_60_5 qb_60_5 bit_60_5 bitb_60_5 word60_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_5 q_61_5 qb_61_5 bit_61_5 bitb_61_5 word61_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_5 q_62_5 qb_62_5 bit_62_5 bitb_62_5 word62_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_5 q_63_5 qb_63_5 bit_63_5 bitb_63_5 word63_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_5 q_64_5 qb_64_5 bit_64_5 bitb_64_5 word64_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_5 q_65_5 qb_65_5 bit_65_5 bitb_65_5 word65_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_5 q_66_5 qb_66_5 bit_66_5 bitb_66_5 word66_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_5 q_67_5 qb_67_5 bit_67_5 bitb_67_5 word67_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_5 q_68_5 qb_68_5 bit_68_5 bitb_68_5 word68_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_5 q_69_5 qb_69_5 bit_69_5 bitb_69_5 word69_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_5 q_70_5 qb_70_5 bit_70_5 bitb_70_5 word70_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_5 q_71_5 qb_71_5 bit_71_5 bitb_71_5 word71_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_5 q_72_5 qb_72_5 bit_72_5 bitb_72_5 word72_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_5 q_73_5 qb_73_5 bit_73_5 bitb_73_5 word73_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_5 q_74_5 qb_74_5 bit_74_5 bitb_74_5 word74_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_5 q_75_5 qb_75_5 bit_75_5 bitb_75_5 word75_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_5 q_76_5 qb_76_5 bit_76_5 bitb_76_5 word76_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_5 q_77_5 qb_77_5 bit_77_5 bitb_77_5 word77_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_5 q_78_5 qb_78_5 bit_78_5 bitb_78_5 word78_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_5 q_79_5 qb_79_5 bit_79_5 bitb_79_5 word79_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_5 q_80_5 qb_80_5 bit_80_5 bitb_80_5 word80_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_5 q_81_5 qb_81_5 bit_81_5 bitb_81_5 word81_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_5 q_82_5 qb_82_5 bit_82_5 bitb_82_5 word82_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_5 q_83_5 qb_83_5 bit_83_5 bitb_83_5 word83_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_5 q_84_5 qb_84_5 bit_84_5 bitb_84_5 word84_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_5 q_85_5 qb_85_5 bit_85_5 bitb_85_5 word85_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_5 q_86_5 qb_86_5 bit_86_5 bitb_86_5 word86_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_5 q_87_5 qb_87_5 bit_87_5 bitb_87_5 word87_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_5 q_88_5 qb_88_5 bit_88_5 bitb_88_5 word88_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_5 q_89_5 qb_89_5 bit_89_5 bitb_89_5 word89_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_5 q_90_5 qb_90_5 bit_90_5 bitb_90_5 word90_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_5 q_91_5 qb_91_5 bit_91_5 bitb_91_5 word91_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_5 q_92_5 qb_92_5 bit_92_5 bitb_92_5 word92_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_5 q_93_5 qb_93_5 bit_93_5 bitb_93_5 word93_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_5 q_94_5 qb_94_5 bit_94_5 bitb_94_5 word94_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_5 q_95_5 qb_95_5 bit_95_5 bitb_95_5 word95_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_5 q_96_5 qb_96_5 bit_96_5 bitb_96_5 word96_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_5 q_97_5 qb_97_5 bit_97_5 bitb_97_5 word97_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_5 q_98_5 qb_98_5 bit_98_5 bitb_98_5 word98_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_5 q_99_5 qb_99_5 bit_99_5 bitb_99_5 word99_5 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_6 q_0_6 qb_0_6 bit_0_6 bitb_0_6 word0_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_6 q_1_6 qb_1_6 bit_1_6 bitb_1_6 word1_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_6 q_2_6 qb_2_6 bit_2_6 bitb_2_6 word2_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_6 q_3_6 qb_3_6 bit_3_6 bitb_3_6 word3_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_6 q_4_6 qb_4_6 bit_4_6 bitb_4_6 word4_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_6 q_5_6 qb_5_6 bit_5_6 bitb_5_6 word5_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_6 q_6_6 qb_6_6 bit_6_6 bitb_6_6 word6_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_6 q_7_6 qb_7_6 bit_7_6 bitb_7_6 word7_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_6 q_8_6 qb_8_6 bit_8_6 bitb_8_6 word8_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_6 q_9_6 qb_9_6 bit_9_6 bitb_9_6 word9_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_6 q_10_6 qb_10_6 bit_10_6 bitb_10_6 word10_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_6 q_11_6 qb_11_6 bit_11_6 bitb_11_6 word11_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_6 q_12_6 qb_12_6 bit_12_6 bitb_12_6 word12_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_6 q_13_6 qb_13_6 bit_13_6 bitb_13_6 word13_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_6 q_14_6 qb_14_6 bit_14_6 bitb_14_6 word14_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_6 q_15_6 qb_15_6 bit_15_6 bitb_15_6 word15_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_6 q_16_6 qb_16_6 bit_16_6 bitb_16_6 word16_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_6 q_17_6 qb_17_6 bit_17_6 bitb_17_6 word17_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_6 q_18_6 qb_18_6 bit_18_6 bitb_18_6 word18_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_6 q_19_6 qb_19_6 bit_19_6 bitb_19_6 word19_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_6 q_20_6 qb_20_6 bit_20_6 bitb_20_6 word20_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_6 q_21_6 qb_21_6 bit_21_6 bitb_21_6 word21_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_6 q_22_6 qb_22_6 bit_22_6 bitb_22_6 word22_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_6 q_23_6 qb_23_6 bit_23_6 bitb_23_6 word23_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_6 q_24_6 qb_24_6 bit_24_6 bitb_24_6 word24_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_6 q_25_6 qb_25_6 bit_25_6 bitb_25_6 word25_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_6 q_26_6 qb_26_6 bit_26_6 bitb_26_6 word26_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_6 q_27_6 qb_27_6 bit_27_6 bitb_27_6 word27_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_6 q_28_6 qb_28_6 bit_28_6 bitb_28_6 word28_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_6 q_29_6 qb_29_6 bit_29_6 bitb_29_6 word29_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_6 q_30_6 qb_30_6 bit_30_6 bitb_30_6 word30_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_6 q_31_6 qb_31_6 bit_31_6 bitb_31_6 word31_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_6 q_32_6 qb_32_6 bit_32_6 bitb_32_6 word32_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_6 q_33_6 qb_33_6 bit_33_6 bitb_33_6 word33_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_6 q_34_6 qb_34_6 bit_34_6 bitb_34_6 word34_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_6 q_35_6 qb_35_6 bit_35_6 bitb_35_6 word35_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_6 q_36_6 qb_36_6 bit_36_6 bitb_36_6 word36_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_6 q_37_6 qb_37_6 bit_37_6 bitb_37_6 word37_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_6 q_38_6 qb_38_6 bit_38_6 bitb_38_6 word38_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_6 q_39_6 qb_39_6 bit_39_6 bitb_39_6 word39_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_6 q_40_6 qb_40_6 bit_40_6 bitb_40_6 word40_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_6 q_41_6 qb_41_6 bit_41_6 bitb_41_6 word41_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_6 q_42_6 qb_42_6 bit_42_6 bitb_42_6 word42_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_6 q_43_6 qb_43_6 bit_43_6 bitb_43_6 word43_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_6 q_44_6 qb_44_6 bit_44_6 bitb_44_6 word44_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_6 q_45_6 qb_45_6 bit_45_6 bitb_45_6 word45_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_6 q_46_6 qb_46_6 bit_46_6 bitb_46_6 word46_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_6 q_47_6 qb_47_6 bit_47_6 bitb_47_6 word47_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_6 q_48_6 qb_48_6 bit_48_6 bitb_48_6 word48_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_6 q_49_6 qb_49_6 bit_49_6 bitb_49_6 word49_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_6 q_50_6 qb_50_6 bit_50_6 bitb_50_6 word50_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_6 q_51_6 qb_51_6 bit_51_6 bitb_51_6 word51_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_6 q_52_6 qb_52_6 bit_52_6 bitb_52_6 word52_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_6 q_53_6 qb_53_6 bit_53_6 bitb_53_6 word53_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_6 q_54_6 qb_54_6 bit_54_6 bitb_54_6 word54_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_6 q_55_6 qb_55_6 bit_55_6 bitb_55_6 word55_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_6 q_56_6 qb_56_6 bit_56_6 bitb_56_6 word56_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_6 q_57_6 qb_57_6 bit_57_6 bitb_57_6 word57_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_6 q_58_6 qb_58_6 bit_58_6 bitb_58_6 word58_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_6 q_59_6 qb_59_6 bit_59_6 bitb_59_6 word59_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_6 q_60_6 qb_60_6 bit_60_6 bitb_60_6 word60_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_6 q_61_6 qb_61_6 bit_61_6 bitb_61_6 word61_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_6 q_62_6 qb_62_6 bit_62_6 bitb_62_6 word62_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_6 q_63_6 qb_63_6 bit_63_6 bitb_63_6 word63_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_6 q_64_6 qb_64_6 bit_64_6 bitb_64_6 word64_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_6 q_65_6 qb_65_6 bit_65_6 bitb_65_6 word65_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_6 q_66_6 qb_66_6 bit_66_6 bitb_66_6 word66_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_6 q_67_6 qb_67_6 bit_67_6 bitb_67_6 word67_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_6 q_68_6 qb_68_6 bit_68_6 bitb_68_6 word68_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_6 q_69_6 qb_69_6 bit_69_6 bitb_69_6 word69_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_6 q_70_6 qb_70_6 bit_70_6 bitb_70_6 word70_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_6 q_71_6 qb_71_6 bit_71_6 bitb_71_6 word71_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_6 q_72_6 qb_72_6 bit_72_6 bitb_72_6 word72_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_6 q_73_6 qb_73_6 bit_73_6 bitb_73_6 word73_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_6 q_74_6 qb_74_6 bit_74_6 bitb_74_6 word74_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_6 q_75_6 qb_75_6 bit_75_6 bitb_75_6 word75_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_6 q_76_6 qb_76_6 bit_76_6 bitb_76_6 word76_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_6 q_77_6 qb_77_6 bit_77_6 bitb_77_6 word77_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_6 q_78_6 qb_78_6 bit_78_6 bitb_78_6 word78_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_6 q_79_6 qb_79_6 bit_79_6 bitb_79_6 word79_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_6 q_80_6 qb_80_6 bit_80_6 bitb_80_6 word80_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_6 q_81_6 qb_81_6 bit_81_6 bitb_81_6 word81_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_6 q_82_6 qb_82_6 bit_82_6 bitb_82_6 word82_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_6 q_83_6 qb_83_6 bit_83_6 bitb_83_6 word83_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_6 q_84_6 qb_84_6 bit_84_6 bitb_84_6 word84_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_6 q_85_6 qb_85_6 bit_85_6 bitb_85_6 word85_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_6 q_86_6 qb_86_6 bit_86_6 bitb_86_6 word86_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_6 q_87_6 qb_87_6 bit_87_6 bitb_87_6 word87_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_6 q_88_6 qb_88_6 bit_88_6 bitb_88_6 word88_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_6 q_89_6 qb_89_6 bit_89_6 bitb_89_6 word89_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_6 q_90_6 qb_90_6 bit_90_6 bitb_90_6 word90_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_6 q_91_6 qb_91_6 bit_91_6 bitb_91_6 word91_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_6 q_92_6 qb_92_6 bit_92_6 bitb_92_6 word92_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_6 q_93_6 qb_93_6 bit_93_6 bitb_93_6 word93_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_6 q_94_6 qb_94_6 bit_94_6 bitb_94_6 word94_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_6 q_95_6 qb_95_6 bit_95_6 bitb_95_6 word95_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_6 q_96_6 qb_96_6 bit_96_6 bitb_96_6 word96_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_6 q_97_6 qb_97_6 bit_97_6 bitb_97_6 word97_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_6 q_98_6 qb_98_6 bit_98_6 bitb_98_6 word98_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_6 q_99_6 qb_99_6 bit_99_6 bitb_99_6 word99_6 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_7 q_0_7 qb_0_7 bit_0_7 bitb_0_7 word0_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_7 q_1_7 qb_1_7 bit_1_7 bitb_1_7 word1_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_7 q_2_7 qb_2_7 bit_2_7 bitb_2_7 word2_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_7 q_3_7 qb_3_7 bit_3_7 bitb_3_7 word3_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_7 q_4_7 qb_4_7 bit_4_7 bitb_4_7 word4_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_7 q_5_7 qb_5_7 bit_5_7 bitb_5_7 word5_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_7 q_6_7 qb_6_7 bit_6_7 bitb_6_7 word6_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_7 q_7_7 qb_7_7 bit_7_7 bitb_7_7 word7_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_7 q_8_7 qb_8_7 bit_8_7 bitb_8_7 word8_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_7 q_9_7 qb_9_7 bit_9_7 bitb_9_7 word9_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_7 q_10_7 qb_10_7 bit_10_7 bitb_10_7 word10_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_7 q_11_7 qb_11_7 bit_11_7 bitb_11_7 word11_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_7 q_12_7 qb_12_7 bit_12_7 bitb_12_7 word12_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_7 q_13_7 qb_13_7 bit_13_7 bitb_13_7 word13_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_7 q_14_7 qb_14_7 bit_14_7 bitb_14_7 word14_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_7 q_15_7 qb_15_7 bit_15_7 bitb_15_7 word15_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_7 q_16_7 qb_16_7 bit_16_7 bitb_16_7 word16_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_7 q_17_7 qb_17_7 bit_17_7 bitb_17_7 word17_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_7 q_18_7 qb_18_7 bit_18_7 bitb_18_7 word18_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_7 q_19_7 qb_19_7 bit_19_7 bitb_19_7 word19_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_7 q_20_7 qb_20_7 bit_20_7 bitb_20_7 word20_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_7 q_21_7 qb_21_7 bit_21_7 bitb_21_7 word21_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_7 q_22_7 qb_22_7 bit_22_7 bitb_22_7 word22_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_7 q_23_7 qb_23_7 bit_23_7 bitb_23_7 word23_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_7 q_24_7 qb_24_7 bit_24_7 bitb_24_7 word24_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_7 q_25_7 qb_25_7 bit_25_7 bitb_25_7 word25_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_7 q_26_7 qb_26_7 bit_26_7 bitb_26_7 word26_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_7 q_27_7 qb_27_7 bit_27_7 bitb_27_7 word27_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_7 q_28_7 qb_28_7 bit_28_7 bitb_28_7 word28_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_7 q_29_7 qb_29_7 bit_29_7 bitb_29_7 word29_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_7 q_30_7 qb_30_7 bit_30_7 bitb_30_7 word30_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_7 q_31_7 qb_31_7 bit_31_7 bitb_31_7 word31_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_7 q_32_7 qb_32_7 bit_32_7 bitb_32_7 word32_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_7 q_33_7 qb_33_7 bit_33_7 bitb_33_7 word33_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_7 q_34_7 qb_34_7 bit_34_7 bitb_34_7 word34_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_7 q_35_7 qb_35_7 bit_35_7 bitb_35_7 word35_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_7 q_36_7 qb_36_7 bit_36_7 bitb_36_7 word36_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_7 q_37_7 qb_37_7 bit_37_7 bitb_37_7 word37_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_7 q_38_7 qb_38_7 bit_38_7 bitb_38_7 word38_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_7 q_39_7 qb_39_7 bit_39_7 bitb_39_7 word39_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_7 q_40_7 qb_40_7 bit_40_7 bitb_40_7 word40_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_7 q_41_7 qb_41_7 bit_41_7 bitb_41_7 word41_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_7 q_42_7 qb_42_7 bit_42_7 bitb_42_7 word42_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_7 q_43_7 qb_43_7 bit_43_7 bitb_43_7 word43_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_7 q_44_7 qb_44_7 bit_44_7 bitb_44_7 word44_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_7 q_45_7 qb_45_7 bit_45_7 bitb_45_7 word45_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_7 q_46_7 qb_46_7 bit_46_7 bitb_46_7 word46_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_7 q_47_7 qb_47_7 bit_47_7 bitb_47_7 word47_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_7 q_48_7 qb_48_7 bit_48_7 bitb_48_7 word48_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_7 q_49_7 qb_49_7 bit_49_7 bitb_49_7 word49_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_7 q_50_7 qb_50_7 bit_50_7 bitb_50_7 word50_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_7 q_51_7 qb_51_7 bit_51_7 bitb_51_7 word51_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_7 q_52_7 qb_52_7 bit_52_7 bitb_52_7 word52_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_7 q_53_7 qb_53_7 bit_53_7 bitb_53_7 word53_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_7 q_54_7 qb_54_7 bit_54_7 bitb_54_7 word54_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_7 q_55_7 qb_55_7 bit_55_7 bitb_55_7 word55_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_7 q_56_7 qb_56_7 bit_56_7 bitb_56_7 word56_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_7 q_57_7 qb_57_7 bit_57_7 bitb_57_7 word57_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_7 q_58_7 qb_58_7 bit_58_7 bitb_58_7 word58_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_7 q_59_7 qb_59_7 bit_59_7 bitb_59_7 word59_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_7 q_60_7 qb_60_7 bit_60_7 bitb_60_7 word60_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_7 q_61_7 qb_61_7 bit_61_7 bitb_61_7 word61_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_7 q_62_7 qb_62_7 bit_62_7 bitb_62_7 word62_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_7 q_63_7 qb_63_7 bit_63_7 bitb_63_7 word63_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_7 q_64_7 qb_64_7 bit_64_7 bitb_64_7 word64_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_7 q_65_7 qb_65_7 bit_65_7 bitb_65_7 word65_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_7 q_66_7 qb_66_7 bit_66_7 bitb_66_7 word66_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_7 q_67_7 qb_67_7 bit_67_7 bitb_67_7 word67_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_7 q_68_7 qb_68_7 bit_68_7 bitb_68_7 word68_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_7 q_69_7 qb_69_7 bit_69_7 bitb_69_7 word69_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_7 q_70_7 qb_70_7 bit_70_7 bitb_70_7 word70_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_7 q_71_7 qb_71_7 bit_71_7 bitb_71_7 word71_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_7 q_72_7 qb_72_7 bit_72_7 bitb_72_7 word72_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_7 q_73_7 qb_73_7 bit_73_7 bitb_73_7 word73_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_7 q_74_7 qb_74_7 bit_74_7 bitb_74_7 word74_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_7 q_75_7 qb_75_7 bit_75_7 bitb_75_7 word75_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_7 q_76_7 qb_76_7 bit_76_7 bitb_76_7 word76_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_7 q_77_7 qb_77_7 bit_77_7 bitb_77_7 word77_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_7 q_78_7 qb_78_7 bit_78_7 bitb_78_7 word78_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_7 q_79_7 qb_79_7 bit_79_7 bitb_79_7 word79_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_7 q_80_7 qb_80_7 bit_80_7 bitb_80_7 word80_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_7 q_81_7 qb_81_7 bit_81_7 bitb_81_7 word81_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_7 q_82_7 qb_82_7 bit_82_7 bitb_82_7 word82_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_7 q_83_7 qb_83_7 bit_83_7 bitb_83_7 word83_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_7 q_84_7 qb_84_7 bit_84_7 bitb_84_7 word84_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_7 q_85_7 qb_85_7 bit_85_7 bitb_85_7 word85_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_7 q_86_7 qb_86_7 bit_86_7 bitb_86_7 word86_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_7 q_87_7 qb_87_7 bit_87_7 bitb_87_7 word87_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_7 q_88_7 qb_88_7 bit_88_7 bitb_88_7 word88_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_7 q_89_7 qb_89_7 bit_89_7 bitb_89_7 word89_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_7 q_90_7 qb_90_7 bit_90_7 bitb_90_7 word90_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_7 q_91_7 qb_91_7 bit_91_7 bitb_91_7 word91_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_7 q_92_7 qb_92_7 bit_92_7 bitb_92_7 word92_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_7 q_93_7 qb_93_7 bit_93_7 bitb_93_7 word93_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_7 q_94_7 qb_94_7 bit_94_7 bitb_94_7 word94_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_7 q_95_7 qb_95_7 bit_95_7 bitb_95_7 word95_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_7 q_96_7 qb_96_7 bit_96_7 bitb_96_7 word96_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_7 q_97_7 qb_97_7 bit_97_7 bitb_97_7 word97_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_7 q_98_7 qb_98_7 bit_98_7 bitb_98_7 word98_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_7 q_99_7 qb_99_7 bit_99_7 bitb_99_7 word99_7 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_8 q_0_8 qb_0_8 bit_0_8 bitb_0_8 word0_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_8 q_1_8 qb_1_8 bit_1_8 bitb_1_8 word1_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_8 q_2_8 qb_2_8 bit_2_8 bitb_2_8 word2_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_8 q_3_8 qb_3_8 bit_3_8 bitb_3_8 word3_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_8 q_4_8 qb_4_8 bit_4_8 bitb_4_8 word4_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_8 q_5_8 qb_5_8 bit_5_8 bitb_5_8 word5_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_8 q_6_8 qb_6_8 bit_6_8 bitb_6_8 word6_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_8 q_7_8 qb_7_8 bit_7_8 bitb_7_8 word7_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_8 q_8_8 qb_8_8 bit_8_8 bitb_8_8 word8_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_8 q_9_8 qb_9_8 bit_9_8 bitb_9_8 word9_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_8 q_10_8 qb_10_8 bit_10_8 bitb_10_8 word10_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_8 q_11_8 qb_11_8 bit_11_8 bitb_11_8 word11_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_8 q_12_8 qb_12_8 bit_12_8 bitb_12_8 word12_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_8 q_13_8 qb_13_8 bit_13_8 bitb_13_8 word13_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_8 q_14_8 qb_14_8 bit_14_8 bitb_14_8 word14_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_8 q_15_8 qb_15_8 bit_15_8 bitb_15_8 word15_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_8 q_16_8 qb_16_8 bit_16_8 bitb_16_8 word16_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_8 q_17_8 qb_17_8 bit_17_8 bitb_17_8 word17_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_8 q_18_8 qb_18_8 bit_18_8 bitb_18_8 word18_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_8 q_19_8 qb_19_8 bit_19_8 bitb_19_8 word19_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_8 q_20_8 qb_20_8 bit_20_8 bitb_20_8 word20_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_8 q_21_8 qb_21_8 bit_21_8 bitb_21_8 word21_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_8 q_22_8 qb_22_8 bit_22_8 bitb_22_8 word22_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_8 q_23_8 qb_23_8 bit_23_8 bitb_23_8 word23_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_8 q_24_8 qb_24_8 bit_24_8 bitb_24_8 word24_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_8 q_25_8 qb_25_8 bit_25_8 bitb_25_8 word25_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_8 q_26_8 qb_26_8 bit_26_8 bitb_26_8 word26_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_8 q_27_8 qb_27_8 bit_27_8 bitb_27_8 word27_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_8 q_28_8 qb_28_8 bit_28_8 bitb_28_8 word28_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_8 q_29_8 qb_29_8 bit_29_8 bitb_29_8 word29_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_8 q_30_8 qb_30_8 bit_30_8 bitb_30_8 word30_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_8 q_31_8 qb_31_8 bit_31_8 bitb_31_8 word31_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_8 q_32_8 qb_32_8 bit_32_8 bitb_32_8 word32_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_8 q_33_8 qb_33_8 bit_33_8 bitb_33_8 word33_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_8 q_34_8 qb_34_8 bit_34_8 bitb_34_8 word34_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_8 q_35_8 qb_35_8 bit_35_8 bitb_35_8 word35_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_8 q_36_8 qb_36_8 bit_36_8 bitb_36_8 word36_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_8 q_37_8 qb_37_8 bit_37_8 bitb_37_8 word37_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_8 q_38_8 qb_38_8 bit_38_8 bitb_38_8 word38_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_8 q_39_8 qb_39_8 bit_39_8 bitb_39_8 word39_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_8 q_40_8 qb_40_8 bit_40_8 bitb_40_8 word40_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_8 q_41_8 qb_41_8 bit_41_8 bitb_41_8 word41_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_8 q_42_8 qb_42_8 bit_42_8 bitb_42_8 word42_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_8 q_43_8 qb_43_8 bit_43_8 bitb_43_8 word43_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_8 q_44_8 qb_44_8 bit_44_8 bitb_44_8 word44_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_8 q_45_8 qb_45_8 bit_45_8 bitb_45_8 word45_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_8 q_46_8 qb_46_8 bit_46_8 bitb_46_8 word46_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_8 q_47_8 qb_47_8 bit_47_8 bitb_47_8 word47_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_8 q_48_8 qb_48_8 bit_48_8 bitb_48_8 word48_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_8 q_49_8 qb_49_8 bit_49_8 bitb_49_8 word49_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_8 q_50_8 qb_50_8 bit_50_8 bitb_50_8 word50_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_8 q_51_8 qb_51_8 bit_51_8 bitb_51_8 word51_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_8 q_52_8 qb_52_8 bit_52_8 bitb_52_8 word52_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_8 q_53_8 qb_53_8 bit_53_8 bitb_53_8 word53_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_8 q_54_8 qb_54_8 bit_54_8 bitb_54_8 word54_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_8 q_55_8 qb_55_8 bit_55_8 bitb_55_8 word55_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_8 q_56_8 qb_56_8 bit_56_8 bitb_56_8 word56_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_8 q_57_8 qb_57_8 bit_57_8 bitb_57_8 word57_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_8 q_58_8 qb_58_8 bit_58_8 bitb_58_8 word58_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_8 q_59_8 qb_59_8 bit_59_8 bitb_59_8 word59_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_8 q_60_8 qb_60_8 bit_60_8 bitb_60_8 word60_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_8 q_61_8 qb_61_8 bit_61_8 bitb_61_8 word61_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_8 q_62_8 qb_62_8 bit_62_8 bitb_62_8 word62_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_8 q_63_8 qb_63_8 bit_63_8 bitb_63_8 word63_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_8 q_64_8 qb_64_8 bit_64_8 bitb_64_8 word64_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_8 q_65_8 qb_65_8 bit_65_8 bitb_65_8 word65_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_8 q_66_8 qb_66_8 bit_66_8 bitb_66_8 word66_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_8 q_67_8 qb_67_8 bit_67_8 bitb_67_8 word67_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_8 q_68_8 qb_68_8 bit_68_8 bitb_68_8 word68_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_8 q_69_8 qb_69_8 bit_69_8 bitb_69_8 word69_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_8 q_70_8 qb_70_8 bit_70_8 bitb_70_8 word70_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_8 q_71_8 qb_71_8 bit_71_8 bitb_71_8 word71_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_8 q_72_8 qb_72_8 bit_72_8 bitb_72_8 word72_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_8 q_73_8 qb_73_8 bit_73_8 bitb_73_8 word73_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_8 q_74_8 qb_74_8 bit_74_8 bitb_74_8 word74_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_8 q_75_8 qb_75_8 bit_75_8 bitb_75_8 word75_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_8 q_76_8 qb_76_8 bit_76_8 bitb_76_8 word76_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_8 q_77_8 qb_77_8 bit_77_8 bitb_77_8 word77_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_8 q_78_8 qb_78_8 bit_78_8 bitb_78_8 word78_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_8 q_79_8 qb_79_8 bit_79_8 bitb_79_8 word79_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_8 q_80_8 qb_80_8 bit_80_8 bitb_80_8 word80_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_8 q_81_8 qb_81_8 bit_81_8 bitb_81_8 word81_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_8 q_82_8 qb_82_8 bit_82_8 bitb_82_8 word82_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_8 q_83_8 qb_83_8 bit_83_8 bitb_83_8 word83_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_8 q_84_8 qb_84_8 bit_84_8 bitb_84_8 word84_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_8 q_85_8 qb_85_8 bit_85_8 bitb_85_8 word85_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_8 q_86_8 qb_86_8 bit_86_8 bitb_86_8 word86_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_8 q_87_8 qb_87_8 bit_87_8 bitb_87_8 word87_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_8 q_88_8 qb_88_8 bit_88_8 bitb_88_8 word88_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_8 q_89_8 qb_89_8 bit_89_8 bitb_89_8 word89_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_8 q_90_8 qb_90_8 bit_90_8 bitb_90_8 word90_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_8 q_91_8 qb_91_8 bit_91_8 bitb_91_8 word91_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_8 q_92_8 qb_92_8 bit_92_8 bitb_92_8 word92_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_8 q_93_8 qb_93_8 bit_93_8 bitb_93_8 word93_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_8 q_94_8 qb_94_8 bit_94_8 bitb_94_8 word94_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_8 q_95_8 qb_95_8 bit_95_8 bitb_95_8 word95_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_8 q_96_8 qb_96_8 bit_96_8 bitb_96_8 word96_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_8 q_97_8 qb_97_8 bit_97_8 bitb_97_8 word97_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_8 q_98_8 qb_98_8 bit_98_8 bitb_98_8 word98_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_8 q_99_8 qb_99_8 bit_99_8 bitb_99_8 word99_8 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_9 q_0_9 qb_0_9 bit_0_9 bitb_0_9 word0_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_9 q_1_9 qb_1_9 bit_1_9 bitb_1_9 word1_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_9 q_2_9 qb_2_9 bit_2_9 bitb_2_9 word2_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_9 q_3_9 qb_3_9 bit_3_9 bitb_3_9 word3_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_9 q_4_9 qb_4_9 bit_4_9 bitb_4_9 word4_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_9 q_5_9 qb_5_9 bit_5_9 bitb_5_9 word5_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_9 q_6_9 qb_6_9 bit_6_9 bitb_6_9 word6_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_9 q_7_9 qb_7_9 bit_7_9 bitb_7_9 word7_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_9 q_8_9 qb_8_9 bit_8_9 bitb_8_9 word8_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_9 q_9_9 qb_9_9 bit_9_9 bitb_9_9 word9_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_9 q_10_9 qb_10_9 bit_10_9 bitb_10_9 word10_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_9 q_11_9 qb_11_9 bit_11_9 bitb_11_9 word11_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_9 q_12_9 qb_12_9 bit_12_9 bitb_12_9 word12_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_9 q_13_9 qb_13_9 bit_13_9 bitb_13_9 word13_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_9 q_14_9 qb_14_9 bit_14_9 bitb_14_9 word14_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_9 q_15_9 qb_15_9 bit_15_9 bitb_15_9 word15_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_9 q_16_9 qb_16_9 bit_16_9 bitb_16_9 word16_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_9 q_17_9 qb_17_9 bit_17_9 bitb_17_9 word17_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_9 q_18_9 qb_18_9 bit_18_9 bitb_18_9 word18_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_9 q_19_9 qb_19_9 bit_19_9 bitb_19_9 word19_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_9 q_20_9 qb_20_9 bit_20_9 bitb_20_9 word20_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_9 q_21_9 qb_21_9 bit_21_9 bitb_21_9 word21_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_9 q_22_9 qb_22_9 bit_22_9 bitb_22_9 word22_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_9 q_23_9 qb_23_9 bit_23_9 bitb_23_9 word23_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_9 q_24_9 qb_24_9 bit_24_9 bitb_24_9 word24_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_9 q_25_9 qb_25_9 bit_25_9 bitb_25_9 word25_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_9 q_26_9 qb_26_9 bit_26_9 bitb_26_9 word26_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_9 q_27_9 qb_27_9 bit_27_9 bitb_27_9 word27_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_9 q_28_9 qb_28_9 bit_28_9 bitb_28_9 word28_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_9 q_29_9 qb_29_9 bit_29_9 bitb_29_9 word29_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_9 q_30_9 qb_30_9 bit_30_9 bitb_30_9 word30_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_9 q_31_9 qb_31_9 bit_31_9 bitb_31_9 word31_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_9 q_32_9 qb_32_9 bit_32_9 bitb_32_9 word32_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_9 q_33_9 qb_33_9 bit_33_9 bitb_33_9 word33_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_9 q_34_9 qb_34_9 bit_34_9 bitb_34_9 word34_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_9 q_35_9 qb_35_9 bit_35_9 bitb_35_9 word35_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_9 q_36_9 qb_36_9 bit_36_9 bitb_36_9 word36_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_9 q_37_9 qb_37_9 bit_37_9 bitb_37_9 word37_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_9 q_38_9 qb_38_9 bit_38_9 bitb_38_9 word38_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_9 q_39_9 qb_39_9 bit_39_9 bitb_39_9 word39_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_9 q_40_9 qb_40_9 bit_40_9 bitb_40_9 word40_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_9 q_41_9 qb_41_9 bit_41_9 bitb_41_9 word41_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_9 q_42_9 qb_42_9 bit_42_9 bitb_42_9 word42_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_9 q_43_9 qb_43_9 bit_43_9 bitb_43_9 word43_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_9 q_44_9 qb_44_9 bit_44_9 bitb_44_9 word44_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_9 q_45_9 qb_45_9 bit_45_9 bitb_45_9 word45_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_9 q_46_9 qb_46_9 bit_46_9 bitb_46_9 word46_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_9 q_47_9 qb_47_9 bit_47_9 bitb_47_9 word47_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_9 q_48_9 qb_48_9 bit_48_9 bitb_48_9 word48_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_9 q_49_9 qb_49_9 bit_49_9 bitb_49_9 word49_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_9 q_50_9 qb_50_9 bit_50_9 bitb_50_9 word50_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_9 q_51_9 qb_51_9 bit_51_9 bitb_51_9 word51_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_9 q_52_9 qb_52_9 bit_52_9 bitb_52_9 word52_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_9 q_53_9 qb_53_9 bit_53_9 bitb_53_9 word53_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_9 q_54_9 qb_54_9 bit_54_9 bitb_54_9 word54_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_9 q_55_9 qb_55_9 bit_55_9 bitb_55_9 word55_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_9 q_56_9 qb_56_9 bit_56_9 bitb_56_9 word56_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_9 q_57_9 qb_57_9 bit_57_9 bitb_57_9 word57_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_9 q_58_9 qb_58_9 bit_58_9 bitb_58_9 word58_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_9 q_59_9 qb_59_9 bit_59_9 bitb_59_9 word59_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_9 q_60_9 qb_60_9 bit_60_9 bitb_60_9 word60_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_9 q_61_9 qb_61_9 bit_61_9 bitb_61_9 word61_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_9 q_62_9 qb_62_9 bit_62_9 bitb_62_9 word62_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_9 q_63_9 qb_63_9 bit_63_9 bitb_63_9 word63_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_9 q_64_9 qb_64_9 bit_64_9 bitb_64_9 word64_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_9 q_65_9 qb_65_9 bit_65_9 bitb_65_9 word65_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_9 q_66_9 qb_66_9 bit_66_9 bitb_66_9 word66_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_9 q_67_9 qb_67_9 bit_67_9 bitb_67_9 word67_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_9 q_68_9 qb_68_9 bit_68_9 bitb_68_9 word68_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_9 q_69_9 qb_69_9 bit_69_9 bitb_69_9 word69_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_9 q_70_9 qb_70_9 bit_70_9 bitb_70_9 word70_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_9 q_71_9 qb_71_9 bit_71_9 bitb_71_9 word71_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_9 q_72_9 qb_72_9 bit_72_9 bitb_72_9 word72_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_9 q_73_9 qb_73_9 bit_73_9 bitb_73_9 word73_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_9 q_74_9 qb_74_9 bit_74_9 bitb_74_9 word74_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_9 q_75_9 qb_75_9 bit_75_9 bitb_75_9 word75_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_9 q_76_9 qb_76_9 bit_76_9 bitb_76_9 word76_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_9 q_77_9 qb_77_9 bit_77_9 bitb_77_9 word77_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_9 q_78_9 qb_78_9 bit_78_9 bitb_78_9 word78_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_9 q_79_9 qb_79_9 bit_79_9 bitb_79_9 word79_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_9 q_80_9 qb_80_9 bit_80_9 bitb_80_9 word80_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_9 q_81_9 qb_81_9 bit_81_9 bitb_81_9 word81_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_9 q_82_9 qb_82_9 bit_82_9 bitb_82_9 word82_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_9 q_83_9 qb_83_9 bit_83_9 bitb_83_9 word83_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_9 q_84_9 qb_84_9 bit_84_9 bitb_84_9 word84_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_9 q_85_9 qb_85_9 bit_85_9 bitb_85_9 word85_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_9 q_86_9 qb_86_9 bit_86_9 bitb_86_9 word86_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_9 q_87_9 qb_87_9 bit_87_9 bitb_87_9 word87_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_9 q_88_9 qb_88_9 bit_88_9 bitb_88_9 word88_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_9 q_89_9 qb_89_9 bit_89_9 bitb_89_9 word89_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_9 q_90_9 qb_90_9 bit_90_9 bitb_90_9 word90_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_9 q_91_9 qb_91_9 bit_91_9 bitb_91_9 word91_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_9 q_92_9 qb_92_9 bit_92_9 bitb_92_9 word92_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_9 q_93_9 qb_93_9 bit_93_9 bitb_93_9 word93_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_9 q_94_9 qb_94_9 bit_94_9 bitb_94_9 word94_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_9 q_95_9 qb_95_9 bit_95_9 bitb_95_9 word95_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_9 q_96_9 qb_96_9 bit_96_9 bitb_96_9 word96_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_9 q_97_9 qb_97_9 bit_97_9 bitb_97_9 word97_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_9 q_98_9 qb_98_9 bit_98_9 bitb_98_9 word98_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_9 q_99_9 qb_99_9 bit_99_9 bitb_99_9 word99_9 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_10 q_0_10 qb_0_10 bit_0_10 bitb_0_10 word0_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_10 q_1_10 qb_1_10 bit_1_10 bitb_1_10 word1_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_10 q_2_10 qb_2_10 bit_2_10 bitb_2_10 word2_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_10 q_3_10 qb_3_10 bit_3_10 bitb_3_10 word3_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_10 q_4_10 qb_4_10 bit_4_10 bitb_4_10 word4_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_10 q_5_10 qb_5_10 bit_5_10 bitb_5_10 word5_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_10 q_6_10 qb_6_10 bit_6_10 bitb_6_10 word6_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_10 q_7_10 qb_7_10 bit_7_10 bitb_7_10 word7_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_10 q_8_10 qb_8_10 bit_8_10 bitb_8_10 word8_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_10 q_9_10 qb_9_10 bit_9_10 bitb_9_10 word9_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_10 q_10_10 qb_10_10 bit_10_10 bitb_10_10 word10_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_10 q_11_10 qb_11_10 bit_11_10 bitb_11_10 word11_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_10 q_12_10 qb_12_10 bit_12_10 bitb_12_10 word12_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_10 q_13_10 qb_13_10 bit_13_10 bitb_13_10 word13_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_10 q_14_10 qb_14_10 bit_14_10 bitb_14_10 word14_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_10 q_15_10 qb_15_10 bit_15_10 bitb_15_10 word15_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_10 q_16_10 qb_16_10 bit_16_10 bitb_16_10 word16_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_10 q_17_10 qb_17_10 bit_17_10 bitb_17_10 word17_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_10 q_18_10 qb_18_10 bit_18_10 bitb_18_10 word18_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_10 q_19_10 qb_19_10 bit_19_10 bitb_19_10 word19_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_10 q_20_10 qb_20_10 bit_20_10 bitb_20_10 word20_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_10 q_21_10 qb_21_10 bit_21_10 bitb_21_10 word21_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_10 q_22_10 qb_22_10 bit_22_10 bitb_22_10 word22_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_10 q_23_10 qb_23_10 bit_23_10 bitb_23_10 word23_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_10 q_24_10 qb_24_10 bit_24_10 bitb_24_10 word24_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_10 q_25_10 qb_25_10 bit_25_10 bitb_25_10 word25_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_10 q_26_10 qb_26_10 bit_26_10 bitb_26_10 word26_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_10 q_27_10 qb_27_10 bit_27_10 bitb_27_10 word27_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_10 q_28_10 qb_28_10 bit_28_10 bitb_28_10 word28_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_10 q_29_10 qb_29_10 bit_29_10 bitb_29_10 word29_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_10 q_30_10 qb_30_10 bit_30_10 bitb_30_10 word30_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_10 q_31_10 qb_31_10 bit_31_10 bitb_31_10 word31_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_10 q_32_10 qb_32_10 bit_32_10 bitb_32_10 word32_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_10 q_33_10 qb_33_10 bit_33_10 bitb_33_10 word33_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_10 q_34_10 qb_34_10 bit_34_10 bitb_34_10 word34_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_10 q_35_10 qb_35_10 bit_35_10 bitb_35_10 word35_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_10 q_36_10 qb_36_10 bit_36_10 bitb_36_10 word36_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_10 q_37_10 qb_37_10 bit_37_10 bitb_37_10 word37_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_10 q_38_10 qb_38_10 bit_38_10 bitb_38_10 word38_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_10 q_39_10 qb_39_10 bit_39_10 bitb_39_10 word39_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_10 q_40_10 qb_40_10 bit_40_10 bitb_40_10 word40_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_10 q_41_10 qb_41_10 bit_41_10 bitb_41_10 word41_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_10 q_42_10 qb_42_10 bit_42_10 bitb_42_10 word42_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_10 q_43_10 qb_43_10 bit_43_10 bitb_43_10 word43_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_10 q_44_10 qb_44_10 bit_44_10 bitb_44_10 word44_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_10 q_45_10 qb_45_10 bit_45_10 bitb_45_10 word45_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_10 q_46_10 qb_46_10 bit_46_10 bitb_46_10 word46_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_10 q_47_10 qb_47_10 bit_47_10 bitb_47_10 word47_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_10 q_48_10 qb_48_10 bit_48_10 bitb_48_10 word48_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_10 q_49_10 qb_49_10 bit_49_10 bitb_49_10 word49_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_10 q_50_10 qb_50_10 bit_50_10 bitb_50_10 word50_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_10 q_51_10 qb_51_10 bit_51_10 bitb_51_10 word51_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_10 q_52_10 qb_52_10 bit_52_10 bitb_52_10 word52_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_10 q_53_10 qb_53_10 bit_53_10 bitb_53_10 word53_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_10 q_54_10 qb_54_10 bit_54_10 bitb_54_10 word54_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_10 q_55_10 qb_55_10 bit_55_10 bitb_55_10 word55_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_10 q_56_10 qb_56_10 bit_56_10 bitb_56_10 word56_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_10 q_57_10 qb_57_10 bit_57_10 bitb_57_10 word57_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_10 q_58_10 qb_58_10 bit_58_10 bitb_58_10 word58_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_10 q_59_10 qb_59_10 bit_59_10 bitb_59_10 word59_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_10 q_60_10 qb_60_10 bit_60_10 bitb_60_10 word60_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_10 q_61_10 qb_61_10 bit_61_10 bitb_61_10 word61_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_10 q_62_10 qb_62_10 bit_62_10 bitb_62_10 word62_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_10 q_63_10 qb_63_10 bit_63_10 bitb_63_10 word63_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_10 q_64_10 qb_64_10 bit_64_10 bitb_64_10 word64_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_10 q_65_10 qb_65_10 bit_65_10 bitb_65_10 word65_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_10 q_66_10 qb_66_10 bit_66_10 bitb_66_10 word66_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_10 q_67_10 qb_67_10 bit_67_10 bitb_67_10 word67_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_10 q_68_10 qb_68_10 bit_68_10 bitb_68_10 word68_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_10 q_69_10 qb_69_10 bit_69_10 bitb_69_10 word69_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_10 q_70_10 qb_70_10 bit_70_10 bitb_70_10 word70_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_10 q_71_10 qb_71_10 bit_71_10 bitb_71_10 word71_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_10 q_72_10 qb_72_10 bit_72_10 bitb_72_10 word72_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_10 q_73_10 qb_73_10 bit_73_10 bitb_73_10 word73_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_10 q_74_10 qb_74_10 bit_74_10 bitb_74_10 word74_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_10 q_75_10 qb_75_10 bit_75_10 bitb_75_10 word75_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_10 q_76_10 qb_76_10 bit_76_10 bitb_76_10 word76_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_10 q_77_10 qb_77_10 bit_77_10 bitb_77_10 word77_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_10 q_78_10 qb_78_10 bit_78_10 bitb_78_10 word78_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_10 q_79_10 qb_79_10 bit_79_10 bitb_79_10 word79_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_10 q_80_10 qb_80_10 bit_80_10 bitb_80_10 word80_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_10 q_81_10 qb_81_10 bit_81_10 bitb_81_10 word81_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_10 q_82_10 qb_82_10 bit_82_10 bitb_82_10 word82_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_10 q_83_10 qb_83_10 bit_83_10 bitb_83_10 word83_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_10 q_84_10 qb_84_10 bit_84_10 bitb_84_10 word84_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_10 q_85_10 qb_85_10 bit_85_10 bitb_85_10 word85_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_10 q_86_10 qb_86_10 bit_86_10 bitb_86_10 word86_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_10 q_87_10 qb_87_10 bit_87_10 bitb_87_10 word87_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_10 q_88_10 qb_88_10 bit_88_10 bitb_88_10 word88_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_10 q_89_10 qb_89_10 bit_89_10 bitb_89_10 word89_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_10 q_90_10 qb_90_10 bit_90_10 bitb_90_10 word90_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_10 q_91_10 qb_91_10 bit_91_10 bitb_91_10 word91_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_10 q_92_10 qb_92_10 bit_92_10 bitb_92_10 word92_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_10 q_93_10 qb_93_10 bit_93_10 bitb_93_10 word93_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_10 q_94_10 qb_94_10 bit_94_10 bitb_94_10 word94_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_10 q_95_10 qb_95_10 bit_95_10 bitb_95_10 word95_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_10 q_96_10 qb_96_10 bit_96_10 bitb_96_10 word96_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_10 q_97_10 qb_97_10 bit_97_10 bitb_97_10 word97_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_10 q_98_10 qb_98_10 bit_98_10 bitb_98_10 word98_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_10 q_99_10 qb_99_10 bit_99_10 bitb_99_10 word99_10 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_11 q_0_11 qb_0_11 bit_0_11 bitb_0_11 word0_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_11 q_1_11 qb_1_11 bit_1_11 bitb_1_11 word1_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_11 q_2_11 qb_2_11 bit_2_11 bitb_2_11 word2_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_11 q_3_11 qb_3_11 bit_3_11 bitb_3_11 word3_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_11 q_4_11 qb_4_11 bit_4_11 bitb_4_11 word4_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_11 q_5_11 qb_5_11 bit_5_11 bitb_5_11 word5_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_11 q_6_11 qb_6_11 bit_6_11 bitb_6_11 word6_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_11 q_7_11 qb_7_11 bit_7_11 bitb_7_11 word7_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_11 q_8_11 qb_8_11 bit_8_11 bitb_8_11 word8_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_11 q_9_11 qb_9_11 bit_9_11 bitb_9_11 word9_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_11 q_10_11 qb_10_11 bit_10_11 bitb_10_11 word10_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_11 q_11_11 qb_11_11 bit_11_11 bitb_11_11 word11_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_11 q_12_11 qb_12_11 bit_12_11 bitb_12_11 word12_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_11 q_13_11 qb_13_11 bit_13_11 bitb_13_11 word13_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_11 q_14_11 qb_14_11 bit_14_11 bitb_14_11 word14_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_11 q_15_11 qb_15_11 bit_15_11 bitb_15_11 word15_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_11 q_16_11 qb_16_11 bit_16_11 bitb_16_11 word16_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_11 q_17_11 qb_17_11 bit_17_11 bitb_17_11 word17_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_11 q_18_11 qb_18_11 bit_18_11 bitb_18_11 word18_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_11 q_19_11 qb_19_11 bit_19_11 bitb_19_11 word19_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_11 q_20_11 qb_20_11 bit_20_11 bitb_20_11 word20_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_11 q_21_11 qb_21_11 bit_21_11 bitb_21_11 word21_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_11 q_22_11 qb_22_11 bit_22_11 bitb_22_11 word22_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_11 q_23_11 qb_23_11 bit_23_11 bitb_23_11 word23_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_11 q_24_11 qb_24_11 bit_24_11 bitb_24_11 word24_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_11 q_25_11 qb_25_11 bit_25_11 bitb_25_11 word25_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_11 q_26_11 qb_26_11 bit_26_11 bitb_26_11 word26_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_11 q_27_11 qb_27_11 bit_27_11 bitb_27_11 word27_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_11 q_28_11 qb_28_11 bit_28_11 bitb_28_11 word28_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_11 q_29_11 qb_29_11 bit_29_11 bitb_29_11 word29_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_11 q_30_11 qb_30_11 bit_30_11 bitb_30_11 word30_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_11 q_31_11 qb_31_11 bit_31_11 bitb_31_11 word31_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_11 q_32_11 qb_32_11 bit_32_11 bitb_32_11 word32_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_11 q_33_11 qb_33_11 bit_33_11 bitb_33_11 word33_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_11 q_34_11 qb_34_11 bit_34_11 bitb_34_11 word34_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_11 q_35_11 qb_35_11 bit_35_11 bitb_35_11 word35_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_11 q_36_11 qb_36_11 bit_36_11 bitb_36_11 word36_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_11 q_37_11 qb_37_11 bit_37_11 bitb_37_11 word37_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_11 q_38_11 qb_38_11 bit_38_11 bitb_38_11 word38_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_11 q_39_11 qb_39_11 bit_39_11 bitb_39_11 word39_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_11 q_40_11 qb_40_11 bit_40_11 bitb_40_11 word40_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_11 q_41_11 qb_41_11 bit_41_11 bitb_41_11 word41_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_11 q_42_11 qb_42_11 bit_42_11 bitb_42_11 word42_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_11 q_43_11 qb_43_11 bit_43_11 bitb_43_11 word43_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_11 q_44_11 qb_44_11 bit_44_11 bitb_44_11 word44_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_11 q_45_11 qb_45_11 bit_45_11 bitb_45_11 word45_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_11 q_46_11 qb_46_11 bit_46_11 bitb_46_11 word46_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_11 q_47_11 qb_47_11 bit_47_11 bitb_47_11 word47_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_11 q_48_11 qb_48_11 bit_48_11 bitb_48_11 word48_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_11 q_49_11 qb_49_11 bit_49_11 bitb_49_11 word49_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_11 q_50_11 qb_50_11 bit_50_11 bitb_50_11 word50_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_11 q_51_11 qb_51_11 bit_51_11 bitb_51_11 word51_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_11 q_52_11 qb_52_11 bit_52_11 bitb_52_11 word52_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_11 q_53_11 qb_53_11 bit_53_11 bitb_53_11 word53_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_11 q_54_11 qb_54_11 bit_54_11 bitb_54_11 word54_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_11 q_55_11 qb_55_11 bit_55_11 bitb_55_11 word55_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_11 q_56_11 qb_56_11 bit_56_11 bitb_56_11 word56_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_11 q_57_11 qb_57_11 bit_57_11 bitb_57_11 word57_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_11 q_58_11 qb_58_11 bit_58_11 bitb_58_11 word58_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_11 q_59_11 qb_59_11 bit_59_11 bitb_59_11 word59_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_11 q_60_11 qb_60_11 bit_60_11 bitb_60_11 word60_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_11 q_61_11 qb_61_11 bit_61_11 bitb_61_11 word61_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_11 q_62_11 qb_62_11 bit_62_11 bitb_62_11 word62_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_11 q_63_11 qb_63_11 bit_63_11 bitb_63_11 word63_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_11 q_64_11 qb_64_11 bit_64_11 bitb_64_11 word64_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_11 q_65_11 qb_65_11 bit_65_11 bitb_65_11 word65_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_11 q_66_11 qb_66_11 bit_66_11 bitb_66_11 word66_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_11 q_67_11 qb_67_11 bit_67_11 bitb_67_11 word67_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_11 q_68_11 qb_68_11 bit_68_11 bitb_68_11 word68_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_11 q_69_11 qb_69_11 bit_69_11 bitb_69_11 word69_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_11 q_70_11 qb_70_11 bit_70_11 bitb_70_11 word70_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_11 q_71_11 qb_71_11 bit_71_11 bitb_71_11 word71_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_11 q_72_11 qb_72_11 bit_72_11 bitb_72_11 word72_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_11 q_73_11 qb_73_11 bit_73_11 bitb_73_11 word73_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_11 q_74_11 qb_74_11 bit_74_11 bitb_74_11 word74_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_11 q_75_11 qb_75_11 bit_75_11 bitb_75_11 word75_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_11 q_76_11 qb_76_11 bit_76_11 bitb_76_11 word76_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_11 q_77_11 qb_77_11 bit_77_11 bitb_77_11 word77_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_11 q_78_11 qb_78_11 bit_78_11 bitb_78_11 word78_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_11 q_79_11 qb_79_11 bit_79_11 bitb_79_11 word79_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_11 q_80_11 qb_80_11 bit_80_11 bitb_80_11 word80_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_11 q_81_11 qb_81_11 bit_81_11 bitb_81_11 word81_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_11 q_82_11 qb_82_11 bit_82_11 bitb_82_11 word82_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_11 q_83_11 qb_83_11 bit_83_11 bitb_83_11 word83_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_11 q_84_11 qb_84_11 bit_84_11 bitb_84_11 word84_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_11 q_85_11 qb_85_11 bit_85_11 bitb_85_11 word85_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_11 q_86_11 qb_86_11 bit_86_11 bitb_86_11 word86_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_11 q_87_11 qb_87_11 bit_87_11 bitb_87_11 word87_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_11 q_88_11 qb_88_11 bit_88_11 bitb_88_11 word88_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_11 q_89_11 qb_89_11 bit_89_11 bitb_89_11 word89_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_11 q_90_11 qb_90_11 bit_90_11 bitb_90_11 word90_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_11 q_91_11 qb_91_11 bit_91_11 bitb_91_11 word91_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_11 q_92_11 qb_92_11 bit_92_11 bitb_92_11 word92_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_11 q_93_11 qb_93_11 bit_93_11 bitb_93_11 word93_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_11 q_94_11 qb_94_11 bit_94_11 bitb_94_11 word94_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_11 q_95_11 qb_95_11 bit_95_11 bitb_95_11 word95_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_11 q_96_11 qb_96_11 bit_96_11 bitb_96_11 word96_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_11 q_97_11 qb_97_11 bit_97_11 bitb_97_11 word97_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_11 q_98_11 qb_98_11 bit_98_11 bitb_98_11 word98_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_11 q_99_11 qb_99_11 bit_99_11 bitb_99_11 word99_11 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_12 q_0_12 qb_0_12 bit_0_12 bitb_0_12 word0_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_12 q_1_12 qb_1_12 bit_1_12 bitb_1_12 word1_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_12 q_2_12 qb_2_12 bit_2_12 bitb_2_12 word2_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_12 q_3_12 qb_3_12 bit_3_12 bitb_3_12 word3_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_12 q_4_12 qb_4_12 bit_4_12 bitb_4_12 word4_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_12 q_5_12 qb_5_12 bit_5_12 bitb_5_12 word5_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_12 q_6_12 qb_6_12 bit_6_12 bitb_6_12 word6_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_12 q_7_12 qb_7_12 bit_7_12 bitb_7_12 word7_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_12 q_8_12 qb_8_12 bit_8_12 bitb_8_12 word8_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_12 q_9_12 qb_9_12 bit_9_12 bitb_9_12 word9_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_12 q_10_12 qb_10_12 bit_10_12 bitb_10_12 word10_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_12 q_11_12 qb_11_12 bit_11_12 bitb_11_12 word11_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_12 q_12_12 qb_12_12 bit_12_12 bitb_12_12 word12_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_12 q_13_12 qb_13_12 bit_13_12 bitb_13_12 word13_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_12 q_14_12 qb_14_12 bit_14_12 bitb_14_12 word14_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_12 q_15_12 qb_15_12 bit_15_12 bitb_15_12 word15_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_12 q_16_12 qb_16_12 bit_16_12 bitb_16_12 word16_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_12 q_17_12 qb_17_12 bit_17_12 bitb_17_12 word17_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_12 q_18_12 qb_18_12 bit_18_12 bitb_18_12 word18_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_12 q_19_12 qb_19_12 bit_19_12 bitb_19_12 word19_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_12 q_20_12 qb_20_12 bit_20_12 bitb_20_12 word20_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_12 q_21_12 qb_21_12 bit_21_12 bitb_21_12 word21_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_12 q_22_12 qb_22_12 bit_22_12 bitb_22_12 word22_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_12 q_23_12 qb_23_12 bit_23_12 bitb_23_12 word23_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_12 q_24_12 qb_24_12 bit_24_12 bitb_24_12 word24_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_12 q_25_12 qb_25_12 bit_25_12 bitb_25_12 word25_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_12 q_26_12 qb_26_12 bit_26_12 bitb_26_12 word26_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_12 q_27_12 qb_27_12 bit_27_12 bitb_27_12 word27_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_12 q_28_12 qb_28_12 bit_28_12 bitb_28_12 word28_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_12 q_29_12 qb_29_12 bit_29_12 bitb_29_12 word29_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_12 q_30_12 qb_30_12 bit_30_12 bitb_30_12 word30_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_12 q_31_12 qb_31_12 bit_31_12 bitb_31_12 word31_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_12 q_32_12 qb_32_12 bit_32_12 bitb_32_12 word32_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_12 q_33_12 qb_33_12 bit_33_12 bitb_33_12 word33_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_12 q_34_12 qb_34_12 bit_34_12 bitb_34_12 word34_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_12 q_35_12 qb_35_12 bit_35_12 bitb_35_12 word35_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_12 q_36_12 qb_36_12 bit_36_12 bitb_36_12 word36_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_12 q_37_12 qb_37_12 bit_37_12 bitb_37_12 word37_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_12 q_38_12 qb_38_12 bit_38_12 bitb_38_12 word38_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_12 q_39_12 qb_39_12 bit_39_12 bitb_39_12 word39_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_12 q_40_12 qb_40_12 bit_40_12 bitb_40_12 word40_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_12 q_41_12 qb_41_12 bit_41_12 bitb_41_12 word41_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_12 q_42_12 qb_42_12 bit_42_12 bitb_42_12 word42_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_12 q_43_12 qb_43_12 bit_43_12 bitb_43_12 word43_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_12 q_44_12 qb_44_12 bit_44_12 bitb_44_12 word44_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_12 q_45_12 qb_45_12 bit_45_12 bitb_45_12 word45_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_12 q_46_12 qb_46_12 bit_46_12 bitb_46_12 word46_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_12 q_47_12 qb_47_12 bit_47_12 bitb_47_12 word47_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_12 q_48_12 qb_48_12 bit_48_12 bitb_48_12 word48_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_12 q_49_12 qb_49_12 bit_49_12 bitb_49_12 word49_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_12 q_50_12 qb_50_12 bit_50_12 bitb_50_12 word50_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_12 q_51_12 qb_51_12 bit_51_12 bitb_51_12 word51_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_12 q_52_12 qb_52_12 bit_52_12 bitb_52_12 word52_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_12 q_53_12 qb_53_12 bit_53_12 bitb_53_12 word53_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_12 q_54_12 qb_54_12 bit_54_12 bitb_54_12 word54_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_12 q_55_12 qb_55_12 bit_55_12 bitb_55_12 word55_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_12 q_56_12 qb_56_12 bit_56_12 bitb_56_12 word56_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_12 q_57_12 qb_57_12 bit_57_12 bitb_57_12 word57_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_12 q_58_12 qb_58_12 bit_58_12 bitb_58_12 word58_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_12 q_59_12 qb_59_12 bit_59_12 bitb_59_12 word59_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_12 q_60_12 qb_60_12 bit_60_12 bitb_60_12 word60_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_12 q_61_12 qb_61_12 bit_61_12 bitb_61_12 word61_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_12 q_62_12 qb_62_12 bit_62_12 bitb_62_12 word62_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_12 q_63_12 qb_63_12 bit_63_12 bitb_63_12 word63_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_12 q_64_12 qb_64_12 bit_64_12 bitb_64_12 word64_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_12 q_65_12 qb_65_12 bit_65_12 bitb_65_12 word65_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_12 q_66_12 qb_66_12 bit_66_12 bitb_66_12 word66_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_12 q_67_12 qb_67_12 bit_67_12 bitb_67_12 word67_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_12 q_68_12 qb_68_12 bit_68_12 bitb_68_12 word68_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_12 q_69_12 qb_69_12 bit_69_12 bitb_69_12 word69_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_12 q_70_12 qb_70_12 bit_70_12 bitb_70_12 word70_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_12 q_71_12 qb_71_12 bit_71_12 bitb_71_12 word71_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_12 q_72_12 qb_72_12 bit_72_12 bitb_72_12 word72_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_12 q_73_12 qb_73_12 bit_73_12 bitb_73_12 word73_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_12 q_74_12 qb_74_12 bit_74_12 bitb_74_12 word74_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_12 q_75_12 qb_75_12 bit_75_12 bitb_75_12 word75_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_12 q_76_12 qb_76_12 bit_76_12 bitb_76_12 word76_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_12 q_77_12 qb_77_12 bit_77_12 bitb_77_12 word77_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_12 q_78_12 qb_78_12 bit_78_12 bitb_78_12 word78_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_12 q_79_12 qb_79_12 bit_79_12 bitb_79_12 word79_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_12 q_80_12 qb_80_12 bit_80_12 bitb_80_12 word80_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_12 q_81_12 qb_81_12 bit_81_12 bitb_81_12 word81_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_12 q_82_12 qb_82_12 bit_82_12 bitb_82_12 word82_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_12 q_83_12 qb_83_12 bit_83_12 bitb_83_12 word83_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_12 q_84_12 qb_84_12 bit_84_12 bitb_84_12 word84_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_12 q_85_12 qb_85_12 bit_85_12 bitb_85_12 word85_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_12 q_86_12 qb_86_12 bit_86_12 bitb_86_12 word86_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_12 q_87_12 qb_87_12 bit_87_12 bitb_87_12 word87_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_12 q_88_12 qb_88_12 bit_88_12 bitb_88_12 word88_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_12 q_89_12 qb_89_12 bit_89_12 bitb_89_12 word89_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_12 q_90_12 qb_90_12 bit_90_12 bitb_90_12 word90_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_12 q_91_12 qb_91_12 bit_91_12 bitb_91_12 word91_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_12 q_92_12 qb_92_12 bit_92_12 bitb_92_12 word92_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_12 q_93_12 qb_93_12 bit_93_12 bitb_93_12 word93_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_12 q_94_12 qb_94_12 bit_94_12 bitb_94_12 word94_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_12 q_95_12 qb_95_12 bit_95_12 bitb_95_12 word95_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_12 q_96_12 qb_96_12 bit_96_12 bitb_96_12 word96_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_12 q_97_12 qb_97_12 bit_97_12 bitb_97_12 word97_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_12 q_98_12 qb_98_12 bit_98_12 bitb_98_12 word98_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_12 q_99_12 qb_99_12 bit_99_12 bitb_99_12 word99_12 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_13 q_0_13 qb_0_13 bit_0_13 bitb_0_13 word0_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_13 q_1_13 qb_1_13 bit_1_13 bitb_1_13 word1_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_13 q_2_13 qb_2_13 bit_2_13 bitb_2_13 word2_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_13 q_3_13 qb_3_13 bit_3_13 bitb_3_13 word3_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_13 q_4_13 qb_4_13 bit_4_13 bitb_4_13 word4_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_13 q_5_13 qb_5_13 bit_5_13 bitb_5_13 word5_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_13 q_6_13 qb_6_13 bit_6_13 bitb_6_13 word6_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_13 q_7_13 qb_7_13 bit_7_13 bitb_7_13 word7_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_13 q_8_13 qb_8_13 bit_8_13 bitb_8_13 word8_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_13 q_9_13 qb_9_13 bit_9_13 bitb_9_13 word9_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_13 q_10_13 qb_10_13 bit_10_13 bitb_10_13 word10_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_13 q_11_13 qb_11_13 bit_11_13 bitb_11_13 word11_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_13 q_12_13 qb_12_13 bit_12_13 bitb_12_13 word12_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_13 q_13_13 qb_13_13 bit_13_13 bitb_13_13 word13_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_13 q_14_13 qb_14_13 bit_14_13 bitb_14_13 word14_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_13 q_15_13 qb_15_13 bit_15_13 bitb_15_13 word15_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_13 q_16_13 qb_16_13 bit_16_13 bitb_16_13 word16_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_13 q_17_13 qb_17_13 bit_17_13 bitb_17_13 word17_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_13 q_18_13 qb_18_13 bit_18_13 bitb_18_13 word18_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_13 q_19_13 qb_19_13 bit_19_13 bitb_19_13 word19_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_13 q_20_13 qb_20_13 bit_20_13 bitb_20_13 word20_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_13 q_21_13 qb_21_13 bit_21_13 bitb_21_13 word21_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_13 q_22_13 qb_22_13 bit_22_13 bitb_22_13 word22_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_13 q_23_13 qb_23_13 bit_23_13 bitb_23_13 word23_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_13 q_24_13 qb_24_13 bit_24_13 bitb_24_13 word24_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_13 q_25_13 qb_25_13 bit_25_13 bitb_25_13 word25_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_13 q_26_13 qb_26_13 bit_26_13 bitb_26_13 word26_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_13 q_27_13 qb_27_13 bit_27_13 bitb_27_13 word27_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_13 q_28_13 qb_28_13 bit_28_13 bitb_28_13 word28_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_13 q_29_13 qb_29_13 bit_29_13 bitb_29_13 word29_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_13 q_30_13 qb_30_13 bit_30_13 bitb_30_13 word30_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_13 q_31_13 qb_31_13 bit_31_13 bitb_31_13 word31_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_13 q_32_13 qb_32_13 bit_32_13 bitb_32_13 word32_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_13 q_33_13 qb_33_13 bit_33_13 bitb_33_13 word33_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_13 q_34_13 qb_34_13 bit_34_13 bitb_34_13 word34_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_13 q_35_13 qb_35_13 bit_35_13 bitb_35_13 word35_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_13 q_36_13 qb_36_13 bit_36_13 bitb_36_13 word36_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_13 q_37_13 qb_37_13 bit_37_13 bitb_37_13 word37_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_13 q_38_13 qb_38_13 bit_38_13 bitb_38_13 word38_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_13 q_39_13 qb_39_13 bit_39_13 bitb_39_13 word39_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_13 q_40_13 qb_40_13 bit_40_13 bitb_40_13 word40_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_13 q_41_13 qb_41_13 bit_41_13 bitb_41_13 word41_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_13 q_42_13 qb_42_13 bit_42_13 bitb_42_13 word42_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_13 q_43_13 qb_43_13 bit_43_13 bitb_43_13 word43_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_13 q_44_13 qb_44_13 bit_44_13 bitb_44_13 word44_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_13 q_45_13 qb_45_13 bit_45_13 bitb_45_13 word45_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_13 q_46_13 qb_46_13 bit_46_13 bitb_46_13 word46_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_13 q_47_13 qb_47_13 bit_47_13 bitb_47_13 word47_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_13 q_48_13 qb_48_13 bit_48_13 bitb_48_13 word48_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_13 q_49_13 qb_49_13 bit_49_13 bitb_49_13 word49_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_13 q_50_13 qb_50_13 bit_50_13 bitb_50_13 word50_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_13 q_51_13 qb_51_13 bit_51_13 bitb_51_13 word51_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_13 q_52_13 qb_52_13 bit_52_13 bitb_52_13 word52_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_13 q_53_13 qb_53_13 bit_53_13 bitb_53_13 word53_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_13 q_54_13 qb_54_13 bit_54_13 bitb_54_13 word54_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_13 q_55_13 qb_55_13 bit_55_13 bitb_55_13 word55_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_13 q_56_13 qb_56_13 bit_56_13 bitb_56_13 word56_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_13 q_57_13 qb_57_13 bit_57_13 bitb_57_13 word57_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_13 q_58_13 qb_58_13 bit_58_13 bitb_58_13 word58_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_13 q_59_13 qb_59_13 bit_59_13 bitb_59_13 word59_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_13 q_60_13 qb_60_13 bit_60_13 bitb_60_13 word60_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_13 q_61_13 qb_61_13 bit_61_13 bitb_61_13 word61_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_13 q_62_13 qb_62_13 bit_62_13 bitb_62_13 word62_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_13 q_63_13 qb_63_13 bit_63_13 bitb_63_13 word63_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_13 q_64_13 qb_64_13 bit_64_13 bitb_64_13 word64_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_13 q_65_13 qb_65_13 bit_65_13 bitb_65_13 word65_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_13 q_66_13 qb_66_13 bit_66_13 bitb_66_13 word66_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_13 q_67_13 qb_67_13 bit_67_13 bitb_67_13 word67_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_13 q_68_13 qb_68_13 bit_68_13 bitb_68_13 word68_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_13 q_69_13 qb_69_13 bit_69_13 bitb_69_13 word69_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_13 q_70_13 qb_70_13 bit_70_13 bitb_70_13 word70_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_13 q_71_13 qb_71_13 bit_71_13 bitb_71_13 word71_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_13 q_72_13 qb_72_13 bit_72_13 bitb_72_13 word72_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_13 q_73_13 qb_73_13 bit_73_13 bitb_73_13 word73_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_13 q_74_13 qb_74_13 bit_74_13 bitb_74_13 word74_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_13 q_75_13 qb_75_13 bit_75_13 bitb_75_13 word75_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_13 q_76_13 qb_76_13 bit_76_13 bitb_76_13 word76_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_13 q_77_13 qb_77_13 bit_77_13 bitb_77_13 word77_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_13 q_78_13 qb_78_13 bit_78_13 bitb_78_13 word78_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_13 q_79_13 qb_79_13 bit_79_13 bitb_79_13 word79_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_13 q_80_13 qb_80_13 bit_80_13 bitb_80_13 word80_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_13 q_81_13 qb_81_13 bit_81_13 bitb_81_13 word81_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_13 q_82_13 qb_82_13 bit_82_13 bitb_82_13 word82_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_13 q_83_13 qb_83_13 bit_83_13 bitb_83_13 word83_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_13 q_84_13 qb_84_13 bit_84_13 bitb_84_13 word84_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_13 q_85_13 qb_85_13 bit_85_13 bitb_85_13 word85_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_13 q_86_13 qb_86_13 bit_86_13 bitb_86_13 word86_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_13 q_87_13 qb_87_13 bit_87_13 bitb_87_13 word87_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_13 q_88_13 qb_88_13 bit_88_13 bitb_88_13 word88_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_13 q_89_13 qb_89_13 bit_89_13 bitb_89_13 word89_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_13 q_90_13 qb_90_13 bit_90_13 bitb_90_13 word90_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_13 q_91_13 qb_91_13 bit_91_13 bitb_91_13 word91_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_13 q_92_13 qb_92_13 bit_92_13 bitb_92_13 word92_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_13 q_93_13 qb_93_13 bit_93_13 bitb_93_13 word93_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_13 q_94_13 qb_94_13 bit_94_13 bitb_94_13 word94_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_13 q_95_13 qb_95_13 bit_95_13 bitb_95_13 word95_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_13 q_96_13 qb_96_13 bit_96_13 bitb_96_13 word96_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_13 q_97_13 qb_97_13 bit_97_13 bitb_97_13 word97_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_13 q_98_13 qb_98_13 bit_98_13 bitb_98_13 word98_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_13 q_99_13 qb_99_13 bit_99_13 bitb_99_13 word99_13 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_14 q_0_14 qb_0_14 bit_0_14 bitb_0_14 word0_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_14 q_1_14 qb_1_14 bit_1_14 bitb_1_14 word1_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_14 q_2_14 qb_2_14 bit_2_14 bitb_2_14 word2_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_14 q_3_14 qb_3_14 bit_3_14 bitb_3_14 word3_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_14 q_4_14 qb_4_14 bit_4_14 bitb_4_14 word4_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_14 q_5_14 qb_5_14 bit_5_14 bitb_5_14 word5_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_14 q_6_14 qb_6_14 bit_6_14 bitb_6_14 word6_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_14 q_7_14 qb_7_14 bit_7_14 bitb_7_14 word7_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_14 q_8_14 qb_8_14 bit_8_14 bitb_8_14 word8_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_14 q_9_14 qb_9_14 bit_9_14 bitb_9_14 word9_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_14 q_10_14 qb_10_14 bit_10_14 bitb_10_14 word10_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_14 q_11_14 qb_11_14 bit_11_14 bitb_11_14 word11_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_14 q_12_14 qb_12_14 bit_12_14 bitb_12_14 word12_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_14 q_13_14 qb_13_14 bit_13_14 bitb_13_14 word13_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_14 q_14_14 qb_14_14 bit_14_14 bitb_14_14 word14_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_14 q_15_14 qb_15_14 bit_15_14 bitb_15_14 word15_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_14 q_16_14 qb_16_14 bit_16_14 bitb_16_14 word16_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_14 q_17_14 qb_17_14 bit_17_14 bitb_17_14 word17_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_14 q_18_14 qb_18_14 bit_18_14 bitb_18_14 word18_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_14 q_19_14 qb_19_14 bit_19_14 bitb_19_14 word19_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_14 q_20_14 qb_20_14 bit_20_14 bitb_20_14 word20_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_14 q_21_14 qb_21_14 bit_21_14 bitb_21_14 word21_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_14 q_22_14 qb_22_14 bit_22_14 bitb_22_14 word22_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_14 q_23_14 qb_23_14 bit_23_14 bitb_23_14 word23_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_14 q_24_14 qb_24_14 bit_24_14 bitb_24_14 word24_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_14 q_25_14 qb_25_14 bit_25_14 bitb_25_14 word25_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_14 q_26_14 qb_26_14 bit_26_14 bitb_26_14 word26_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_14 q_27_14 qb_27_14 bit_27_14 bitb_27_14 word27_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_14 q_28_14 qb_28_14 bit_28_14 bitb_28_14 word28_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_14 q_29_14 qb_29_14 bit_29_14 bitb_29_14 word29_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_14 q_30_14 qb_30_14 bit_30_14 bitb_30_14 word30_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_14 q_31_14 qb_31_14 bit_31_14 bitb_31_14 word31_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_14 q_32_14 qb_32_14 bit_32_14 bitb_32_14 word32_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_14 q_33_14 qb_33_14 bit_33_14 bitb_33_14 word33_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_14 q_34_14 qb_34_14 bit_34_14 bitb_34_14 word34_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_14 q_35_14 qb_35_14 bit_35_14 bitb_35_14 word35_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_14 q_36_14 qb_36_14 bit_36_14 bitb_36_14 word36_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_14 q_37_14 qb_37_14 bit_37_14 bitb_37_14 word37_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_14 q_38_14 qb_38_14 bit_38_14 bitb_38_14 word38_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_14 q_39_14 qb_39_14 bit_39_14 bitb_39_14 word39_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_14 q_40_14 qb_40_14 bit_40_14 bitb_40_14 word40_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_14 q_41_14 qb_41_14 bit_41_14 bitb_41_14 word41_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_14 q_42_14 qb_42_14 bit_42_14 bitb_42_14 word42_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_14 q_43_14 qb_43_14 bit_43_14 bitb_43_14 word43_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_14 q_44_14 qb_44_14 bit_44_14 bitb_44_14 word44_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_14 q_45_14 qb_45_14 bit_45_14 bitb_45_14 word45_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_14 q_46_14 qb_46_14 bit_46_14 bitb_46_14 word46_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_14 q_47_14 qb_47_14 bit_47_14 bitb_47_14 word47_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_14 q_48_14 qb_48_14 bit_48_14 bitb_48_14 word48_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_14 q_49_14 qb_49_14 bit_49_14 bitb_49_14 word49_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_14 q_50_14 qb_50_14 bit_50_14 bitb_50_14 word50_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_14 q_51_14 qb_51_14 bit_51_14 bitb_51_14 word51_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_14 q_52_14 qb_52_14 bit_52_14 bitb_52_14 word52_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_14 q_53_14 qb_53_14 bit_53_14 bitb_53_14 word53_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_14 q_54_14 qb_54_14 bit_54_14 bitb_54_14 word54_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_14 q_55_14 qb_55_14 bit_55_14 bitb_55_14 word55_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_14 q_56_14 qb_56_14 bit_56_14 bitb_56_14 word56_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_14 q_57_14 qb_57_14 bit_57_14 bitb_57_14 word57_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_14 q_58_14 qb_58_14 bit_58_14 bitb_58_14 word58_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_14 q_59_14 qb_59_14 bit_59_14 bitb_59_14 word59_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_14 q_60_14 qb_60_14 bit_60_14 bitb_60_14 word60_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_14 q_61_14 qb_61_14 bit_61_14 bitb_61_14 word61_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_14 q_62_14 qb_62_14 bit_62_14 bitb_62_14 word62_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_14 q_63_14 qb_63_14 bit_63_14 bitb_63_14 word63_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_14 q_64_14 qb_64_14 bit_64_14 bitb_64_14 word64_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_14 q_65_14 qb_65_14 bit_65_14 bitb_65_14 word65_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_14 q_66_14 qb_66_14 bit_66_14 bitb_66_14 word66_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_14 q_67_14 qb_67_14 bit_67_14 bitb_67_14 word67_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_14 q_68_14 qb_68_14 bit_68_14 bitb_68_14 word68_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_14 q_69_14 qb_69_14 bit_69_14 bitb_69_14 word69_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_14 q_70_14 qb_70_14 bit_70_14 bitb_70_14 word70_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_14 q_71_14 qb_71_14 bit_71_14 bitb_71_14 word71_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_14 q_72_14 qb_72_14 bit_72_14 bitb_72_14 word72_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_14 q_73_14 qb_73_14 bit_73_14 bitb_73_14 word73_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_14 q_74_14 qb_74_14 bit_74_14 bitb_74_14 word74_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_14 q_75_14 qb_75_14 bit_75_14 bitb_75_14 word75_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_14 q_76_14 qb_76_14 bit_76_14 bitb_76_14 word76_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_14 q_77_14 qb_77_14 bit_77_14 bitb_77_14 word77_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_14 q_78_14 qb_78_14 bit_78_14 bitb_78_14 word78_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_14 q_79_14 qb_79_14 bit_79_14 bitb_79_14 word79_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_14 q_80_14 qb_80_14 bit_80_14 bitb_80_14 word80_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_14 q_81_14 qb_81_14 bit_81_14 bitb_81_14 word81_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_14 q_82_14 qb_82_14 bit_82_14 bitb_82_14 word82_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_14 q_83_14 qb_83_14 bit_83_14 bitb_83_14 word83_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_14 q_84_14 qb_84_14 bit_84_14 bitb_84_14 word84_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_14 q_85_14 qb_85_14 bit_85_14 bitb_85_14 word85_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_14 q_86_14 qb_86_14 bit_86_14 bitb_86_14 word86_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_14 q_87_14 qb_87_14 bit_87_14 bitb_87_14 word87_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_14 q_88_14 qb_88_14 bit_88_14 bitb_88_14 word88_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_14 q_89_14 qb_89_14 bit_89_14 bitb_89_14 word89_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_14 q_90_14 qb_90_14 bit_90_14 bitb_90_14 word90_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_14 q_91_14 qb_91_14 bit_91_14 bitb_91_14 word91_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_14 q_92_14 qb_92_14 bit_92_14 bitb_92_14 word92_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_14 q_93_14 qb_93_14 bit_93_14 bitb_93_14 word93_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_14 q_94_14 qb_94_14 bit_94_14 bitb_94_14 word94_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_14 q_95_14 qb_95_14 bit_95_14 bitb_95_14 word95_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_14 q_96_14 qb_96_14 bit_96_14 bitb_96_14 word96_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_14 q_97_14 qb_97_14 bit_97_14 bitb_97_14 word97_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_14 q_98_14 qb_98_14 bit_98_14 bitb_98_14 word98_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_14 q_99_14 qb_99_14 bit_99_14 bitb_99_14 word99_14 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_15 q_0_15 qb_0_15 bit_0_15 bitb_0_15 word0_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_15 q_1_15 qb_1_15 bit_1_15 bitb_1_15 word1_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_15 q_2_15 qb_2_15 bit_2_15 bitb_2_15 word2_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_15 q_3_15 qb_3_15 bit_3_15 bitb_3_15 word3_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_15 q_4_15 qb_4_15 bit_4_15 bitb_4_15 word4_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_15 q_5_15 qb_5_15 bit_5_15 bitb_5_15 word5_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_15 q_6_15 qb_6_15 bit_6_15 bitb_6_15 word6_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_15 q_7_15 qb_7_15 bit_7_15 bitb_7_15 word7_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_15 q_8_15 qb_8_15 bit_8_15 bitb_8_15 word8_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_15 q_9_15 qb_9_15 bit_9_15 bitb_9_15 word9_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_15 q_10_15 qb_10_15 bit_10_15 bitb_10_15 word10_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_15 q_11_15 qb_11_15 bit_11_15 bitb_11_15 word11_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_15 q_12_15 qb_12_15 bit_12_15 bitb_12_15 word12_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_15 q_13_15 qb_13_15 bit_13_15 bitb_13_15 word13_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_15 q_14_15 qb_14_15 bit_14_15 bitb_14_15 word14_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_15 q_15_15 qb_15_15 bit_15_15 bitb_15_15 word15_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_15 q_16_15 qb_16_15 bit_16_15 bitb_16_15 word16_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_15 q_17_15 qb_17_15 bit_17_15 bitb_17_15 word17_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_15 q_18_15 qb_18_15 bit_18_15 bitb_18_15 word18_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_15 q_19_15 qb_19_15 bit_19_15 bitb_19_15 word19_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_15 q_20_15 qb_20_15 bit_20_15 bitb_20_15 word20_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_15 q_21_15 qb_21_15 bit_21_15 bitb_21_15 word21_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_15 q_22_15 qb_22_15 bit_22_15 bitb_22_15 word22_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_15 q_23_15 qb_23_15 bit_23_15 bitb_23_15 word23_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_15 q_24_15 qb_24_15 bit_24_15 bitb_24_15 word24_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_15 q_25_15 qb_25_15 bit_25_15 bitb_25_15 word25_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_15 q_26_15 qb_26_15 bit_26_15 bitb_26_15 word26_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_15 q_27_15 qb_27_15 bit_27_15 bitb_27_15 word27_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_15 q_28_15 qb_28_15 bit_28_15 bitb_28_15 word28_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_15 q_29_15 qb_29_15 bit_29_15 bitb_29_15 word29_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_15 q_30_15 qb_30_15 bit_30_15 bitb_30_15 word30_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_15 q_31_15 qb_31_15 bit_31_15 bitb_31_15 word31_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_15 q_32_15 qb_32_15 bit_32_15 bitb_32_15 word32_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_15 q_33_15 qb_33_15 bit_33_15 bitb_33_15 word33_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_15 q_34_15 qb_34_15 bit_34_15 bitb_34_15 word34_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_15 q_35_15 qb_35_15 bit_35_15 bitb_35_15 word35_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_15 q_36_15 qb_36_15 bit_36_15 bitb_36_15 word36_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_15 q_37_15 qb_37_15 bit_37_15 bitb_37_15 word37_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_15 q_38_15 qb_38_15 bit_38_15 bitb_38_15 word38_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_15 q_39_15 qb_39_15 bit_39_15 bitb_39_15 word39_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_15 q_40_15 qb_40_15 bit_40_15 bitb_40_15 word40_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_15 q_41_15 qb_41_15 bit_41_15 bitb_41_15 word41_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_15 q_42_15 qb_42_15 bit_42_15 bitb_42_15 word42_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_15 q_43_15 qb_43_15 bit_43_15 bitb_43_15 word43_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_15 q_44_15 qb_44_15 bit_44_15 bitb_44_15 word44_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_15 q_45_15 qb_45_15 bit_45_15 bitb_45_15 word45_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_15 q_46_15 qb_46_15 bit_46_15 bitb_46_15 word46_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_15 q_47_15 qb_47_15 bit_47_15 bitb_47_15 word47_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_15 q_48_15 qb_48_15 bit_48_15 bitb_48_15 word48_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_15 q_49_15 qb_49_15 bit_49_15 bitb_49_15 word49_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_15 q_50_15 qb_50_15 bit_50_15 bitb_50_15 word50_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_15 q_51_15 qb_51_15 bit_51_15 bitb_51_15 word51_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_15 q_52_15 qb_52_15 bit_52_15 bitb_52_15 word52_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_15 q_53_15 qb_53_15 bit_53_15 bitb_53_15 word53_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_15 q_54_15 qb_54_15 bit_54_15 bitb_54_15 word54_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_15 q_55_15 qb_55_15 bit_55_15 bitb_55_15 word55_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_15 q_56_15 qb_56_15 bit_56_15 bitb_56_15 word56_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_15 q_57_15 qb_57_15 bit_57_15 bitb_57_15 word57_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_15 q_58_15 qb_58_15 bit_58_15 bitb_58_15 word58_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_15 q_59_15 qb_59_15 bit_59_15 bitb_59_15 word59_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_15 q_60_15 qb_60_15 bit_60_15 bitb_60_15 word60_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_15 q_61_15 qb_61_15 bit_61_15 bitb_61_15 word61_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_15 q_62_15 qb_62_15 bit_62_15 bitb_62_15 word62_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_15 q_63_15 qb_63_15 bit_63_15 bitb_63_15 word63_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_15 q_64_15 qb_64_15 bit_64_15 bitb_64_15 word64_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_15 q_65_15 qb_65_15 bit_65_15 bitb_65_15 word65_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_15 q_66_15 qb_66_15 bit_66_15 bitb_66_15 word66_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_15 q_67_15 qb_67_15 bit_67_15 bitb_67_15 word67_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_15 q_68_15 qb_68_15 bit_68_15 bitb_68_15 word68_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_15 q_69_15 qb_69_15 bit_69_15 bitb_69_15 word69_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_15 q_70_15 qb_70_15 bit_70_15 bitb_70_15 word70_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_15 q_71_15 qb_71_15 bit_71_15 bitb_71_15 word71_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_15 q_72_15 qb_72_15 bit_72_15 bitb_72_15 word72_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_15 q_73_15 qb_73_15 bit_73_15 bitb_73_15 word73_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_15 q_74_15 qb_74_15 bit_74_15 bitb_74_15 word74_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_15 q_75_15 qb_75_15 bit_75_15 bitb_75_15 word75_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_15 q_76_15 qb_76_15 bit_76_15 bitb_76_15 word76_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_15 q_77_15 qb_77_15 bit_77_15 bitb_77_15 word77_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_15 q_78_15 qb_78_15 bit_78_15 bitb_78_15 word78_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_15 q_79_15 qb_79_15 bit_79_15 bitb_79_15 word79_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_15 q_80_15 qb_80_15 bit_80_15 bitb_80_15 word80_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_15 q_81_15 qb_81_15 bit_81_15 bitb_81_15 word81_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_15 q_82_15 qb_82_15 bit_82_15 bitb_82_15 word82_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_15 q_83_15 qb_83_15 bit_83_15 bitb_83_15 word83_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_15 q_84_15 qb_84_15 bit_84_15 bitb_84_15 word84_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_15 q_85_15 qb_85_15 bit_85_15 bitb_85_15 word85_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_15 q_86_15 qb_86_15 bit_86_15 bitb_86_15 word86_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_15 q_87_15 qb_87_15 bit_87_15 bitb_87_15 word87_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_15 q_88_15 qb_88_15 bit_88_15 bitb_88_15 word88_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_15 q_89_15 qb_89_15 bit_89_15 bitb_89_15 word89_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_15 q_90_15 qb_90_15 bit_90_15 bitb_90_15 word90_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_15 q_91_15 qb_91_15 bit_91_15 bitb_91_15 word91_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_15 q_92_15 qb_92_15 bit_92_15 bitb_92_15 word92_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_15 q_93_15 qb_93_15 bit_93_15 bitb_93_15 word93_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_15 q_94_15 qb_94_15 bit_94_15 bitb_94_15 word94_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_15 q_95_15 qb_95_15 bit_95_15 bitb_95_15 word95_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_15 q_96_15 qb_96_15 bit_96_15 bitb_96_15 word96_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_15 q_97_15 qb_97_15 bit_97_15 bitb_97_15 word97_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_15 q_98_15 qb_98_15 bit_98_15 bitb_98_15 word98_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_15 q_99_15 qb_99_15 bit_99_15 bitb_99_15 word99_15 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_16 q_0_16 qb_0_16 bit_0_16 bitb_0_16 word0_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_16 q_1_16 qb_1_16 bit_1_16 bitb_1_16 word1_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_16 q_2_16 qb_2_16 bit_2_16 bitb_2_16 word2_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_16 q_3_16 qb_3_16 bit_3_16 bitb_3_16 word3_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_16 q_4_16 qb_4_16 bit_4_16 bitb_4_16 word4_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_16 q_5_16 qb_5_16 bit_5_16 bitb_5_16 word5_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_16 q_6_16 qb_6_16 bit_6_16 bitb_6_16 word6_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_16 q_7_16 qb_7_16 bit_7_16 bitb_7_16 word7_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_16 q_8_16 qb_8_16 bit_8_16 bitb_8_16 word8_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_16 q_9_16 qb_9_16 bit_9_16 bitb_9_16 word9_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_16 q_10_16 qb_10_16 bit_10_16 bitb_10_16 word10_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_16 q_11_16 qb_11_16 bit_11_16 bitb_11_16 word11_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_16 q_12_16 qb_12_16 bit_12_16 bitb_12_16 word12_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_16 q_13_16 qb_13_16 bit_13_16 bitb_13_16 word13_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_16 q_14_16 qb_14_16 bit_14_16 bitb_14_16 word14_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_16 q_15_16 qb_15_16 bit_15_16 bitb_15_16 word15_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_16 q_16_16 qb_16_16 bit_16_16 bitb_16_16 word16_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_16 q_17_16 qb_17_16 bit_17_16 bitb_17_16 word17_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_16 q_18_16 qb_18_16 bit_18_16 bitb_18_16 word18_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_16 q_19_16 qb_19_16 bit_19_16 bitb_19_16 word19_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_16 q_20_16 qb_20_16 bit_20_16 bitb_20_16 word20_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_16 q_21_16 qb_21_16 bit_21_16 bitb_21_16 word21_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_16 q_22_16 qb_22_16 bit_22_16 bitb_22_16 word22_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_16 q_23_16 qb_23_16 bit_23_16 bitb_23_16 word23_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_16 q_24_16 qb_24_16 bit_24_16 bitb_24_16 word24_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_16 q_25_16 qb_25_16 bit_25_16 bitb_25_16 word25_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_16 q_26_16 qb_26_16 bit_26_16 bitb_26_16 word26_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_16 q_27_16 qb_27_16 bit_27_16 bitb_27_16 word27_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_16 q_28_16 qb_28_16 bit_28_16 bitb_28_16 word28_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_16 q_29_16 qb_29_16 bit_29_16 bitb_29_16 word29_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_16 q_30_16 qb_30_16 bit_30_16 bitb_30_16 word30_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_16 q_31_16 qb_31_16 bit_31_16 bitb_31_16 word31_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_16 q_32_16 qb_32_16 bit_32_16 bitb_32_16 word32_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_16 q_33_16 qb_33_16 bit_33_16 bitb_33_16 word33_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_16 q_34_16 qb_34_16 bit_34_16 bitb_34_16 word34_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_16 q_35_16 qb_35_16 bit_35_16 bitb_35_16 word35_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_16 q_36_16 qb_36_16 bit_36_16 bitb_36_16 word36_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_16 q_37_16 qb_37_16 bit_37_16 bitb_37_16 word37_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_16 q_38_16 qb_38_16 bit_38_16 bitb_38_16 word38_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_16 q_39_16 qb_39_16 bit_39_16 bitb_39_16 word39_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_16 q_40_16 qb_40_16 bit_40_16 bitb_40_16 word40_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_16 q_41_16 qb_41_16 bit_41_16 bitb_41_16 word41_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_16 q_42_16 qb_42_16 bit_42_16 bitb_42_16 word42_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_16 q_43_16 qb_43_16 bit_43_16 bitb_43_16 word43_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_16 q_44_16 qb_44_16 bit_44_16 bitb_44_16 word44_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_16 q_45_16 qb_45_16 bit_45_16 bitb_45_16 word45_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_16 q_46_16 qb_46_16 bit_46_16 bitb_46_16 word46_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_16 q_47_16 qb_47_16 bit_47_16 bitb_47_16 word47_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_16 q_48_16 qb_48_16 bit_48_16 bitb_48_16 word48_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_16 q_49_16 qb_49_16 bit_49_16 bitb_49_16 word49_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_16 q_50_16 qb_50_16 bit_50_16 bitb_50_16 word50_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_16 q_51_16 qb_51_16 bit_51_16 bitb_51_16 word51_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_16 q_52_16 qb_52_16 bit_52_16 bitb_52_16 word52_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_16 q_53_16 qb_53_16 bit_53_16 bitb_53_16 word53_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_16 q_54_16 qb_54_16 bit_54_16 bitb_54_16 word54_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_16 q_55_16 qb_55_16 bit_55_16 bitb_55_16 word55_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_16 q_56_16 qb_56_16 bit_56_16 bitb_56_16 word56_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_16 q_57_16 qb_57_16 bit_57_16 bitb_57_16 word57_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_16 q_58_16 qb_58_16 bit_58_16 bitb_58_16 word58_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_16 q_59_16 qb_59_16 bit_59_16 bitb_59_16 word59_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_16 q_60_16 qb_60_16 bit_60_16 bitb_60_16 word60_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_16 q_61_16 qb_61_16 bit_61_16 bitb_61_16 word61_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_16 q_62_16 qb_62_16 bit_62_16 bitb_62_16 word62_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_16 q_63_16 qb_63_16 bit_63_16 bitb_63_16 word63_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_16 q_64_16 qb_64_16 bit_64_16 bitb_64_16 word64_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_16 q_65_16 qb_65_16 bit_65_16 bitb_65_16 word65_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_16 q_66_16 qb_66_16 bit_66_16 bitb_66_16 word66_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_16 q_67_16 qb_67_16 bit_67_16 bitb_67_16 word67_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_16 q_68_16 qb_68_16 bit_68_16 bitb_68_16 word68_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_16 q_69_16 qb_69_16 bit_69_16 bitb_69_16 word69_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_16 q_70_16 qb_70_16 bit_70_16 bitb_70_16 word70_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_16 q_71_16 qb_71_16 bit_71_16 bitb_71_16 word71_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_16 q_72_16 qb_72_16 bit_72_16 bitb_72_16 word72_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_16 q_73_16 qb_73_16 bit_73_16 bitb_73_16 word73_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_16 q_74_16 qb_74_16 bit_74_16 bitb_74_16 word74_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_16 q_75_16 qb_75_16 bit_75_16 bitb_75_16 word75_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_16 q_76_16 qb_76_16 bit_76_16 bitb_76_16 word76_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_16 q_77_16 qb_77_16 bit_77_16 bitb_77_16 word77_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_16 q_78_16 qb_78_16 bit_78_16 bitb_78_16 word78_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_16 q_79_16 qb_79_16 bit_79_16 bitb_79_16 word79_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_16 q_80_16 qb_80_16 bit_80_16 bitb_80_16 word80_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_16 q_81_16 qb_81_16 bit_81_16 bitb_81_16 word81_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_16 q_82_16 qb_82_16 bit_82_16 bitb_82_16 word82_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_16 q_83_16 qb_83_16 bit_83_16 bitb_83_16 word83_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_16 q_84_16 qb_84_16 bit_84_16 bitb_84_16 word84_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_16 q_85_16 qb_85_16 bit_85_16 bitb_85_16 word85_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_16 q_86_16 qb_86_16 bit_86_16 bitb_86_16 word86_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_16 q_87_16 qb_87_16 bit_87_16 bitb_87_16 word87_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_16 q_88_16 qb_88_16 bit_88_16 bitb_88_16 word88_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_16 q_89_16 qb_89_16 bit_89_16 bitb_89_16 word89_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_16 q_90_16 qb_90_16 bit_90_16 bitb_90_16 word90_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_16 q_91_16 qb_91_16 bit_91_16 bitb_91_16 word91_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_16 q_92_16 qb_92_16 bit_92_16 bitb_92_16 word92_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_16 q_93_16 qb_93_16 bit_93_16 bitb_93_16 word93_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_16 q_94_16 qb_94_16 bit_94_16 bitb_94_16 word94_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_16 q_95_16 qb_95_16 bit_95_16 bitb_95_16 word95_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_16 q_96_16 qb_96_16 bit_96_16 bitb_96_16 word96_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_16 q_97_16 qb_97_16 bit_97_16 bitb_97_16 word97_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_16 q_98_16 qb_98_16 bit_98_16 bitb_98_16 word98_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_16 q_99_16 qb_99_16 bit_99_16 bitb_99_16 word99_16 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_17 q_0_17 qb_0_17 bit_0_17 bitb_0_17 word0_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_17 q_1_17 qb_1_17 bit_1_17 bitb_1_17 word1_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_17 q_2_17 qb_2_17 bit_2_17 bitb_2_17 word2_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_17 q_3_17 qb_3_17 bit_3_17 bitb_3_17 word3_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_17 q_4_17 qb_4_17 bit_4_17 bitb_4_17 word4_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_17 q_5_17 qb_5_17 bit_5_17 bitb_5_17 word5_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_17 q_6_17 qb_6_17 bit_6_17 bitb_6_17 word6_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_17 q_7_17 qb_7_17 bit_7_17 bitb_7_17 word7_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_17 q_8_17 qb_8_17 bit_8_17 bitb_8_17 word8_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_17 q_9_17 qb_9_17 bit_9_17 bitb_9_17 word9_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_17 q_10_17 qb_10_17 bit_10_17 bitb_10_17 word10_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_17 q_11_17 qb_11_17 bit_11_17 bitb_11_17 word11_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_17 q_12_17 qb_12_17 bit_12_17 bitb_12_17 word12_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_17 q_13_17 qb_13_17 bit_13_17 bitb_13_17 word13_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_17 q_14_17 qb_14_17 bit_14_17 bitb_14_17 word14_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_17 q_15_17 qb_15_17 bit_15_17 bitb_15_17 word15_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_17 q_16_17 qb_16_17 bit_16_17 bitb_16_17 word16_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_17 q_17_17 qb_17_17 bit_17_17 bitb_17_17 word17_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_17 q_18_17 qb_18_17 bit_18_17 bitb_18_17 word18_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_17 q_19_17 qb_19_17 bit_19_17 bitb_19_17 word19_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_17 q_20_17 qb_20_17 bit_20_17 bitb_20_17 word20_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_17 q_21_17 qb_21_17 bit_21_17 bitb_21_17 word21_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_17 q_22_17 qb_22_17 bit_22_17 bitb_22_17 word22_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_17 q_23_17 qb_23_17 bit_23_17 bitb_23_17 word23_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_17 q_24_17 qb_24_17 bit_24_17 bitb_24_17 word24_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_17 q_25_17 qb_25_17 bit_25_17 bitb_25_17 word25_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_17 q_26_17 qb_26_17 bit_26_17 bitb_26_17 word26_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_17 q_27_17 qb_27_17 bit_27_17 bitb_27_17 word27_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_17 q_28_17 qb_28_17 bit_28_17 bitb_28_17 word28_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_17 q_29_17 qb_29_17 bit_29_17 bitb_29_17 word29_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_17 q_30_17 qb_30_17 bit_30_17 bitb_30_17 word30_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_17 q_31_17 qb_31_17 bit_31_17 bitb_31_17 word31_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_17 q_32_17 qb_32_17 bit_32_17 bitb_32_17 word32_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_17 q_33_17 qb_33_17 bit_33_17 bitb_33_17 word33_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_17 q_34_17 qb_34_17 bit_34_17 bitb_34_17 word34_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_17 q_35_17 qb_35_17 bit_35_17 bitb_35_17 word35_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_17 q_36_17 qb_36_17 bit_36_17 bitb_36_17 word36_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_17 q_37_17 qb_37_17 bit_37_17 bitb_37_17 word37_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_17 q_38_17 qb_38_17 bit_38_17 bitb_38_17 word38_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_17 q_39_17 qb_39_17 bit_39_17 bitb_39_17 word39_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_17 q_40_17 qb_40_17 bit_40_17 bitb_40_17 word40_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_17 q_41_17 qb_41_17 bit_41_17 bitb_41_17 word41_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_17 q_42_17 qb_42_17 bit_42_17 bitb_42_17 word42_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_17 q_43_17 qb_43_17 bit_43_17 bitb_43_17 word43_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_17 q_44_17 qb_44_17 bit_44_17 bitb_44_17 word44_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_17 q_45_17 qb_45_17 bit_45_17 bitb_45_17 word45_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_17 q_46_17 qb_46_17 bit_46_17 bitb_46_17 word46_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_17 q_47_17 qb_47_17 bit_47_17 bitb_47_17 word47_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_17 q_48_17 qb_48_17 bit_48_17 bitb_48_17 word48_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_17 q_49_17 qb_49_17 bit_49_17 bitb_49_17 word49_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_17 q_50_17 qb_50_17 bit_50_17 bitb_50_17 word50_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_17 q_51_17 qb_51_17 bit_51_17 bitb_51_17 word51_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_17 q_52_17 qb_52_17 bit_52_17 bitb_52_17 word52_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_17 q_53_17 qb_53_17 bit_53_17 bitb_53_17 word53_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_17 q_54_17 qb_54_17 bit_54_17 bitb_54_17 word54_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_17 q_55_17 qb_55_17 bit_55_17 bitb_55_17 word55_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_17 q_56_17 qb_56_17 bit_56_17 bitb_56_17 word56_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_17 q_57_17 qb_57_17 bit_57_17 bitb_57_17 word57_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_17 q_58_17 qb_58_17 bit_58_17 bitb_58_17 word58_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_17 q_59_17 qb_59_17 bit_59_17 bitb_59_17 word59_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_17 q_60_17 qb_60_17 bit_60_17 bitb_60_17 word60_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_17 q_61_17 qb_61_17 bit_61_17 bitb_61_17 word61_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_17 q_62_17 qb_62_17 bit_62_17 bitb_62_17 word62_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_17 q_63_17 qb_63_17 bit_63_17 bitb_63_17 word63_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_17 q_64_17 qb_64_17 bit_64_17 bitb_64_17 word64_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_17 q_65_17 qb_65_17 bit_65_17 bitb_65_17 word65_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_17 q_66_17 qb_66_17 bit_66_17 bitb_66_17 word66_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_17 q_67_17 qb_67_17 bit_67_17 bitb_67_17 word67_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_17 q_68_17 qb_68_17 bit_68_17 bitb_68_17 word68_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_17 q_69_17 qb_69_17 bit_69_17 bitb_69_17 word69_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_17 q_70_17 qb_70_17 bit_70_17 bitb_70_17 word70_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_17 q_71_17 qb_71_17 bit_71_17 bitb_71_17 word71_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_17 q_72_17 qb_72_17 bit_72_17 bitb_72_17 word72_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_17 q_73_17 qb_73_17 bit_73_17 bitb_73_17 word73_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_17 q_74_17 qb_74_17 bit_74_17 bitb_74_17 word74_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_17 q_75_17 qb_75_17 bit_75_17 bitb_75_17 word75_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_17 q_76_17 qb_76_17 bit_76_17 bitb_76_17 word76_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_17 q_77_17 qb_77_17 bit_77_17 bitb_77_17 word77_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_17 q_78_17 qb_78_17 bit_78_17 bitb_78_17 word78_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_17 q_79_17 qb_79_17 bit_79_17 bitb_79_17 word79_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_17 q_80_17 qb_80_17 bit_80_17 bitb_80_17 word80_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_17 q_81_17 qb_81_17 bit_81_17 bitb_81_17 word81_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_17 q_82_17 qb_82_17 bit_82_17 bitb_82_17 word82_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_17 q_83_17 qb_83_17 bit_83_17 bitb_83_17 word83_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_17 q_84_17 qb_84_17 bit_84_17 bitb_84_17 word84_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_17 q_85_17 qb_85_17 bit_85_17 bitb_85_17 word85_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_17 q_86_17 qb_86_17 bit_86_17 bitb_86_17 word86_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_17 q_87_17 qb_87_17 bit_87_17 bitb_87_17 word87_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_17 q_88_17 qb_88_17 bit_88_17 bitb_88_17 word88_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_17 q_89_17 qb_89_17 bit_89_17 bitb_89_17 word89_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_17 q_90_17 qb_90_17 bit_90_17 bitb_90_17 word90_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_17 q_91_17 qb_91_17 bit_91_17 bitb_91_17 word91_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_17 q_92_17 qb_92_17 bit_92_17 bitb_92_17 word92_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_17 q_93_17 qb_93_17 bit_93_17 bitb_93_17 word93_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_17 q_94_17 qb_94_17 bit_94_17 bitb_94_17 word94_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_17 q_95_17 qb_95_17 bit_95_17 bitb_95_17 word95_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_17 q_96_17 qb_96_17 bit_96_17 bitb_96_17 word96_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_17 q_97_17 qb_97_17 bit_97_17 bitb_97_17 word97_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_17 q_98_17 qb_98_17 bit_98_17 bitb_98_17 word98_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_17 q_99_17 qb_99_17 bit_99_17 bitb_99_17 word99_17 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_18 q_0_18 qb_0_18 bit_0_18 bitb_0_18 word0_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_18 q_1_18 qb_1_18 bit_1_18 bitb_1_18 word1_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_18 q_2_18 qb_2_18 bit_2_18 bitb_2_18 word2_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_18 q_3_18 qb_3_18 bit_3_18 bitb_3_18 word3_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_18 q_4_18 qb_4_18 bit_4_18 bitb_4_18 word4_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_18 q_5_18 qb_5_18 bit_5_18 bitb_5_18 word5_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_18 q_6_18 qb_6_18 bit_6_18 bitb_6_18 word6_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_18 q_7_18 qb_7_18 bit_7_18 bitb_7_18 word7_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_18 q_8_18 qb_8_18 bit_8_18 bitb_8_18 word8_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_18 q_9_18 qb_9_18 bit_9_18 bitb_9_18 word9_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_18 q_10_18 qb_10_18 bit_10_18 bitb_10_18 word10_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_18 q_11_18 qb_11_18 bit_11_18 bitb_11_18 word11_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_18 q_12_18 qb_12_18 bit_12_18 bitb_12_18 word12_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_18 q_13_18 qb_13_18 bit_13_18 bitb_13_18 word13_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_18 q_14_18 qb_14_18 bit_14_18 bitb_14_18 word14_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_18 q_15_18 qb_15_18 bit_15_18 bitb_15_18 word15_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_18 q_16_18 qb_16_18 bit_16_18 bitb_16_18 word16_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_18 q_17_18 qb_17_18 bit_17_18 bitb_17_18 word17_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_18 q_18_18 qb_18_18 bit_18_18 bitb_18_18 word18_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_18 q_19_18 qb_19_18 bit_19_18 bitb_19_18 word19_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_18 q_20_18 qb_20_18 bit_20_18 bitb_20_18 word20_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_18 q_21_18 qb_21_18 bit_21_18 bitb_21_18 word21_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_18 q_22_18 qb_22_18 bit_22_18 bitb_22_18 word22_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_18 q_23_18 qb_23_18 bit_23_18 bitb_23_18 word23_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_18 q_24_18 qb_24_18 bit_24_18 bitb_24_18 word24_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_18 q_25_18 qb_25_18 bit_25_18 bitb_25_18 word25_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_18 q_26_18 qb_26_18 bit_26_18 bitb_26_18 word26_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_18 q_27_18 qb_27_18 bit_27_18 bitb_27_18 word27_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_18 q_28_18 qb_28_18 bit_28_18 bitb_28_18 word28_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_18 q_29_18 qb_29_18 bit_29_18 bitb_29_18 word29_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_18 q_30_18 qb_30_18 bit_30_18 bitb_30_18 word30_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_18 q_31_18 qb_31_18 bit_31_18 bitb_31_18 word31_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_18 q_32_18 qb_32_18 bit_32_18 bitb_32_18 word32_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_18 q_33_18 qb_33_18 bit_33_18 bitb_33_18 word33_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_18 q_34_18 qb_34_18 bit_34_18 bitb_34_18 word34_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_18 q_35_18 qb_35_18 bit_35_18 bitb_35_18 word35_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_18 q_36_18 qb_36_18 bit_36_18 bitb_36_18 word36_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_18 q_37_18 qb_37_18 bit_37_18 bitb_37_18 word37_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_18 q_38_18 qb_38_18 bit_38_18 bitb_38_18 word38_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_18 q_39_18 qb_39_18 bit_39_18 bitb_39_18 word39_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_18 q_40_18 qb_40_18 bit_40_18 bitb_40_18 word40_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_18 q_41_18 qb_41_18 bit_41_18 bitb_41_18 word41_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_18 q_42_18 qb_42_18 bit_42_18 bitb_42_18 word42_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_18 q_43_18 qb_43_18 bit_43_18 bitb_43_18 word43_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_18 q_44_18 qb_44_18 bit_44_18 bitb_44_18 word44_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_18 q_45_18 qb_45_18 bit_45_18 bitb_45_18 word45_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_18 q_46_18 qb_46_18 bit_46_18 bitb_46_18 word46_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_18 q_47_18 qb_47_18 bit_47_18 bitb_47_18 word47_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_18 q_48_18 qb_48_18 bit_48_18 bitb_48_18 word48_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_18 q_49_18 qb_49_18 bit_49_18 bitb_49_18 word49_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_18 q_50_18 qb_50_18 bit_50_18 bitb_50_18 word50_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_18 q_51_18 qb_51_18 bit_51_18 bitb_51_18 word51_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_18 q_52_18 qb_52_18 bit_52_18 bitb_52_18 word52_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_18 q_53_18 qb_53_18 bit_53_18 bitb_53_18 word53_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_18 q_54_18 qb_54_18 bit_54_18 bitb_54_18 word54_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_18 q_55_18 qb_55_18 bit_55_18 bitb_55_18 word55_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_18 q_56_18 qb_56_18 bit_56_18 bitb_56_18 word56_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_18 q_57_18 qb_57_18 bit_57_18 bitb_57_18 word57_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_18 q_58_18 qb_58_18 bit_58_18 bitb_58_18 word58_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_18 q_59_18 qb_59_18 bit_59_18 bitb_59_18 word59_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_18 q_60_18 qb_60_18 bit_60_18 bitb_60_18 word60_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_18 q_61_18 qb_61_18 bit_61_18 bitb_61_18 word61_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_18 q_62_18 qb_62_18 bit_62_18 bitb_62_18 word62_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_18 q_63_18 qb_63_18 bit_63_18 bitb_63_18 word63_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_18 q_64_18 qb_64_18 bit_64_18 bitb_64_18 word64_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_18 q_65_18 qb_65_18 bit_65_18 bitb_65_18 word65_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_18 q_66_18 qb_66_18 bit_66_18 bitb_66_18 word66_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_18 q_67_18 qb_67_18 bit_67_18 bitb_67_18 word67_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_18 q_68_18 qb_68_18 bit_68_18 bitb_68_18 word68_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_18 q_69_18 qb_69_18 bit_69_18 bitb_69_18 word69_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_18 q_70_18 qb_70_18 bit_70_18 bitb_70_18 word70_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_18 q_71_18 qb_71_18 bit_71_18 bitb_71_18 word71_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_18 q_72_18 qb_72_18 bit_72_18 bitb_72_18 word72_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_18 q_73_18 qb_73_18 bit_73_18 bitb_73_18 word73_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_18 q_74_18 qb_74_18 bit_74_18 bitb_74_18 word74_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_18 q_75_18 qb_75_18 bit_75_18 bitb_75_18 word75_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_18 q_76_18 qb_76_18 bit_76_18 bitb_76_18 word76_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_18 q_77_18 qb_77_18 bit_77_18 bitb_77_18 word77_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_18 q_78_18 qb_78_18 bit_78_18 bitb_78_18 word78_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_18 q_79_18 qb_79_18 bit_79_18 bitb_79_18 word79_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_18 q_80_18 qb_80_18 bit_80_18 bitb_80_18 word80_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_18 q_81_18 qb_81_18 bit_81_18 bitb_81_18 word81_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_18 q_82_18 qb_82_18 bit_82_18 bitb_82_18 word82_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_18 q_83_18 qb_83_18 bit_83_18 bitb_83_18 word83_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_18 q_84_18 qb_84_18 bit_84_18 bitb_84_18 word84_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_18 q_85_18 qb_85_18 bit_85_18 bitb_85_18 word85_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_18 q_86_18 qb_86_18 bit_86_18 bitb_86_18 word86_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_18 q_87_18 qb_87_18 bit_87_18 bitb_87_18 word87_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_18 q_88_18 qb_88_18 bit_88_18 bitb_88_18 word88_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_18 q_89_18 qb_89_18 bit_89_18 bitb_89_18 word89_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_18 q_90_18 qb_90_18 bit_90_18 bitb_90_18 word90_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_18 q_91_18 qb_91_18 bit_91_18 bitb_91_18 word91_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_18 q_92_18 qb_92_18 bit_92_18 bitb_92_18 word92_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_18 q_93_18 qb_93_18 bit_93_18 bitb_93_18 word93_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_18 q_94_18 qb_94_18 bit_94_18 bitb_94_18 word94_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_18 q_95_18 qb_95_18 bit_95_18 bitb_95_18 word95_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_18 q_96_18 qb_96_18 bit_96_18 bitb_96_18 word96_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_18 q_97_18 qb_97_18 bit_97_18 bitb_97_18 word97_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_18 q_98_18 qb_98_18 bit_98_18 bitb_98_18 word98_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_18 q_99_18 qb_99_18 bit_99_18 bitb_99_18 word99_18 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_19 q_0_19 qb_0_19 bit_0_19 bitb_0_19 word0_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_19 q_1_19 qb_1_19 bit_1_19 bitb_1_19 word1_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_19 q_2_19 qb_2_19 bit_2_19 bitb_2_19 word2_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_19 q_3_19 qb_3_19 bit_3_19 bitb_3_19 word3_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_19 q_4_19 qb_4_19 bit_4_19 bitb_4_19 word4_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_19 q_5_19 qb_5_19 bit_5_19 bitb_5_19 word5_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_19 q_6_19 qb_6_19 bit_6_19 bitb_6_19 word6_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_19 q_7_19 qb_7_19 bit_7_19 bitb_7_19 word7_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_19 q_8_19 qb_8_19 bit_8_19 bitb_8_19 word8_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_19 q_9_19 qb_9_19 bit_9_19 bitb_9_19 word9_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_19 q_10_19 qb_10_19 bit_10_19 bitb_10_19 word10_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_19 q_11_19 qb_11_19 bit_11_19 bitb_11_19 word11_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_19 q_12_19 qb_12_19 bit_12_19 bitb_12_19 word12_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_19 q_13_19 qb_13_19 bit_13_19 bitb_13_19 word13_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_19 q_14_19 qb_14_19 bit_14_19 bitb_14_19 word14_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_19 q_15_19 qb_15_19 bit_15_19 bitb_15_19 word15_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_19 q_16_19 qb_16_19 bit_16_19 bitb_16_19 word16_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_19 q_17_19 qb_17_19 bit_17_19 bitb_17_19 word17_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_19 q_18_19 qb_18_19 bit_18_19 bitb_18_19 word18_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_19 q_19_19 qb_19_19 bit_19_19 bitb_19_19 word19_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_19 q_20_19 qb_20_19 bit_20_19 bitb_20_19 word20_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_19 q_21_19 qb_21_19 bit_21_19 bitb_21_19 word21_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_19 q_22_19 qb_22_19 bit_22_19 bitb_22_19 word22_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_19 q_23_19 qb_23_19 bit_23_19 bitb_23_19 word23_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_19 q_24_19 qb_24_19 bit_24_19 bitb_24_19 word24_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_19 q_25_19 qb_25_19 bit_25_19 bitb_25_19 word25_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_19 q_26_19 qb_26_19 bit_26_19 bitb_26_19 word26_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_19 q_27_19 qb_27_19 bit_27_19 bitb_27_19 word27_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_19 q_28_19 qb_28_19 bit_28_19 bitb_28_19 word28_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_19 q_29_19 qb_29_19 bit_29_19 bitb_29_19 word29_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_19 q_30_19 qb_30_19 bit_30_19 bitb_30_19 word30_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_19 q_31_19 qb_31_19 bit_31_19 bitb_31_19 word31_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_19 q_32_19 qb_32_19 bit_32_19 bitb_32_19 word32_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_19 q_33_19 qb_33_19 bit_33_19 bitb_33_19 word33_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_19 q_34_19 qb_34_19 bit_34_19 bitb_34_19 word34_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_19 q_35_19 qb_35_19 bit_35_19 bitb_35_19 word35_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_19 q_36_19 qb_36_19 bit_36_19 bitb_36_19 word36_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_19 q_37_19 qb_37_19 bit_37_19 bitb_37_19 word37_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_19 q_38_19 qb_38_19 bit_38_19 bitb_38_19 word38_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_19 q_39_19 qb_39_19 bit_39_19 bitb_39_19 word39_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_19 q_40_19 qb_40_19 bit_40_19 bitb_40_19 word40_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_19 q_41_19 qb_41_19 bit_41_19 bitb_41_19 word41_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_19 q_42_19 qb_42_19 bit_42_19 bitb_42_19 word42_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_19 q_43_19 qb_43_19 bit_43_19 bitb_43_19 word43_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_19 q_44_19 qb_44_19 bit_44_19 bitb_44_19 word44_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_19 q_45_19 qb_45_19 bit_45_19 bitb_45_19 word45_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_19 q_46_19 qb_46_19 bit_46_19 bitb_46_19 word46_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_19 q_47_19 qb_47_19 bit_47_19 bitb_47_19 word47_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_19 q_48_19 qb_48_19 bit_48_19 bitb_48_19 word48_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_19 q_49_19 qb_49_19 bit_49_19 bitb_49_19 word49_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_19 q_50_19 qb_50_19 bit_50_19 bitb_50_19 word50_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_19 q_51_19 qb_51_19 bit_51_19 bitb_51_19 word51_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_19 q_52_19 qb_52_19 bit_52_19 bitb_52_19 word52_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_19 q_53_19 qb_53_19 bit_53_19 bitb_53_19 word53_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_19 q_54_19 qb_54_19 bit_54_19 bitb_54_19 word54_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_19 q_55_19 qb_55_19 bit_55_19 bitb_55_19 word55_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_19 q_56_19 qb_56_19 bit_56_19 bitb_56_19 word56_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_19 q_57_19 qb_57_19 bit_57_19 bitb_57_19 word57_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_19 q_58_19 qb_58_19 bit_58_19 bitb_58_19 word58_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_19 q_59_19 qb_59_19 bit_59_19 bitb_59_19 word59_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_19 q_60_19 qb_60_19 bit_60_19 bitb_60_19 word60_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_19 q_61_19 qb_61_19 bit_61_19 bitb_61_19 word61_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_19 q_62_19 qb_62_19 bit_62_19 bitb_62_19 word62_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_19 q_63_19 qb_63_19 bit_63_19 bitb_63_19 word63_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_19 q_64_19 qb_64_19 bit_64_19 bitb_64_19 word64_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_19 q_65_19 qb_65_19 bit_65_19 bitb_65_19 word65_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_19 q_66_19 qb_66_19 bit_66_19 bitb_66_19 word66_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_19 q_67_19 qb_67_19 bit_67_19 bitb_67_19 word67_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_19 q_68_19 qb_68_19 bit_68_19 bitb_68_19 word68_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_19 q_69_19 qb_69_19 bit_69_19 bitb_69_19 word69_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_19 q_70_19 qb_70_19 bit_70_19 bitb_70_19 word70_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_19 q_71_19 qb_71_19 bit_71_19 bitb_71_19 word71_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_19 q_72_19 qb_72_19 bit_72_19 bitb_72_19 word72_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_19 q_73_19 qb_73_19 bit_73_19 bitb_73_19 word73_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_19 q_74_19 qb_74_19 bit_74_19 bitb_74_19 word74_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_19 q_75_19 qb_75_19 bit_75_19 bitb_75_19 word75_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_19 q_76_19 qb_76_19 bit_76_19 bitb_76_19 word76_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_19 q_77_19 qb_77_19 bit_77_19 bitb_77_19 word77_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_19 q_78_19 qb_78_19 bit_78_19 bitb_78_19 word78_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_19 q_79_19 qb_79_19 bit_79_19 bitb_79_19 word79_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_19 q_80_19 qb_80_19 bit_80_19 bitb_80_19 word80_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_19 q_81_19 qb_81_19 bit_81_19 bitb_81_19 word81_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_19 q_82_19 qb_82_19 bit_82_19 bitb_82_19 word82_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_19 q_83_19 qb_83_19 bit_83_19 bitb_83_19 word83_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_19 q_84_19 qb_84_19 bit_84_19 bitb_84_19 word84_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_19 q_85_19 qb_85_19 bit_85_19 bitb_85_19 word85_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_19 q_86_19 qb_86_19 bit_86_19 bitb_86_19 word86_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_19 q_87_19 qb_87_19 bit_87_19 bitb_87_19 word87_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_19 q_88_19 qb_88_19 bit_88_19 bitb_88_19 word88_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_19 q_89_19 qb_89_19 bit_89_19 bitb_89_19 word89_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_19 q_90_19 qb_90_19 bit_90_19 bitb_90_19 word90_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_19 q_91_19 qb_91_19 bit_91_19 bitb_91_19 word91_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_19 q_92_19 qb_92_19 bit_92_19 bitb_92_19 word92_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_19 q_93_19 qb_93_19 bit_93_19 bitb_93_19 word93_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_19 q_94_19 qb_94_19 bit_94_19 bitb_94_19 word94_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_19 q_95_19 qb_95_19 bit_95_19 bitb_95_19 word95_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_19 q_96_19 qb_96_19 bit_96_19 bitb_96_19 word96_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_19 q_97_19 qb_97_19 bit_97_19 bitb_97_19 word97_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_19 q_98_19 qb_98_19 bit_98_19 bitb_98_19 word98_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_19 q_99_19 qb_99_19 bit_99_19 bitb_99_19 word99_19 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_20 q_0_20 qb_0_20 bit_0_20 bitb_0_20 word0_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_20 q_1_20 qb_1_20 bit_1_20 bitb_1_20 word1_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_20 q_2_20 qb_2_20 bit_2_20 bitb_2_20 word2_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_20 q_3_20 qb_3_20 bit_3_20 bitb_3_20 word3_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_20 q_4_20 qb_4_20 bit_4_20 bitb_4_20 word4_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_20 q_5_20 qb_5_20 bit_5_20 bitb_5_20 word5_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_20 q_6_20 qb_6_20 bit_6_20 bitb_6_20 word6_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_20 q_7_20 qb_7_20 bit_7_20 bitb_7_20 word7_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_20 q_8_20 qb_8_20 bit_8_20 bitb_8_20 word8_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_20 q_9_20 qb_9_20 bit_9_20 bitb_9_20 word9_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_20 q_10_20 qb_10_20 bit_10_20 bitb_10_20 word10_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_20 q_11_20 qb_11_20 bit_11_20 bitb_11_20 word11_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_20 q_12_20 qb_12_20 bit_12_20 bitb_12_20 word12_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_20 q_13_20 qb_13_20 bit_13_20 bitb_13_20 word13_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_20 q_14_20 qb_14_20 bit_14_20 bitb_14_20 word14_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_20 q_15_20 qb_15_20 bit_15_20 bitb_15_20 word15_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_20 q_16_20 qb_16_20 bit_16_20 bitb_16_20 word16_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_20 q_17_20 qb_17_20 bit_17_20 bitb_17_20 word17_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_20 q_18_20 qb_18_20 bit_18_20 bitb_18_20 word18_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_20 q_19_20 qb_19_20 bit_19_20 bitb_19_20 word19_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_20 q_20_20 qb_20_20 bit_20_20 bitb_20_20 word20_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_20 q_21_20 qb_21_20 bit_21_20 bitb_21_20 word21_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_20 q_22_20 qb_22_20 bit_22_20 bitb_22_20 word22_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_20 q_23_20 qb_23_20 bit_23_20 bitb_23_20 word23_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_20 q_24_20 qb_24_20 bit_24_20 bitb_24_20 word24_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_20 q_25_20 qb_25_20 bit_25_20 bitb_25_20 word25_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_20 q_26_20 qb_26_20 bit_26_20 bitb_26_20 word26_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_20 q_27_20 qb_27_20 bit_27_20 bitb_27_20 word27_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_20 q_28_20 qb_28_20 bit_28_20 bitb_28_20 word28_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_20 q_29_20 qb_29_20 bit_29_20 bitb_29_20 word29_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_20 q_30_20 qb_30_20 bit_30_20 bitb_30_20 word30_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_20 q_31_20 qb_31_20 bit_31_20 bitb_31_20 word31_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_20 q_32_20 qb_32_20 bit_32_20 bitb_32_20 word32_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_20 q_33_20 qb_33_20 bit_33_20 bitb_33_20 word33_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_20 q_34_20 qb_34_20 bit_34_20 bitb_34_20 word34_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_20 q_35_20 qb_35_20 bit_35_20 bitb_35_20 word35_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_20 q_36_20 qb_36_20 bit_36_20 bitb_36_20 word36_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_20 q_37_20 qb_37_20 bit_37_20 bitb_37_20 word37_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_20 q_38_20 qb_38_20 bit_38_20 bitb_38_20 word38_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_20 q_39_20 qb_39_20 bit_39_20 bitb_39_20 word39_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_20 q_40_20 qb_40_20 bit_40_20 bitb_40_20 word40_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_20 q_41_20 qb_41_20 bit_41_20 bitb_41_20 word41_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_20 q_42_20 qb_42_20 bit_42_20 bitb_42_20 word42_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_20 q_43_20 qb_43_20 bit_43_20 bitb_43_20 word43_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_20 q_44_20 qb_44_20 bit_44_20 bitb_44_20 word44_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_20 q_45_20 qb_45_20 bit_45_20 bitb_45_20 word45_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_20 q_46_20 qb_46_20 bit_46_20 bitb_46_20 word46_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_20 q_47_20 qb_47_20 bit_47_20 bitb_47_20 word47_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_20 q_48_20 qb_48_20 bit_48_20 bitb_48_20 word48_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_20 q_49_20 qb_49_20 bit_49_20 bitb_49_20 word49_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_20 q_50_20 qb_50_20 bit_50_20 bitb_50_20 word50_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_20 q_51_20 qb_51_20 bit_51_20 bitb_51_20 word51_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_20 q_52_20 qb_52_20 bit_52_20 bitb_52_20 word52_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_20 q_53_20 qb_53_20 bit_53_20 bitb_53_20 word53_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_20 q_54_20 qb_54_20 bit_54_20 bitb_54_20 word54_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_20 q_55_20 qb_55_20 bit_55_20 bitb_55_20 word55_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_20 q_56_20 qb_56_20 bit_56_20 bitb_56_20 word56_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_20 q_57_20 qb_57_20 bit_57_20 bitb_57_20 word57_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_20 q_58_20 qb_58_20 bit_58_20 bitb_58_20 word58_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_20 q_59_20 qb_59_20 bit_59_20 bitb_59_20 word59_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_20 q_60_20 qb_60_20 bit_60_20 bitb_60_20 word60_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_20 q_61_20 qb_61_20 bit_61_20 bitb_61_20 word61_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_20 q_62_20 qb_62_20 bit_62_20 bitb_62_20 word62_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_20 q_63_20 qb_63_20 bit_63_20 bitb_63_20 word63_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_20 q_64_20 qb_64_20 bit_64_20 bitb_64_20 word64_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_20 q_65_20 qb_65_20 bit_65_20 bitb_65_20 word65_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_20 q_66_20 qb_66_20 bit_66_20 bitb_66_20 word66_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_20 q_67_20 qb_67_20 bit_67_20 bitb_67_20 word67_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_20 q_68_20 qb_68_20 bit_68_20 bitb_68_20 word68_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_20 q_69_20 qb_69_20 bit_69_20 bitb_69_20 word69_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_20 q_70_20 qb_70_20 bit_70_20 bitb_70_20 word70_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_20 q_71_20 qb_71_20 bit_71_20 bitb_71_20 word71_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_20 q_72_20 qb_72_20 bit_72_20 bitb_72_20 word72_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_20 q_73_20 qb_73_20 bit_73_20 bitb_73_20 word73_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_20 q_74_20 qb_74_20 bit_74_20 bitb_74_20 word74_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_20 q_75_20 qb_75_20 bit_75_20 bitb_75_20 word75_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_20 q_76_20 qb_76_20 bit_76_20 bitb_76_20 word76_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_20 q_77_20 qb_77_20 bit_77_20 bitb_77_20 word77_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_20 q_78_20 qb_78_20 bit_78_20 bitb_78_20 word78_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_20 q_79_20 qb_79_20 bit_79_20 bitb_79_20 word79_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_20 q_80_20 qb_80_20 bit_80_20 bitb_80_20 word80_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_20 q_81_20 qb_81_20 bit_81_20 bitb_81_20 word81_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_20 q_82_20 qb_82_20 bit_82_20 bitb_82_20 word82_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_20 q_83_20 qb_83_20 bit_83_20 bitb_83_20 word83_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_20 q_84_20 qb_84_20 bit_84_20 bitb_84_20 word84_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_20 q_85_20 qb_85_20 bit_85_20 bitb_85_20 word85_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_20 q_86_20 qb_86_20 bit_86_20 bitb_86_20 word86_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_20 q_87_20 qb_87_20 bit_87_20 bitb_87_20 word87_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_20 q_88_20 qb_88_20 bit_88_20 bitb_88_20 word88_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_20 q_89_20 qb_89_20 bit_89_20 bitb_89_20 word89_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_20 q_90_20 qb_90_20 bit_90_20 bitb_90_20 word90_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_20 q_91_20 qb_91_20 bit_91_20 bitb_91_20 word91_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_20 q_92_20 qb_92_20 bit_92_20 bitb_92_20 word92_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_20 q_93_20 qb_93_20 bit_93_20 bitb_93_20 word93_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_20 q_94_20 qb_94_20 bit_94_20 bitb_94_20 word94_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_20 q_95_20 qb_95_20 bit_95_20 bitb_95_20 word95_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_20 q_96_20 qb_96_20 bit_96_20 bitb_96_20 word96_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_20 q_97_20 qb_97_20 bit_97_20 bitb_97_20 word97_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_20 q_98_20 qb_98_20 bit_98_20 bitb_98_20 word98_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_20 q_99_20 qb_99_20 bit_99_20 bitb_99_20 word99_20 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_21 q_0_21 qb_0_21 bit_0_21 bitb_0_21 word0_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_21 q_1_21 qb_1_21 bit_1_21 bitb_1_21 word1_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_21 q_2_21 qb_2_21 bit_2_21 bitb_2_21 word2_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_21 q_3_21 qb_3_21 bit_3_21 bitb_3_21 word3_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_21 q_4_21 qb_4_21 bit_4_21 bitb_4_21 word4_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_21 q_5_21 qb_5_21 bit_5_21 bitb_5_21 word5_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_21 q_6_21 qb_6_21 bit_6_21 bitb_6_21 word6_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_21 q_7_21 qb_7_21 bit_7_21 bitb_7_21 word7_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_21 q_8_21 qb_8_21 bit_8_21 bitb_8_21 word8_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_21 q_9_21 qb_9_21 bit_9_21 bitb_9_21 word9_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_21 q_10_21 qb_10_21 bit_10_21 bitb_10_21 word10_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_21 q_11_21 qb_11_21 bit_11_21 bitb_11_21 word11_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_21 q_12_21 qb_12_21 bit_12_21 bitb_12_21 word12_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_21 q_13_21 qb_13_21 bit_13_21 bitb_13_21 word13_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_21 q_14_21 qb_14_21 bit_14_21 bitb_14_21 word14_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_21 q_15_21 qb_15_21 bit_15_21 bitb_15_21 word15_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_21 q_16_21 qb_16_21 bit_16_21 bitb_16_21 word16_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_21 q_17_21 qb_17_21 bit_17_21 bitb_17_21 word17_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_21 q_18_21 qb_18_21 bit_18_21 bitb_18_21 word18_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_21 q_19_21 qb_19_21 bit_19_21 bitb_19_21 word19_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_21 q_20_21 qb_20_21 bit_20_21 bitb_20_21 word20_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_21 q_21_21 qb_21_21 bit_21_21 bitb_21_21 word21_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_21 q_22_21 qb_22_21 bit_22_21 bitb_22_21 word22_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_21 q_23_21 qb_23_21 bit_23_21 bitb_23_21 word23_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_21 q_24_21 qb_24_21 bit_24_21 bitb_24_21 word24_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_21 q_25_21 qb_25_21 bit_25_21 bitb_25_21 word25_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_21 q_26_21 qb_26_21 bit_26_21 bitb_26_21 word26_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_21 q_27_21 qb_27_21 bit_27_21 bitb_27_21 word27_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_21 q_28_21 qb_28_21 bit_28_21 bitb_28_21 word28_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_21 q_29_21 qb_29_21 bit_29_21 bitb_29_21 word29_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_21 q_30_21 qb_30_21 bit_30_21 bitb_30_21 word30_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_21 q_31_21 qb_31_21 bit_31_21 bitb_31_21 word31_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_21 q_32_21 qb_32_21 bit_32_21 bitb_32_21 word32_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_21 q_33_21 qb_33_21 bit_33_21 bitb_33_21 word33_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_21 q_34_21 qb_34_21 bit_34_21 bitb_34_21 word34_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_21 q_35_21 qb_35_21 bit_35_21 bitb_35_21 word35_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_21 q_36_21 qb_36_21 bit_36_21 bitb_36_21 word36_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_21 q_37_21 qb_37_21 bit_37_21 bitb_37_21 word37_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_21 q_38_21 qb_38_21 bit_38_21 bitb_38_21 word38_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_21 q_39_21 qb_39_21 bit_39_21 bitb_39_21 word39_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_21 q_40_21 qb_40_21 bit_40_21 bitb_40_21 word40_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_21 q_41_21 qb_41_21 bit_41_21 bitb_41_21 word41_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_21 q_42_21 qb_42_21 bit_42_21 bitb_42_21 word42_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_21 q_43_21 qb_43_21 bit_43_21 bitb_43_21 word43_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_21 q_44_21 qb_44_21 bit_44_21 bitb_44_21 word44_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_21 q_45_21 qb_45_21 bit_45_21 bitb_45_21 word45_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_21 q_46_21 qb_46_21 bit_46_21 bitb_46_21 word46_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_21 q_47_21 qb_47_21 bit_47_21 bitb_47_21 word47_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_21 q_48_21 qb_48_21 bit_48_21 bitb_48_21 word48_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_21 q_49_21 qb_49_21 bit_49_21 bitb_49_21 word49_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_21 q_50_21 qb_50_21 bit_50_21 bitb_50_21 word50_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_21 q_51_21 qb_51_21 bit_51_21 bitb_51_21 word51_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_21 q_52_21 qb_52_21 bit_52_21 bitb_52_21 word52_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_21 q_53_21 qb_53_21 bit_53_21 bitb_53_21 word53_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_21 q_54_21 qb_54_21 bit_54_21 bitb_54_21 word54_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_21 q_55_21 qb_55_21 bit_55_21 bitb_55_21 word55_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_21 q_56_21 qb_56_21 bit_56_21 bitb_56_21 word56_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_21 q_57_21 qb_57_21 bit_57_21 bitb_57_21 word57_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_21 q_58_21 qb_58_21 bit_58_21 bitb_58_21 word58_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_21 q_59_21 qb_59_21 bit_59_21 bitb_59_21 word59_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_21 q_60_21 qb_60_21 bit_60_21 bitb_60_21 word60_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_21 q_61_21 qb_61_21 bit_61_21 bitb_61_21 word61_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_21 q_62_21 qb_62_21 bit_62_21 bitb_62_21 word62_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_21 q_63_21 qb_63_21 bit_63_21 bitb_63_21 word63_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_21 q_64_21 qb_64_21 bit_64_21 bitb_64_21 word64_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_21 q_65_21 qb_65_21 bit_65_21 bitb_65_21 word65_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_21 q_66_21 qb_66_21 bit_66_21 bitb_66_21 word66_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_21 q_67_21 qb_67_21 bit_67_21 bitb_67_21 word67_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_21 q_68_21 qb_68_21 bit_68_21 bitb_68_21 word68_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_21 q_69_21 qb_69_21 bit_69_21 bitb_69_21 word69_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_21 q_70_21 qb_70_21 bit_70_21 bitb_70_21 word70_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_21 q_71_21 qb_71_21 bit_71_21 bitb_71_21 word71_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_21 q_72_21 qb_72_21 bit_72_21 bitb_72_21 word72_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_21 q_73_21 qb_73_21 bit_73_21 bitb_73_21 word73_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_21 q_74_21 qb_74_21 bit_74_21 bitb_74_21 word74_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_21 q_75_21 qb_75_21 bit_75_21 bitb_75_21 word75_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_21 q_76_21 qb_76_21 bit_76_21 bitb_76_21 word76_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_21 q_77_21 qb_77_21 bit_77_21 bitb_77_21 word77_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_21 q_78_21 qb_78_21 bit_78_21 bitb_78_21 word78_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_21 q_79_21 qb_79_21 bit_79_21 bitb_79_21 word79_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_21 q_80_21 qb_80_21 bit_80_21 bitb_80_21 word80_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_21 q_81_21 qb_81_21 bit_81_21 bitb_81_21 word81_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_21 q_82_21 qb_82_21 bit_82_21 bitb_82_21 word82_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_21 q_83_21 qb_83_21 bit_83_21 bitb_83_21 word83_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_21 q_84_21 qb_84_21 bit_84_21 bitb_84_21 word84_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_21 q_85_21 qb_85_21 bit_85_21 bitb_85_21 word85_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_21 q_86_21 qb_86_21 bit_86_21 bitb_86_21 word86_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_21 q_87_21 qb_87_21 bit_87_21 bitb_87_21 word87_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_21 q_88_21 qb_88_21 bit_88_21 bitb_88_21 word88_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_21 q_89_21 qb_89_21 bit_89_21 bitb_89_21 word89_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_21 q_90_21 qb_90_21 bit_90_21 bitb_90_21 word90_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_21 q_91_21 qb_91_21 bit_91_21 bitb_91_21 word91_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_21 q_92_21 qb_92_21 bit_92_21 bitb_92_21 word92_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_21 q_93_21 qb_93_21 bit_93_21 bitb_93_21 word93_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_21 q_94_21 qb_94_21 bit_94_21 bitb_94_21 word94_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_21 q_95_21 qb_95_21 bit_95_21 bitb_95_21 word95_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_21 q_96_21 qb_96_21 bit_96_21 bitb_96_21 word96_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_21 q_97_21 qb_97_21 bit_97_21 bitb_97_21 word97_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_21 q_98_21 qb_98_21 bit_98_21 bitb_98_21 word98_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_21 q_99_21 qb_99_21 bit_99_21 bitb_99_21 word99_21 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_22 q_0_22 qb_0_22 bit_0_22 bitb_0_22 word0_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_22 q_1_22 qb_1_22 bit_1_22 bitb_1_22 word1_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_22 q_2_22 qb_2_22 bit_2_22 bitb_2_22 word2_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_22 q_3_22 qb_3_22 bit_3_22 bitb_3_22 word3_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_22 q_4_22 qb_4_22 bit_4_22 bitb_4_22 word4_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_22 q_5_22 qb_5_22 bit_5_22 bitb_5_22 word5_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_22 q_6_22 qb_6_22 bit_6_22 bitb_6_22 word6_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_22 q_7_22 qb_7_22 bit_7_22 bitb_7_22 word7_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_22 q_8_22 qb_8_22 bit_8_22 bitb_8_22 word8_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_22 q_9_22 qb_9_22 bit_9_22 bitb_9_22 word9_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_22 q_10_22 qb_10_22 bit_10_22 bitb_10_22 word10_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_22 q_11_22 qb_11_22 bit_11_22 bitb_11_22 word11_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_22 q_12_22 qb_12_22 bit_12_22 bitb_12_22 word12_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_22 q_13_22 qb_13_22 bit_13_22 bitb_13_22 word13_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_22 q_14_22 qb_14_22 bit_14_22 bitb_14_22 word14_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_22 q_15_22 qb_15_22 bit_15_22 bitb_15_22 word15_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_22 q_16_22 qb_16_22 bit_16_22 bitb_16_22 word16_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_22 q_17_22 qb_17_22 bit_17_22 bitb_17_22 word17_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_22 q_18_22 qb_18_22 bit_18_22 bitb_18_22 word18_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_22 q_19_22 qb_19_22 bit_19_22 bitb_19_22 word19_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_22 q_20_22 qb_20_22 bit_20_22 bitb_20_22 word20_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_22 q_21_22 qb_21_22 bit_21_22 bitb_21_22 word21_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_22 q_22_22 qb_22_22 bit_22_22 bitb_22_22 word22_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_22 q_23_22 qb_23_22 bit_23_22 bitb_23_22 word23_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_22 q_24_22 qb_24_22 bit_24_22 bitb_24_22 word24_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_22 q_25_22 qb_25_22 bit_25_22 bitb_25_22 word25_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_22 q_26_22 qb_26_22 bit_26_22 bitb_26_22 word26_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_22 q_27_22 qb_27_22 bit_27_22 bitb_27_22 word27_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_22 q_28_22 qb_28_22 bit_28_22 bitb_28_22 word28_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_22 q_29_22 qb_29_22 bit_29_22 bitb_29_22 word29_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_22 q_30_22 qb_30_22 bit_30_22 bitb_30_22 word30_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_22 q_31_22 qb_31_22 bit_31_22 bitb_31_22 word31_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_22 q_32_22 qb_32_22 bit_32_22 bitb_32_22 word32_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_22 q_33_22 qb_33_22 bit_33_22 bitb_33_22 word33_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_22 q_34_22 qb_34_22 bit_34_22 bitb_34_22 word34_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_22 q_35_22 qb_35_22 bit_35_22 bitb_35_22 word35_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_22 q_36_22 qb_36_22 bit_36_22 bitb_36_22 word36_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_22 q_37_22 qb_37_22 bit_37_22 bitb_37_22 word37_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_22 q_38_22 qb_38_22 bit_38_22 bitb_38_22 word38_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_22 q_39_22 qb_39_22 bit_39_22 bitb_39_22 word39_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_22 q_40_22 qb_40_22 bit_40_22 bitb_40_22 word40_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_22 q_41_22 qb_41_22 bit_41_22 bitb_41_22 word41_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_22 q_42_22 qb_42_22 bit_42_22 bitb_42_22 word42_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_22 q_43_22 qb_43_22 bit_43_22 bitb_43_22 word43_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_22 q_44_22 qb_44_22 bit_44_22 bitb_44_22 word44_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_22 q_45_22 qb_45_22 bit_45_22 bitb_45_22 word45_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_22 q_46_22 qb_46_22 bit_46_22 bitb_46_22 word46_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_22 q_47_22 qb_47_22 bit_47_22 bitb_47_22 word47_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_22 q_48_22 qb_48_22 bit_48_22 bitb_48_22 word48_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_22 q_49_22 qb_49_22 bit_49_22 bitb_49_22 word49_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_22 q_50_22 qb_50_22 bit_50_22 bitb_50_22 word50_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_22 q_51_22 qb_51_22 bit_51_22 bitb_51_22 word51_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_22 q_52_22 qb_52_22 bit_52_22 bitb_52_22 word52_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_22 q_53_22 qb_53_22 bit_53_22 bitb_53_22 word53_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_22 q_54_22 qb_54_22 bit_54_22 bitb_54_22 word54_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_22 q_55_22 qb_55_22 bit_55_22 bitb_55_22 word55_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_22 q_56_22 qb_56_22 bit_56_22 bitb_56_22 word56_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_22 q_57_22 qb_57_22 bit_57_22 bitb_57_22 word57_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_22 q_58_22 qb_58_22 bit_58_22 bitb_58_22 word58_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_22 q_59_22 qb_59_22 bit_59_22 bitb_59_22 word59_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_22 q_60_22 qb_60_22 bit_60_22 bitb_60_22 word60_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_22 q_61_22 qb_61_22 bit_61_22 bitb_61_22 word61_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_22 q_62_22 qb_62_22 bit_62_22 bitb_62_22 word62_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_22 q_63_22 qb_63_22 bit_63_22 bitb_63_22 word63_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_22 q_64_22 qb_64_22 bit_64_22 bitb_64_22 word64_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_22 q_65_22 qb_65_22 bit_65_22 bitb_65_22 word65_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_22 q_66_22 qb_66_22 bit_66_22 bitb_66_22 word66_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_22 q_67_22 qb_67_22 bit_67_22 bitb_67_22 word67_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_22 q_68_22 qb_68_22 bit_68_22 bitb_68_22 word68_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_22 q_69_22 qb_69_22 bit_69_22 bitb_69_22 word69_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_22 q_70_22 qb_70_22 bit_70_22 bitb_70_22 word70_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_22 q_71_22 qb_71_22 bit_71_22 bitb_71_22 word71_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_22 q_72_22 qb_72_22 bit_72_22 bitb_72_22 word72_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_22 q_73_22 qb_73_22 bit_73_22 bitb_73_22 word73_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_22 q_74_22 qb_74_22 bit_74_22 bitb_74_22 word74_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_22 q_75_22 qb_75_22 bit_75_22 bitb_75_22 word75_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_22 q_76_22 qb_76_22 bit_76_22 bitb_76_22 word76_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_22 q_77_22 qb_77_22 bit_77_22 bitb_77_22 word77_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_22 q_78_22 qb_78_22 bit_78_22 bitb_78_22 word78_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_22 q_79_22 qb_79_22 bit_79_22 bitb_79_22 word79_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_22 q_80_22 qb_80_22 bit_80_22 bitb_80_22 word80_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_22 q_81_22 qb_81_22 bit_81_22 bitb_81_22 word81_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_22 q_82_22 qb_82_22 bit_82_22 bitb_82_22 word82_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_22 q_83_22 qb_83_22 bit_83_22 bitb_83_22 word83_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_22 q_84_22 qb_84_22 bit_84_22 bitb_84_22 word84_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_22 q_85_22 qb_85_22 bit_85_22 bitb_85_22 word85_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_22 q_86_22 qb_86_22 bit_86_22 bitb_86_22 word86_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_22 q_87_22 qb_87_22 bit_87_22 bitb_87_22 word87_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_22 q_88_22 qb_88_22 bit_88_22 bitb_88_22 word88_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_22 q_89_22 qb_89_22 bit_89_22 bitb_89_22 word89_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_22 q_90_22 qb_90_22 bit_90_22 bitb_90_22 word90_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_22 q_91_22 qb_91_22 bit_91_22 bitb_91_22 word91_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_22 q_92_22 qb_92_22 bit_92_22 bitb_92_22 word92_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_22 q_93_22 qb_93_22 bit_93_22 bitb_93_22 word93_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_22 q_94_22 qb_94_22 bit_94_22 bitb_94_22 word94_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_22 q_95_22 qb_95_22 bit_95_22 bitb_95_22 word95_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_22 q_96_22 qb_96_22 bit_96_22 bitb_96_22 word96_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_22 q_97_22 qb_97_22 bit_97_22 bitb_97_22 word97_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_22 q_98_22 qb_98_22 bit_98_22 bitb_98_22 word98_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_22 q_99_22 qb_99_22 bit_99_22 bitb_99_22 word99_22 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_23 q_0_23 qb_0_23 bit_0_23 bitb_0_23 word0_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_23 q_1_23 qb_1_23 bit_1_23 bitb_1_23 word1_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_23 q_2_23 qb_2_23 bit_2_23 bitb_2_23 word2_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_23 q_3_23 qb_3_23 bit_3_23 bitb_3_23 word3_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_23 q_4_23 qb_4_23 bit_4_23 bitb_4_23 word4_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_23 q_5_23 qb_5_23 bit_5_23 bitb_5_23 word5_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_23 q_6_23 qb_6_23 bit_6_23 bitb_6_23 word6_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_23 q_7_23 qb_7_23 bit_7_23 bitb_7_23 word7_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_23 q_8_23 qb_8_23 bit_8_23 bitb_8_23 word8_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_23 q_9_23 qb_9_23 bit_9_23 bitb_9_23 word9_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_23 q_10_23 qb_10_23 bit_10_23 bitb_10_23 word10_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_23 q_11_23 qb_11_23 bit_11_23 bitb_11_23 word11_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_23 q_12_23 qb_12_23 bit_12_23 bitb_12_23 word12_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_23 q_13_23 qb_13_23 bit_13_23 bitb_13_23 word13_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_23 q_14_23 qb_14_23 bit_14_23 bitb_14_23 word14_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_23 q_15_23 qb_15_23 bit_15_23 bitb_15_23 word15_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_23 q_16_23 qb_16_23 bit_16_23 bitb_16_23 word16_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_23 q_17_23 qb_17_23 bit_17_23 bitb_17_23 word17_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_23 q_18_23 qb_18_23 bit_18_23 bitb_18_23 word18_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_23 q_19_23 qb_19_23 bit_19_23 bitb_19_23 word19_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_23 q_20_23 qb_20_23 bit_20_23 bitb_20_23 word20_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_23 q_21_23 qb_21_23 bit_21_23 bitb_21_23 word21_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_23 q_22_23 qb_22_23 bit_22_23 bitb_22_23 word22_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_23 q_23_23 qb_23_23 bit_23_23 bitb_23_23 word23_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_23 q_24_23 qb_24_23 bit_24_23 bitb_24_23 word24_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_23 q_25_23 qb_25_23 bit_25_23 bitb_25_23 word25_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_23 q_26_23 qb_26_23 bit_26_23 bitb_26_23 word26_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_23 q_27_23 qb_27_23 bit_27_23 bitb_27_23 word27_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_23 q_28_23 qb_28_23 bit_28_23 bitb_28_23 word28_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_23 q_29_23 qb_29_23 bit_29_23 bitb_29_23 word29_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_23 q_30_23 qb_30_23 bit_30_23 bitb_30_23 word30_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_23 q_31_23 qb_31_23 bit_31_23 bitb_31_23 word31_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_23 q_32_23 qb_32_23 bit_32_23 bitb_32_23 word32_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_23 q_33_23 qb_33_23 bit_33_23 bitb_33_23 word33_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_23 q_34_23 qb_34_23 bit_34_23 bitb_34_23 word34_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_23 q_35_23 qb_35_23 bit_35_23 bitb_35_23 word35_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_23 q_36_23 qb_36_23 bit_36_23 bitb_36_23 word36_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_23 q_37_23 qb_37_23 bit_37_23 bitb_37_23 word37_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_23 q_38_23 qb_38_23 bit_38_23 bitb_38_23 word38_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_23 q_39_23 qb_39_23 bit_39_23 bitb_39_23 word39_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_23 q_40_23 qb_40_23 bit_40_23 bitb_40_23 word40_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_23 q_41_23 qb_41_23 bit_41_23 bitb_41_23 word41_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_23 q_42_23 qb_42_23 bit_42_23 bitb_42_23 word42_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_23 q_43_23 qb_43_23 bit_43_23 bitb_43_23 word43_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_23 q_44_23 qb_44_23 bit_44_23 bitb_44_23 word44_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_23 q_45_23 qb_45_23 bit_45_23 bitb_45_23 word45_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_23 q_46_23 qb_46_23 bit_46_23 bitb_46_23 word46_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_23 q_47_23 qb_47_23 bit_47_23 bitb_47_23 word47_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_23 q_48_23 qb_48_23 bit_48_23 bitb_48_23 word48_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_23 q_49_23 qb_49_23 bit_49_23 bitb_49_23 word49_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_23 q_50_23 qb_50_23 bit_50_23 bitb_50_23 word50_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_23 q_51_23 qb_51_23 bit_51_23 bitb_51_23 word51_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_23 q_52_23 qb_52_23 bit_52_23 bitb_52_23 word52_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_23 q_53_23 qb_53_23 bit_53_23 bitb_53_23 word53_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_23 q_54_23 qb_54_23 bit_54_23 bitb_54_23 word54_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_23 q_55_23 qb_55_23 bit_55_23 bitb_55_23 word55_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_23 q_56_23 qb_56_23 bit_56_23 bitb_56_23 word56_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_23 q_57_23 qb_57_23 bit_57_23 bitb_57_23 word57_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_23 q_58_23 qb_58_23 bit_58_23 bitb_58_23 word58_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_23 q_59_23 qb_59_23 bit_59_23 bitb_59_23 word59_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_23 q_60_23 qb_60_23 bit_60_23 bitb_60_23 word60_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_23 q_61_23 qb_61_23 bit_61_23 bitb_61_23 word61_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_23 q_62_23 qb_62_23 bit_62_23 bitb_62_23 word62_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_23 q_63_23 qb_63_23 bit_63_23 bitb_63_23 word63_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_23 q_64_23 qb_64_23 bit_64_23 bitb_64_23 word64_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_23 q_65_23 qb_65_23 bit_65_23 bitb_65_23 word65_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_23 q_66_23 qb_66_23 bit_66_23 bitb_66_23 word66_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_23 q_67_23 qb_67_23 bit_67_23 bitb_67_23 word67_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_23 q_68_23 qb_68_23 bit_68_23 bitb_68_23 word68_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_23 q_69_23 qb_69_23 bit_69_23 bitb_69_23 word69_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_23 q_70_23 qb_70_23 bit_70_23 bitb_70_23 word70_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_23 q_71_23 qb_71_23 bit_71_23 bitb_71_23 word71_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_23 q_72_23 qb_72_23 bit_72_23 bitb_72_23 word72_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_23 q_73_23 qb_73_23 bit_73_23 bitb_73_23 word73_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_23 q_74_23 qb_74_23 bit_74_23 bitb_74_23 word74_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_23 q_75_23 qb_75_23 bit_75_23 bitb_75_23 word75_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_23 q_76_23 qb_76_23 bit_76_23 bitb_76_23 word76_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_23 q_77_23 qb_77_23 bit_77_23 bitb_77_23 word77_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_23 q_78_23 qb_78_23 bit_78_23 bitb_78_23 word78_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_23 q_79_23 qb_79_23 bit_79_23 bitb_79_23 word79_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_23 q_80_23 qb_80_23 bit_80_23 bitb_80_23 word80_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_23 q_81_23 qb_81_23 bit_81_23 bitb_81_23 word81_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_23 q_82_23 qb_82_23 bit_82_23 bitb_82_23 word82_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_23 q_83_23 qb_83_23 bit_83_23 bitb_83_23 word83_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_23 q_84_23 qb_84_23 bit_84_23 bitb_84_23 word84_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_23 q_85_23 qb_85_23 bit_85_23 bitb_85_23 word85_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_23 q_86_23 qb_86_23 bit_86_23 bitb_86_23 word86_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_23 q_87_23 qb_87_23 bit_87_23 bitb_87_23 word87_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_23 q_88_23 qb_88_23 bit_88_23 bitb_88_23 word88_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_23 q_89_23 qb_89_23 bit_89_23 bitb_89_23 word89_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_23 q_90_23 qb_90_23 bit_90_23 bitb_90_23 word90_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_23 q_91_23 qb_91_23 bit_91_23 bitb_91_23 word91_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_23 q_92_23 qb_92_23 bit_92_23 bitb_92_23 word92_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_23 q_93_23 qb_93_23 bit_93_23 bitb_93_23 word93_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_23 q_94_23 qb_94_23 bit_94_23 bitb_94_23 word94_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_23 q_95_23 qb_95_23 bit_95_23 bitb_95_23 word95_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_23 q_96_23 qb_96_23 bit_96_23 bitb_96_23 word96_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_23 q_97_23 qb_97_23 bit_97_23 bitb_97_23 word97_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_23 q_98_23 qb_98_23 bit_98_23 bitb_98_23 word98_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_23 q_99_23 qb_99_23 bit_99_23 bitb_99_23 word99_23 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_24 q_0_24 qb_0_24 bit_0_24 bitb_0_24 word0_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_24 q_1_24 qb_1_24 bit_1_24 bitb_1_24 word1_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_24 q_2_24 qb_2_24 bit_2_24 bitb_2_24 word2_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_24 q_3_24 qb_3_24 bit_3_24 bitb_3_24 word3_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_24 q_4_24 qb_4_24 bit_4_24 bitb_4_24 word4_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_24 q_5_24 qb_5_24 bit_5_24 bitb_5_24 word5_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_24 q_6_24 qb_6_24 bit_6_24 bitb_6_24 word6_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_24 q_7_24 qb_7_24 bit_7_24 bitb_7_24 word7_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_24 q_8_24 qb_8_24 bit_8_24 bitb_8_24 word8_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_24 q_9_24 qb_9_24 bit_9_24 bitb_9_24 word9_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_24 q_10_24 qb_10_24 bit_10_24 bitb_10_24 word10_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_24 q_11_24 qb_11_24 bit_11_24 bitb_11_24 word11_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_24 q_12_24 qb_12_24 bit_12_24 bitb_12_24 word12_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_24 q_13_24 qb_13_24 bit_13_24 bitb_13_24 word13_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_24 q_14_24 qb_14_24 bit_14_24 bitb_14_24 word14_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_24 q_15_24 qb_15_24 bit_15_24 bitb_15_24 word15_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_24 q_16_24 qb_16_24 bit_16_24 bitb_16_24 word16_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_24 q_17_24 qb_17_24 bit_17_24 bitb_17_24 word17_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_24 q_18_24 qb_18_24 bit_18_24 bitb_18_24 word18_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_24 q_19_24 qb_19_24 bit_19_24 bitb_19_24 word19_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_24 q_20_24 qb_20_24 bit_20_24 bitb_20_24 word20_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_24 q_21_24 qb_21_24 bit_21_24 bitb_21_24 word21_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_24 q_22_24 qb_22_24 bit_22_24 bitb_22_24 word22_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_24 q_23_24 qb_23_24 bit_23_24 bitb_23_24 word23_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_24 q_24_24 qb_24_24 bit_24_24 bitb_24_24 word24_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_24 q_25_24 qb_25_24 bit_25_24 bitb_25_24 word25_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_24 q_26_24 qb_26_24 bit_26_24 bitb_26_24 word26_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_24 q_27_24 qb_27_24 bit_27_24 bitb_27_24 word27_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_24 q_28_24 qb_28_24 bit_28_24 bitb_28_24 word28_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_24 q_29_24 qb_29_24 bit_29_24 bitb_29_24 word29_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_24 q_30_24 qb_30_24 bit_30_24 bitb_30_24 word30_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_24 q_31_24 qb_31_24 bit_31_24 bitb_31_24 word31_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_24 q_32_24 qb_32_24 bit_32_24 bitb_32_24 word32_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_24 q_33_24 qb_33_24 bit_33_24 bitb_33_24 word33_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_24 q_34_24 qb_34_24 bit_34_24 bitb_34_24 word34_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_24 q_35_24 qb_35_24 bit_35_24 bitb_35_24 word35_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_24 q_36_24 qb_36_24 bit_36_24 bitb_36_24 word36_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_24 q_37_24 qb_37_24 bit_37_24 bitb_37_24 word37_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_24 q_38_24 qb_38_24 bit_38_24 bitb_38_24 word38_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_24 q_39_24 qb_39_24 bit_39_24 bitb_39_24 word39_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_24 q_40_24 qb_40_24 bit_40_24 bitb_40_24 word40_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_24 q_41_24 qb_41_24 bit_41_24 bitb_41_24 word41_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_24 q_42_24 qb_42_24 bit_42_24 bitb_42_24 word42_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_24 q_43_24 qb_43_24 bit_43_24 bitb_43_24 word43_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_24 q_44_24 qb_44_24 bit_44_24 bitb_44_24 word44_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_24 q_45_24 qb_45_24 bit_45_24 bitb_45_24 word45_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_24 q_46_24 qb_46_24 bit_46_24 bitb_46_24 word46_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_24 q_47_24 qb_47_24 bit_47_24 bitb_47_24 word47_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_24 q_48_24 qb_48_24 bit_48_24 bitb_48_24 word48_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_24 q_49_24 qb_49_24 bit_49_24 bitb_49_24 word49_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_24 q_50_24 qb_50_24 bit_50_24 bitb_50_24 word50_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_24 q_51_24 qb_51_24 bit_51_24 bitb_51_24 word51_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_24 q_52_24 qb_52_24 bit_52_24 bitb_52_24 word52_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_24 q_53_24 qb_53_24 bit_53_24 bitb_53_24 word53_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_24 q_54_24 qb_54_24 bit_54_24 bitb_54_24 word54_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_24 q_55_24 qb_55_24 bit_55_24 bitb_55_24 word55_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_24 q_56_24 qb_56_24 bit_56_24 bitb_56_24 word56_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_24 q_57_24 qb_57_24 bit_57_24 bitb_57_24 word57_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_24 q_58_24 qb_58_24 bit_58_24 bitb_58_24 word58_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_24 q_59_24 qb_59_24 bit_59_24 bitb_59_24 word59_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_24 q_60_24 qb_60_24 bit_60_24 bitb_60_24 word60_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_24 q_61_24 qb_61_24 bit_61_24 bitb_61_24 word61_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_24 q_62_24 qb_62_24 bit_62_24 bitb_62_24 word62_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_24 q_63_24 qb_63_24 bit_63_24 bitb_63_24 word63_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_24 q_64_24 qb_64_24 bit_64_24 bitb_64_24 word64_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_24 q_65_24 qb_65_24 bit_65_24 bitb_65_24 word65_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_24 q_66_24 qb_66_24 bit_66_24 bitb_66_24 word66_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_24 q_67_24 qb_67_24 bit_67_24 bitb_67_24 word67_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_24 q_68_24 qb_68_24 bit_68_24 bitb_68_24 word68_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_24 q_69_24 qb_69_24 bit_69_24 bitb_69_24 word69_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_24 q_70_24 qb_70_24 bit_70_24 bitb_70_24 word70_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_24 q_71_24 qb_71_24 bit_71_24 bitb_71_24 word71_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_24 q_72_24 qb_72_24 bit_72_24 bitb_72_24 word72_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_24 q_73_24 qb_73_24 bit_73_24 bitb_73_24 word73_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_24 q_74_24 qb_74_24 bit_74_24 bitb_74_24 word74_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_24 q_75_24 qb_75_24 bit_75_24 bitb_75_24 word75_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_24 q_76_24 qb_76_24 bit_76_24 bitb_76_24 word76_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_24 q_77_24 qb_77_24 bit_77_24 bitb_77_24 word77_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_24 q_78_24 qb_78_24 bit_78_24 bitb_78_24 word78_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_24 q_79_24 qb_79_24 bit_79_24 bitb_79_24 word79_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_24 q_80_24 qb_80_24 bit_80_24 bitb_80_24 word80_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_24 q_81_24 qb_81_24 bit_81_24 bitb_81_24 word81_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_24 q_82_24 qb_82_24 bit_82_24 bitb_82_24 word82_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_24 q_83_24 qb_83_24 bit_83_24 bitb_83_24 word83_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_24 q_84_24 qb_84_24 bit_84_24 bitb_84_24 word84_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_24 q_85_24 qb_85_24 bit_85_24 bitb_85_24 word85_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_24 q_86_24 qb_86_24 bit_86_24 bitb_86_24 word86_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_24 q_87_24 qb_87_24 bit_87_24 bitb_87_24 word87_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_24 q_88_24 qb_88_24 bit_88_24 bitb_88_24 word88_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_24 q_89_24 qb_89_24 bit_89_24 bitb_89_24 word89_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_24 q_90_24 qb_90_24 bit_90_24 bitb_90_24 word90_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_24 q_91_24 qb_91_24 bit_91_24 bitb_91_24 word91_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_24 q_92_24 qb_92_24 bit_92_24 bitb_92_24 word92_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_24 q_93_24 qb_93_24 bit_93_24 bitb_93_24 word93_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_24 q_94_24 qb_94_24 bit_94_24 bitb_94_24 word94_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_24 q_95_24 qb_95_24 bit_95_24 bitb_95_24 word95_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_24 q_96_24 qb_96_24 bit_96_24 bitb_96_24 word96_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_24 q_97_24 qb_97_24 bit_97_24 bitb_97_24 word97_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_24 q_98_24 qb_98_24 bit_98_24 bitb_98_24 word98_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_24 q_99_24 qb_99_24 bit_99_24 bitb_99_24 word99_24 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_25 q_0_25 qb_0_25 bit_0_25 bitb_0_25 word0_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_25 q_1_25 qb_1_25 bit_1_25 bitb_1_25 word1_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_25 q_2_25 qb_2_25 bit_2_25 bitb_2_25 word2_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_25 q_3_25 qb_3_25 bit_3_25 bitb_3_25 word3_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_25 q_4_25 qb_4_25 bit_4_25 bitb_4_25 word4_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_25 q_5_25 qb_5_25 bit_5_25 bitb_5_25 word5_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_25 q_6_25 qb_6_25 bit_6_25 bitb_6_25 word6_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_25 q_7_25 qb_7_25 bit_7_25 bitb_7_25 word7_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_25 q_8_25 qb_8_25 bit_8_25 bitb_8_25 word8_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_25 q_9_25 qb_9_25 bit_9_25 bitb_9_25 word9_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_25 q_10_25 qb_10_25 bit_10_25 bitb_10_25 word10_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_25 q_11_25 qb_11_25 bit_11_25 bitb_11_25 word11_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_25 q_12_25 qb_12_25 bit_12_25 bitb_12_25 word12_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_25 q_13_25 qb_13_25 bit_13_25 bitb_13_25 word13_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_25 q_14_25 qb_14_25 bit_14_25 bitb_14_25 word14_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_25 q_15_25 qb_15_25 bit_15_25 bitb_15_25 word15_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_25 q_16_25 qb_16_25 bit_16_25 bitb_16_25 word16_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_25 q_17_25 qb_17_25 bit_17_25 bitb_17_25 word17_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_25 q_18_25 qb_18_25 bit_18_25 bitb_18_25 word18_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_25 q_19_25 qb_19_25 bit_19_25 bitb_19_25 word19_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_25 q_20_25 qb_20_25 bit_20_25 bitb_20_25 word20_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_25 q_21_25 qb_21_25 bit_21_25 bitb_21_25 word21_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_25 q_22_25 qb_22_25 bit_22_25 bitb_22_25 word22_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_25 q_23_25 qb_23_25 bit_23_25 bitb_23_25 word23_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_25 q_24_25 qb_24_25 bit_24_25 bitb_24_25 word24_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_25 q_25_25 qb_25_25 bit_25_25 bitb_25_25 word25_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_25 q_26_25 qb_26_25 bit_26_25 bitb_26_25 word26_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_25 q_27_25 qb_27_25 bit_27_25 bitb_27_25 word27_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_25 q_28_25 qb_28_25 bit_28_25 bitb_28_25 word28_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_25 q_29_25 qb_29_25 bit_29_25 bitb_29_25 word29_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_25 q_30_25 qb_30_25 bit_30_25 bitb_30_25 word30_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_25 q_31_25 qb_31_25 bit_31_25 bitb_31_25 word31_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_25 q_32_25 qb_32_25 bit_32_25 bitb_32_25 word32_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_25 q_33_25 qb_33_25 bit_33_25 bitb_33_25 word33_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_25 q_34_25 qb_34_25 bit_34_25 bitb_34_25 word34_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_25 q_35_25 qb_35_25 bit_35_25 bitb_35_25 word35_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_25 q_36_25 qb_36_25 bit_36_25 bitb_36_25 word36_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_25 q_37_25 qb_37_25 bit_37_25 bitb_37_25 word37_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_25 q_38_25 qb_38_25 bit_38_25 bitb_38_25 word38_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_25 q_39_25 qb_39_25 bit_39_25 bitb_39_25 word39_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_25 q_40_25 qb_40_25 bit_40_25 bitb_40_25 word40_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_25 q_41_25 qb_41_25 bit_41_25 bitb_41_25 word41_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_25 q_42_25 qb_42_25 bit_42_25 bitb_42_25 word42_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_25 q_43_25 qb_43_25 bit_43_25 bitb_43_25 word43_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_25 q_44_25 qb_44_25 bit_44_25 bitb_44_25 word44_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_25 q_45_25 qb_45_25 bit_45_25 bitb_45_25 word45_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_25 q_46_25 qb_46_25 bit_46_25 bitb_46_25 word46_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_25 q_47_25 qb_47_25 bit_47_25 bitb_47_25 word47_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_25 q_48_25 qb_48_25 bit_48_25 bitb_48_25 word48_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_25 q_49_25 qb_49_25 bit_49_25 bitb_49_25 word49_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_25 q_50_25 qb_50_25 bit_50_25 bitb_50_25 word50_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_25 q_51_25 qb_51_25 bit_51_25 bitb_51_25 word51_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_25 q_52_25 qb_52_25 bit_52_25 bitb_52_25 word52_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_25 q_53_25 qb_53_25 bit_53_25 bitb_53_25 word53_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_25 q_54_25 qb_54_25 bit_54_25 bitb_54_25 word54_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_25 q_55_25 qb_55_25 bit_55_25 bitb_55_25 word55_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_25 q_56_25 qb_56_25 bit_56_25 bitb_56_25 word56_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_25 q_57_25 qb_57_25 bit_57_25 bitb_57_25 word57_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_25 q_58_25 qb_58_25 bit_58_25 bitb_58_25 word58_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_25 q_59_25 qb_59_25 bit_59_25 bitb_59_25 word59_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_25 q_60_25 qb_60_25 bit_60_25 bitb_60_25 word60_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_25 q_61_25 qb_61_25 bit_61_25 bitb_61_25 word61_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_25 q_62_25 qb_62_25 bit_62_25 bitb_62_25 word62_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_25 q_63_25 qb_63_25 bit_63_25 bitb_63_25 word63_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_25 q_64_25 qb_64_25 bit_64_25 bitb_64_25 word64_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_25 q_65_25 qb_65_25 bit_65_25 bitb_65_25 word65_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_25 q_66_25 qb_66_25 bit_66_25 bitb_66_25 word66_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_25 q_67_25 qb_67_25 bit_67_25 bitb_67_25 word67_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_25 q_68_25 qb_68_25 bit_68_25 bitb_68_25 word68_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_25 q_69_25 qb_69_25 bit_69_25 bitb_69_25 word69_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_25 q_70_25 qb_70_25 bit_70_25 bitb_70_25 word70_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_25 q_71_25 qb_71_25 bit_71_25 bitb_71_25 word71_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_25 q_72_25 qb_72_25 bit_72_25 bitb_72_25 word72_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_25 q_73_25 qb_73_25 bit_73_25 bitb_73_25 word73_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_25 q_74_25 qb_74_25 bit_74_25 bitb_74_25 word74_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_25 q_75_25 qb_75_25 bit_75_25 bitb_75_25 word75_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_25 q_76_25 qb_76_25 bit_76_25 bitb_76_25 word76_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_25 q_77_25 qb_77_25 bit_77_25 bitb_77_25 word77_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_25 q_78_25 qb_78_25 bit_78_25 bitb_78_25 word78_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_25 q_79_25 qb_79_25 bit_79_25 bitb_79_25 word79_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_25 q_80_25 qb_80_25 bit_80_25 bitb_80_25 word80_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_25 q_81_25 qb_81_25 bit_81_25 bitb_81_25 word81_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_25 q_82_25 qb_82_25 bit_82_25 bitb_82_25 word82_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_25 q_83_25 qb_83_25 bit_83_25 bitb_83_25 word83_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_25 q_84_25 qb_84_25 bit_84_25 bitb_84_25 word84_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_25 q_85_25 qb_85_25 bit_85_25 bitb_85_25 word85_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_25 q_86_25 qb_86_25 bit_86_25 bitb_86_25 word86_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_25 q_87_25 qb_87_25 bit_87_25 bitb_87_25 word87_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_25 q_88_25 qb_88_25 bit_88_25 bitb_88_25 word88_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_25 q_89_25 qb_89_25 bit_89_25 bitb_89_25 word89_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_25 q_90_25 qb_90_25 bit_90_25 bitb_90_25 word90_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_25 q_91_25 qb_91_25 bit_91_25 bitb_91_25 word91_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_25 q_92_25 qb_92_25 bit_92_25 bitb_92_25 word92_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_25 q_93_25 qb_93_25 bit_93_25 bitb_93_25 word93_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_25 q_94_25 qb_94_25 bit_94_25 bitb_94_25 word94_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_25 q_95_25 qb_95_25 bit_95_25 bitb_95_25 word95_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_25 q_96_25 qb_96_25 bit_96_25 bitb_96_25 word96_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_25 q_97_25 qb_97_25 bit_97_25 bitb_97_25 word97_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_25 q_98_25 qb_98_25 bit_98_25 bitb_98_25 word98_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_25 q_99_25 qb_99_25 bit_99_25 bitb_99_25 word99_25 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_26 q_0_26 qb_0_26 bit_0_26 bitb_0_26 word0_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_26 q_1_26 qb_1_26 bit_1_26 bitb_1_26 word1_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_26 q_2_26 qb_2_26 bit_2_26 bitb_2_26 word2_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_26 q_3_26 qb_3_26 bit_3_26 bitb_3_26 word3_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_26 q_4_26 qb_4_26 bit_4_26 bitb_4_26 word4_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_26 q_5_26 qb_5_26 bit_5_26 bitb_5_26 word5_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_26 q_6_26 qb_6_26 bit_6_26 bitb_6_26 word6_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_26 q_7_26 qb_7_26 bit_7_26 bitb_7_26 word7_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_26 q_8_26 qb_8_26 bit_8_26 bitb_8_26 word8_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_26 q_9_26 qb_9_26 bit_9_26 bitb_9_26 word9_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_26 q_10_26 qb_10_26 bit_10_26 bitb_10_26 word10_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_26 q_11_26 qb_11_26 bit_11_26 bitb_11_26 word11_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_26 q_12_26 qb_12_26 bit_12_26 bitb_12_26 word12_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_26 q_13_26 qb_13_26 bit_13_26 bitb_13_26 word13_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_26 q_14_26 qb_14_26 bit_14_26 bitb_14_26 word14_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_26 q_15_26 qb_15_26 bit_15_26 bitb_15_26 word15_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_26 q_16_26 qb_16_26 bit_16_26 bitb_16_26 word16_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_26 q_17_26 qb_17_26 bit_17_26 bitb_17_26 word17_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_26 q_18_26 qb_18_26 bit_18_26 bitb_18_26 word18_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_26 q_19_26 qb_19_26 bit_19_26 bitb_19_26 word19_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_26 q_20_26 qb_20_26 bit_20_26 bitb_20_26 word20_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_26 q_21_26 qb_21_26 bit_21_26 bitb_21_26 word21_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_26 q_22_26 qb_22_26 bit_22_26 bitb_22_26 word22_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_26 q_23_26 qb_23_26 bit_23_26 bitb_23_26 word23_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_26 q_24_26 qb_24_26 bit_24_26 bitb_24_26 word24_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_26 q_25_26 qb_25_26 bit_25_26 bitb_25_26 word25_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_26 q_26_26 qb_26_26 bit_26_26 bitb_26_26 word26_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_26 q_27_26 qb_27_26 bit_27_26 bitb_27_26 word27_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_26 q_28_26 qb_28_26 bit_28_26 bitb_28_26 word28_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_26 q_29_26 qb_29_26 bit_29_26 bitb_29_26 word29_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_26 q_30_26 qb_30_26 bit_30_26 bitb_30_26 word30_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_26 q_31_26 qb_31_26 bit_31_26 bitb_31_26 word31_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_26 q_32_26 qb_32_26 bit_32_26 bitb_32_26 word32_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_26 q_33_26 qb_33_26 bit_33_26 bitb_33_26 word33_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_26 q_34_26 qb_34_26 bit_34_26 bitb_34_26 word34_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_26 q_35_26 qb_35_26 bit_35_26 bitb_35_26 word35_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_26 q_36_26 qb_36_26 bit_36_26 bitb_36_26 word36_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_26 q_37_26 qb_37_26 bit_37_26 bitb_37_26 word37_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_26 q_38_26 qb_38_26 bit_38_26 bitb_38_26 word38_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_26 q_39_26 qb_39_26 bit_39_26 bitb_39_26 word39_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_26 q_40_26 qb_40_26 bit_40_26 bitb_40_26 word40_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_26 q_41_26 qb_41_26 bit_41_26 bitb_41_26 word41_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_26 q_42_26 qb_42_26 bit_42_26 bitb_42_26 word42_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_26 q_43_26 qb_43_26 bit_43_26 bitb_43_26 word43_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_26 q_44_26 qb_44_26 bit_44_26 bitb_44_26 word44_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_26 q_45_26 qb_45_26 bit_45_26 bitb_45_26 word45_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_26 q_46_26 qb_46_26 bit_46_26 bitb_46_26 word46_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_26 q_47_26 qb_47_26 bit_47_26 bitb_47_26 word47_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_26 q_48_26 qb_48_26 bit_48_26 bitb_48_26 word48_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_26 q_49_26 qb_49_26 bit_49_26 bitb_49_26 word49_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_26 q_50_26 qb_50_26 bit_50_26 bitb_50_26 word50_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_26 q_51_26 qb_51_26 bit_51_26 bitb_51_26 word51_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_26 q_52_26 qb_52_26 bit_52_26 bitb_52_26 word52_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_26 q_53_26 qb_53_26 bit_53_26 bitb_53_26 word53_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_26 q_54_26 qb_54_26 bit_54_26 bitb_54_26 word54_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_26 q_55_26 qb_55_26 bit_55_26 bitb_55_26 word55_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_26 q_56_26 qb_56_26 bit_56_26 bitb_56_26 word56_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_26 q_57_26 qb_57_26 bit_57_26 bitb_57_26 word57_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_26 q_58_26 qb_58_26 bit_58_26 bitb_58_26 word58_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_26 q_59_26 qb_59_26 bit_59_26 bitb_59_26 word59_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_26 q_60_26 qb_60_26 bit_60_26 bitb_60_26 word60_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_26 q_61_26 qb_61_26 bit_61_26 bitb_61_26 word61_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_26 q_62_26 qb_62_26 bit_62_26 bitb_62_26 word62_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_26 q_63_26 qb_63_26 bit_63_26 bitb_63_26 word63_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_26 q_64_26 qb_64_26 bit_64_26 bitb_64_26 word64_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_26 q_65_26 qb_65_26 bit_65_26 bitb_65_26 word65_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_26 q_66_26 qb_66_26 bit_66_26 bitb_66_26 word66_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_26 q_67_26 qb_67_26 bit_67_26 bitb_67_26 word67_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_26 q_68_26 qb_68_26 bit_68_26 bitb_68_26 word68_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_26 q_69_26 qb_69_26 bit_69_26 bitb_69_26 word69_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_26 q_70_26 qb_70_26 bit_70_26 bitb_70_26 word70_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_26 q_71_26 qb_71_26 bit_71_26 bitb_71_26 word71_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_26 q_72_26 qb_72_26 bit_72_26 bitb_72_26 word72_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_26 q_73_26 qb_73_26 bit_73_26 bitb_73_26 word73_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_26 q_74_26 qb_74_26 bit_74_26 bitb_74_26 word74_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_26 q_75_26 qb_75_26 bit_75_26 bitb_75_26 word75_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_26 q_76_26 qb_76_26 bit_76_26 bitb_76_26 word76_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_26 q_77_26 qb_77_26 bit_77_26 bitb_77_26 word77_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_26 q_78_26 qb_78_26 bit_78_26 bitb_78_26 word78_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_26 q_79_26 qb_79_26 bit_79_26 bitb_79_26 word79_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_26 q_80_26 qb_80_26 bit_80_26 bitb_80_26 word80_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_26 q_81_26 qb_81_26 bit_81_26 bitb_81_26 word81_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_26 q_82_26 qb_82_26 bit_82_26 bitb_82_26 word82_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_26 q_83_26 qb_83_26 bit_83_26 bitb_83_26 word83_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_26 q_84_26 qb_84_26 bit_84_26 bitb_84_26 word84_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_26 q_85_26 qb_85_26 bit_85_26 bitb_85_26 word85_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_26 q_86_26 qb_86_26 bit_86_26 bitb_86_26 word86_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_26 q_87_26 qb_87_26 bit_87_26 bitb_87_26 word87_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_26 q_88_26 qb_88_26 bit_88_26 bitb_88_26 word88_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_26 q_89_26 qb_89_26 bit_89_26 bitb_89_26 word89_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_26 q_90_26 qb_90_26 bit_90_26 bitb_90_26 word90_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_26 q_91_26 qb_91_26 bit_91_26 bitb_91_26 word91_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_26 q_92_26 qb_92_26 bit_92_26 bitb_92_26 word92_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_26 q_93_26 qb_93_26 bit_93_26 bitb_93_26 word93_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_26 q_94_26 qb_94_26 bit_94_26 bitb_94_26 word94_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_26 q_95_26 qb_95_26 bit_95_26 bitb_95_26 word95_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_26 q_96_26 qb_96_26 bit_96_26 bitb_96_26 word96_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_26 q_97_26 qb_97_26 bit_97_26 bitb_97_26 word97_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_26 q_98_26 qb_98_26 bit_98_26 bitb_98_26 word98_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_26 q_99_26 qb_99_26 bit_99_26 bitb_99_26 word99_26 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_27 q_0_27 qb_0_27 bit_0_27 bitb_0_27 word0_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_27 q_1_27 qb_1_27 bit_1_27 bitb_1_27 word1_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_27 q_2_27 qb_2_27 bit_2_27 bitb_2_27 word2_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_27 q_3_27 qb_3_27 bit_3_27 bitb_3_27 word3_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_27 q_4_27 qb_4_27 bit_4_27 bitb_4_27 word4_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_27 q_5_27 qb_5_27 bit_5_27 bitb_5_27 word5_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_27 q_6_27 qb_6_27 bit_6_27 bitb_6_27 word6_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_27 q_7_27 qb_7_27 bit_7_27 bitb_7_27 word7_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_27 q_8_27 qb_8_27 bit_8_27 bitb_8_27 word8_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_27 q_9_27 qb_9_27 bit_9_27 bitb_9_27 word9_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_27 q_10_27 qb_10_27 bit_10_27 bitb_10_27 word10_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_27 q_11_27 qb_11_27 bit_11_27 bitb_11_27 word11_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_27 q_12_27 qb_12_27 bit_12_27 bitb_12_27 word12_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_27 q_13_27 qb_13_27 bit_13_27 bitb_13_27 word13_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_27 q_14_27 qb_14_27 bit_14_27 bitb_14_27 word14_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_27 q_15_27 qb_15_27 bit_15_27 bitb_15_27 word15_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_27 q_16_27 qb_16_27 bit_16_27 bitb_16_27 word16_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_27 q_17_27 qb_17_27 bit_17_27 bitb_17_27 word17_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_27 q_18_27 qb_18_27 bit_18_27 bitb_18_27 word18_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_27 q_19_27 qb_19_27 bit_19_27 bitb_19_27 word19_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_27 q_20_27 qb_20_27 bit_20_27 bitb_20_27 word20_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_27 q_21_27 qb_21_27 bit_21_27 bitb_21_27 word21_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_27 q_22_27 qb_22_27 bit_22_27 bitb_22_27 word22_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_27 q_23_27 qb_23_27 bit_23_27 bitb_23_27 word23_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_27 q_24_27 qb_24_27 bit_24_27 bitb_24_27 word24_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_27 q_25_27 qb_25_27 bit_25_27 bitb_25_27 word25_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_27 q_26_27 qb_26_27 bit_26_27 bitb_26_27 word26_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_27 q_27_27 qb_27_27 bit_27_27 bitb_27_27 word27_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_27 q_28_27 qb_28_27 bit_28_27 bitb_28_27 word28_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_27 q_29_27 qb_29_27 bit_29_27 bitb_29_27 word29_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_27 q_30_27 qb_30_27 bit_30_27 bitb_30_27 word30_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_27 q_31_27 qb_31_27 bit_31_27 bitb_31_27 word31_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_27 q_32_27 qb_32_27 bit_32_27 bitb_32_27 word32_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_27 q_33_27 qb_33_27 bit_33_27 bitb_33_27 word33_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_27 q_34_27 qb_34_27 bit_34_27 bitb_34_27 word34_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_27 q_35_27 qb_35_27 bit_35_27 bitb_35_27 word35_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_27 q_36_27 qb_36_27 bit_36_27 bitb_36_27 word36_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_27 q_37_27 qb_37_27 bit_37_27 bitb_37_27 word37_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_27 q_38_27 qb_38_27 bit_38_27 bitb_38_27 word38_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_27 q_39_27 qb_39_27 bit_39_27 bitb_39_27 word39_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_27 q_40_27 qb_40_27 bit_40_27 bitb_40_27 word40_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_27 q_41_27 qb_41_27 bit_41_27 bitb_41_27 word41_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_27 q_42_27 qb_42_27 bit_42_27 bitb_42_27 word42_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_27 q_43_27 qb_43_27 bit_43_27 bitb_43_27 word43_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_27 q_44_27 qb_44_27 bit_44_27 bitb_44_27 word44_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_27 q_45_27 qb_45_27 bit_45_27 bitb_45_27 word45_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_27 q_46_27 qb_46_27 bit_46_27 bitb_46_27 word46_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_27 q_47_27 qb_47_27 bit_47_27 bitb_47_27 word47_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_27 q_48_27 qb_48_27 bit_48_27 bitb_48_27 word48_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_27 q_49_27 qb_49_27 bit_49_27 bitb_49_27 word49_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_27 q_50_27 qb_50_27 bit_50_27 bitb_50_27 word50_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_27 q_51_27 qb_51_27 bit_51_27 bitb_51_27 word51_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_27 q_52_27 qb_52_27 bit_52_27 bitb_52_27 word52_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_27 q_53_27 qb_53_27 bit_53_27 bitb_53_27 word53_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_27 q_54_27 qb_54_27 bit_54_27 bitb_54_27 word54_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_27 q_55_27 qb_55_27 bit_55_27 bitb_55_27 word55_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_27 q_56_27 qb_56_27 bit_56_27 bitb_56_27 word56_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_27 q_57_27 qb_57_27 bit_57_27 bitb_57_27 word57_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_27 q_58_27 qb_58_27 bit_58_27 bitb_58_27 word58_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_27 q_59_27 qb_59_27 bit_59_27 bitb_59_27 word59_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_27 q_60_27 qb_60_27 bit_60_27 bitb_60_27 word60_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_27 q_61_27 qb_61_27 bit_61_27 bitb_61_27 word61_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_27 q_62_27 qb_62_27 bit_62_27 bitb_62_27 word62_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_27 q_63_27 qb_63_27 bit_63_27 bitb_63_27 word63_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_27 q_64_27 qb_64_27 bit_64_27 bitb_64_27 word64_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_27 q_65_27 qb_65_27 bit_65_27 bitb_65_27 word65_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_27 q_66_27 qb_66_27 bit_66_27 bitb_66_27 word66_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_27 q_67_27 qb_67_27 bit_67_27 bitb_67_27 word67_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_27 q_68_27 qb_68_27 bit_68_27 bitb_68_27 word68_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_27 q_69_27 qb_69_27 bit_69_27 bitb_69_27 word69_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_27 q_70_27 qb_70_27 bit_70_27 bitb_70_27 word70_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_27 q_71_27 qb_71_27 bit_71_27 bitb_71_27 word71_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_27 q_72_27 qb_72_27 bit_72_27 bitb_72_27 word72_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_27 q_73_27 qb_73_27 bit_73_27 bitb_73_27 word73_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_27 q_74_27 qb_74_27 bit_74_27 bitb_74_27 word74_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_27 q_75_27 qb_75_27 bit_75_27 bitb_75_27 word75_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_27 q_76_27 qb_76_27 bit_76_27 bitb_76_27 word76_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_27 q_77_27 qb_77_27 bit_77_27 bitb_77_27 word77_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_27 q_78_27 qb_78_27 bit_78_27 bitb_78_27 word78_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_27 q_79_27 qb_79_27 bit_79_27 bitb_79_27 word79_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_27 q_80_27 qb_80_27 bit_80_27 bitb_80_27 word80_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_27 q_81_27 qb_81_27 bit_81_27 bitb_81_27 word81_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_27 q_82_27 qb_82_27 bit_82_27 bitb_82_27 word82_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_27 q_83_27 qb_83_27 bit_83_27 bitb_83_27 word83_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_27 q_84_27 qb_84_27 bit_84_27 bitb_84_27 word84_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_27 q_85_27 qb_85_27 bit_85_27 bitb_85_27 word85_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_27 q_86_27 qb_86_27 bit_86_27 bitb_86_27 word86_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_27 q_87_27 qb_87_27 bit_87_27 bitb_87_27 word87_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_27 q_88_27 qb_88_27 bit_88_27 bitb_88_27 word88_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_27 q_89_27 qb_89_27 bit_89_27 bitb_89_27 word89_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_27 q_90_27 qb_90_27 bit_90_27 bitb_90_27 word90_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_27 q_91_27 qb_91_27 bit_91_27 bitb_91_27 word91_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_27 q_92_27 qb_92_27 bit_92_27 bitb_92_27 word92_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_27 q_93_27 qb_93_27 bit_93_27 bitb_93_27 word93_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_27 q_94_27 qb_94_27 bit_94_27 bitb_94_27 word94_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_27 q_95_27 qb_95_27 bit_95_27 bitb_95_27 word95_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_27 q_96_27 qb_96_27 bit_96_27 bitb_96_27 word96_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_27 q_97_27 qb_97_27 bit_97_27 bitb_97_27 word97_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_27 q_98_27 qb_98_27 bit_98_27 bitb_98_27 word98_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_27 q_99_27 qb_99_27 bit_99_27 bitb_99_27 word99_27 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_28 q_0_28 qb_0_28 bit_0_28 bitb_0_28 word0_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_28 q_1_28 qb_1_28 bit_1_28 bitb_1_28 word1_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_28 q_2_28 qb_2_28 bit_2_28 bitb_2_28 word2_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_28 q_3_28 qb_3_28 bit_3_28 bitb_3_28 word3_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_28 q_4_28 qb_4_28 bit_4_28 bitb_4_28 word4_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_28 q_5_28 qb_5_28 bit_5_28 bitb_5_28 word5_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_28 q_6_28 qb_6_28 bit_6_28 bitb_6_28 word6_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_28 q_7_28 qb_7_28 bit_7_28 bitb_7_28 word7_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_28 q_8_28 qb_8_28 bit_8_28 bitb_8_28 word8_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_28 q_9_28 qb_9_28 bit_9_28 bitb_9_28 word9_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_28 q_10_28 qb_10_28 bit_10_28 bitb_10_28 word10_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_28 q_11_28 qb_11_28 bit_11_28 bitb_11_28 word11_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_28 q_12_28 qb_12_28 bit_12_28 bitb_12_28 word12_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_28 q_13_28 qb_13_28 bit_13_28 bitb_13_28 word13_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_28 q_14_28 qb_14_28 bit_14_28 bitb_14_28 word14_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_28 q_15_28 qb_15_28 bit_15_28 bitb_15_28 word15_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_28 q_16_28 qb_16_28 bit_16_28 bitb_16_28 word16_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_28 q_17_28 qb_17_28 bit_17_28 bitb_17_28 word17_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_28 q_18_28 qb_18_28 bit_18_28 bitb_18_28 word18_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_28 q_19_28 qb_19_28 bit_19_28 bitb_19_28 word19_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_28 q_20_28 qb_20_28 bit_20_28 bitb_20_28 word20_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_28 q_21_28 qb_21_28 bit_21_28 bitb_21_28 word21_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_28 q_22_28 qb_22_28 bit_22_28 bitb_22_28 word22_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_28 q_23_28 qb_23_28 bit_23_28 bitb_23_28 word23_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_28 q_24_28 qb_24_28 bit_24_28 bitb_24_28 word24_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_28 q_25_28 qb_25_28 bit_25_28 bitb_25_28 word25_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_28 q_26_28 qb_26_28 bit_26_28 bitb_26_28 word26_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_28 q_27_28 qb_27_28 bit_27_28 bitb_27_28 word27_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_28 q_28_28 qb_28_28 bit_28_28 bitb_28_28 word28_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_28 q_29_28 qb_29_28 bit_29_28 bitb_29_28 word29_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_28 q_30_28 qb_30_28 bit_30_28 bitb_30_28 word30_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_28 q_31_28 qb_31_28 bit_31_28 bitb_31_28 word31_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_28 q_32_28 qb_32_28 bit_32_28 bitb_32_28 word32_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_28 q_33_28 qb_33_28 bit_33_28 bitb_33_28 word33_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_28 q_34_28 qb_34_28 bit_34_28 bitb_34_28 word34_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_28 q_35_28 qb_35_28 bit_35_28 bitb_35_28 word35_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_28 q_36_28 qb_36_28 bit_36_28 bitb_36_28 word36_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_28 q_37_28 qb_37_28 bit_37_28 bitb_37_28 word37_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_28 q_38_28 qb_38_28 bit_38_28 bitb_38_28 word38_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_28 q_39_28 qb_39_28 bit_39_28 bitb_39_28 word39_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_28 q_40_28 qb_40_28 bit_40_28 bitb_40_28 word40_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_28 q_41_28 qb_41_28 bit_41_28 bitb_41_28 word41_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_28 q_42_28 qb_42_28 bit_42_28 bitb_42_28 word42_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_28 q_43_28 qb_43_28 bit_43_28 bitb_43_28 word43_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_28 q_44_28 qb_44_28 bit_44_28 bitb_44_28 word44_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_28 q_45_28 qb_45_28 bit_45_28 bitb_45_28 word45_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_28 q_46_28 qb_46_28 bit_46_28 bitb_46_28 word46_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_28 q_47_28 qb_47_28 bit_47_28 bitb_47_28 word47_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_28 q_48_28 qb_48_28 bit_48_28 bitb_48_28 word48_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_28 q_49_28 qb_49_28 bit_49_28 bitb_49_28 word49_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_28 q_50_28 qb_50_28 bit_50_28 bitb_50_28 word50_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_28 q_51_28 qb_51_28 bit_51_28 bitb_51_28 word51_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_28 q_52_28 qb_52_28 bit_52_28 bitb_52_28 word52_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_28 q_53_28 qb_53_28 bit_53_28 bitb_53_28 word53_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_28 q_54_28 qb_54_28 bit_54_28 bitb_54_28 word54_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_28 q_55_28 qb_55_28 bit_55_28 bitb_55_28 word55_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_28 q_56_28 qb_56_28 bit_56_28 bitb_56_28 word56_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_28 q_57_28 qb_57_28 bit_57_28 bitb_57_28 word57_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_28 q_58_28 qb_58_28 bit_58_28 bitb_58_28 word58_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_28 q_59_28 qb_59_28 bit_59_28 bitb_59_28 word59_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_28 q_60_28 qb_60_28 bit_60_28 bitb_60_28 word60_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_28 q_61_28 qb_61_28 bit_61_28 bitb_61_28 word61_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_28 q_62_28 qb_62_28 bit_62_28 bitb_62_28 word62_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_28 q_63_28 qb_63_28 bit_63_28 bitb_63_28 word63_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_28 q_64_28 qb_64_28 bit_64_28 bitb_64_28 word64_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_28 q_65_28 qb_65_28 bit_65_28 bitb_65_28 word65_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_28 q_66_28 qb_66_28 bit_66_28 bitb_66_28 word66_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_28 q_67_28 qb_67_28 bit_67_28 bitb_67_28 word67_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_28 q_68_28 qb_68_28 bit_68_28 bitb_68_28 word68_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_28 q_69_28 qb_69_28 bit_69_28 bitb_69_28 word69_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_28 q_70_28 qb_70_28 bit_70_28 bitb_70_28 word70_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_28 q_71_28 qb_71_28 bit_71_28 bitb_71_28 word71_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_28 q_72_28 qb_72_28 bit_72_28 bitb_72_28 word72_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_28 q_73_28 qb_73_28 bit_73_28 bitb_73_28 word73_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_28 q_74_28 qb_74_28 bit_74_28 bitb_74_28 word74_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_28 q_75_28 qb_75_28 bit_75_28 bitb_75_28 word75_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_28 q_76_28 qb_76_28 bit_76_28 bitb_76_28 word76_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_28 q_77_28 qb_77_28 bit_77_28 bitb_77_28 word77_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_28 q_78_28 qb_78_28 bit_78_28 bitb_78_28 word78_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_28 q_79_28 qb_79_28 bit_79_28 bitb_79_28 word79_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_28 q_80_28 qb_80_28 bit_80_28 bitb_80_28 word80_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_28 q_81_28 qb_81_28 bit_81_28 bitb_81_28 word81_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_28 q_82_28 qb_82_28 bit_82_28 bitb_82_28 word82_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_28 q_83_28 qb_83_28 bit_83_28 bitb_83_28 word83_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_28 q_84_28 qb_84_28 bit_84_28 bitb_84_28 word84_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_28 q_85_28 qb_85_28 bit_85_28 bitb_85_28 word85_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_28 q_86_28 qb_86_28 bit_86_28 bitb_86_28 word86_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_28 q_87_28 qb_87_28 bit_87_28 bitb_87_28 word87_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_28 q_88_28 qb_88_28 bit_88_28 bitb_88_28 word88_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_28 q_89_28 qb_89_28 bit_89_28 bitb_89_28 word89_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_28 q_90_28 qb_90_28 bit_90_28 bitb_90_28 word90_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_28 q_91_28 qb_91_28 bit_91_28 bitb_91_28 word91_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_28 q_92_28 qb_92_28 bit_92_28 bitb_92_28 word92_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_28 q_93_28 qb_93_28 bit_93_28 bitb_93_28 word93_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_28 q_94_28 qb_94_28 bit_94_28 bitb_94_28 word94_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_28 q_95_28 qb_95_28 bit_95_28 bitb_95_28 word95_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_28 q_96_28 qb_96_28 bit_96_28 bitb_96_28 word96_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_28 q_97_28 qb_97_28 bit_97_28 bitb_97_28 word97_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_28 q_98_28 qb_98_28 bit_98_28 bitb_98_28 word98_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_28 q_99_28 qb_99_28 bit_99_28 bitb_99_28 word99_28 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_29 q_0_29 qb_0_29 bit_0_29 bitb_0_29 word0_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_29 q_1_29 qb_1_29 bit_1_29 bitb_1_29 word1_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_29 q_2_29 qb_2_29 bit_2_29 bitb_2_29 word2_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_29 q_3_29 qb_3_29 bit_3_29 bitb_3_29 word3_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_29 q_4_29 qb_4_29 bit_4_29 bitb_4_29 word4_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_29 q_5_29 qb_5_29 bit_5_29 bitb_5_29 word5_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_29 q_6_29 qb_6_29 bit_6_29 bitb_6_29 word6_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_29 q_7_29 qb_7_29 bit_7_29 bitb_7_29 word7_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_29 q_8_29 qb_8_29 bit_8_29 bitb_8_29 word8_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_29 q_9_29 qb_9_29 bit_9_29 bitb_9_29 word9_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_29 q_10_29 qb_10_29 bit_10_29 bitb_10_29 word10_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_29 q_11_29 qb_11_29 bit_11_29 bitb_11_29 word11_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_29 q_12_29 qb_12_29 bit_12_29 bitb_12_29 word12_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_29 q_13_29 qb_13_29 bit_13_29 bitb_13_29 word13_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_29 q_14_29 qb_14_29 bit_14_29 bitb_14_29 word14_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_29 q_15_29 qb_15_29 bit_15_29 bitb_15_29 word15_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_29 q_16_29 qb_16_29 bit_16_29 bitb_16_29 word16_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_29 q_17_29 qb_17_29 bit_17_29 bitb_17_29 word17_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_29 q_18_29 qb_18_29 bit_18_29 bitb_18_29 word18_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_29 q_19_29 qb_19_29 bit_19_29 bitb_19_29 word19_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_29 q_20_29 qb_20_29 bit_20_29 bitb_20_29 word20_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_29 q_21_29 qb_21_29 bit_21_29 bitb_21_29 word21_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_29 q_22_29 qb_22_29 bit_22_29 bitb_22_29 word22_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_29 q_23_29 qb_23_29 bit_23_29 bitb_23_29 word23_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_29 q_24_29 qb_24_29 bit_24_29 bitb_24_29 word24_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_29 q_25_29 qb_25_29 bit_25_29 bitb_25_29 word25_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_29 q_26_29 qb_26_29 bit_26_29 bitb_26_29 word26_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_29 q_27_29 qb_27_29 bit_27_29 bitb_27_29 word27_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_29 q_28_29 qb_28_29 bit_28_29 bitb_28_29 word28_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_29 q_29_29 qb_29_29 bit_29_29 bitb_29_29 word29_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_29 q_30_29 qb_30_29 bit_30_29 bitb_30_29 word30_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_29 q_31_29 qb_31_29 bit_31_29 bitb_31_29 word31_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_29 q_32_29 qb_32_29 bit_32_29 bitb_32_29 word32_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_29 q_33_29 qb_33_29 bit_33_29 bitb_33_29 word33_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_29 q_34_29 qb_34_29 bit_34_29 bitb_34_29 word34_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_29 q_35_29 qb_35_29 bit_35_29 bitb_35_29 word35_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_29 q_36_29 qb_36_29 bit_36_29 bitb_36_29 word36_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_29 q_37_29 qb_37_29 bit_37_29 bitb_37_29 word37_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_29 q_38_29 qb_38_29 bit_38_29 bitb_38_29 word38_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_29 q_39_29 qb_39_29 bit_39_29 bitb_39_29 word39_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_29 q_40_29 qb_40_29 bit_40_29 bitb_40_29 word40_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_29 q_41_29 qb_41_29 bit_41_29 bitb_41_29 word41_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_29 q_42_29 qb_42_29 bit_42_29 bitb_42_29 word42_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_29 q_43_29 qb_43_29 bit_43_29 bitb_43_29 word43_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_29 q_44_29 qb_44_29 bit_44_29 bitb_44_29 word44_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_29 q_45_29 qb_45_29 bit_45_29 bitb_45_29 word45_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_29 q_46_29 qb_46_29 bit_46_29 bitb_46_29 word46_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_29 q_47_29 qb_47_29 bit_47_29 bitb_47_29 word47_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_29 q_48_29 qb_48_29 bit_48_29 bitb_48_29 word48_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_29 q_49_29 qb_49_29 bit_49_29 bitb_49_29 word49_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_29 q_50_29 qb_50_29 bit_50_29 bitb_50_29 word50_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_29 q_51_29 qb_51_29 bit_51_29 bitb_51_29 word51_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_29 q_52_29 qb_52_29 bit_52_29 bitb_52_29 word52_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_29 q_53_29 qb_53_29 bit_53_29 bitb_53_29 word53_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_29 q_54_29 qb_54_29 bit_54_29 bitb_54_29 word54_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_29 q_55_29 qb_55_29 bit_55_29 bitb_55_29 word55_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_29 q_56_29 qb_56_29 bit_56_29 bitb_56_29 word56_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_29 q_57_29 qb_57_29 bit_57_29 bitb_57_29 word57_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_29 q_58_29 qb_58_29 bit_58_29 bitb_58_29 word58_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_29 q_59_29 qb_59_29 bit_59_29 bitb_59_29 word59_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_29 q_60_29 qb_60_29 bit_60_29 bitb_60_29 word60_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_29 q_61_29 qb_61_29 bit_61_29 bitb_61_29 word61_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_29 q_62_29 qb_62_29 bit_62_29 bitb_62_29 word62_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_29 q_63_29 qb_63_29 bit_63_29 bitb_63_29 word63_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_29 q_64_29 qb_64_29 bit_64_29 bitb_64_29 word64_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_29 q_65_29 qb_65_29 bit_65_29 bitb_65_29 word65_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_29 q_66_29 qb_66_29 bit_66_29 bitb_66_29 word66_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_29 q_67_29 qb_67_29 bit_67_29 bitb_67_29 word67_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_29 q_68_29 qb_68_29 bit_68_29 bitb_68_29 word68_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_29 q_69_29 qb_69_29 bit_69_29 bitb_69_29 word69_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_29 q_70_29 qb_70_29 bit_70_29 bitb_70_29 word70_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_29 q_71_29 qb_71_29 bit_71_29 bitb_71_29 word71_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_29 q_72_29 qb_72_29 bit_72_29 bitb_72_29 word72_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_29 q_73_29 qb_73_29 bit_73_29 bitb_73_29 word73_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_29 q_74_29 qb_74_29 bit_74_29 bitb_74_29 word74_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_29 q_75_29 qb_75_29 bit_75_29 bitb_75_29 word75_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_29 q_76_29 qb_76_29 bit_76_29 bitb_76_29 word76_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_29 q_77_29 qb_77_29 bit_77_29 bitb_77_29 word77_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_29 q_78_29 qb_78_29 bit_78_29 bitb_78_29 word78_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_29 q_79_29 qb_79_29 bit_79_29 bitb_79_29 word79_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_29 q_80_29 qb_80_29 bit_80_29 bitb_80_29 word80_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_29 q_81_29 qb_81_29 bit_81_29 bitb_81_29 word81_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_29 q_82_29 qb_82_29 bit_82_29 bitb_82_29 word82_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_29 q_83_29 qb_83_29 bit_83_29 bitb_83_29 word83_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_29 q_84_29 qb_84_29 bit_84_29 bitb_84_29 word84_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_29 q_85_29 qb_85_29 bit_85_29 bitb_85_29 word85_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_29 q_86_29 qb_86_29 bit_86_29 bitb_86_29 word86_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_29 q_87_29 qb_87_29 bit_87_29 bitb_87_29 word87_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_29 q_88_29 qb_88_29 bit_88_29 bitb_88_29 word88_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_29 q_89_29 qb_89_29 bit_89_29 bitb_89_29 word89_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_29 q_90_29 qb_90_29 bit_90_29 bitb_90_29 word90_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_29 q_91_29 qb_91_29 bit_91_29 bitb_91_29 word91_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_29 q_92_29 qb_92_29 bit_92_29 bitb_92_29 word92_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_29 q_93_29 qb_93_29 bit_93_29 bitb_93_29 word93_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_29 q_94_29 qb_94_29 bit_94_29 bitb_94_29 word94_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_29 q_95_29 qb_95_29 bit_95_29 bitb_95_29 word95_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_29 q_96_29 qb_96_29 bit_96_29 bitb_96_29 word96_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_29 q_97_29 qb_97_29 bit_97_29 bitb_97_29 word97_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_29 q_98_29 qb_98_29 bit_98_29 bitb_98_29 word98_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_29 q_99_29 qb_99_29 bit_99_29 bitb_99_29 word99_29 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_30 q_0_30 qb_0_30 bit_0_30 bitb_0_30 word0_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_30 q_1_30 qb_1_30 bit_1_30 bitb_1_30 word1_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_30 q_2_30 qb_2_30 bit_2_30 bitb_2_30 word2_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_30 q_3_30 qb_3_30 bit_3_30 bitb_3_30 word3_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_30 q_4_30 qb_4_30 bit_4_30 bitb_4_30 word4_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_30 q_5_30 qb_5_30 bit_5_30 bitb_5_30 word5_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_30 q_6_30 qb_6_30 bit_6_30 bitb_6_30 word6_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_30 q_7_30 qb_7_30 bit_7_30 bitb_7_30 word7_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_30 q_8_30 qb_8_30 bit_8_30 bitb_8_30 word8_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_30 q_9_30 qb_9_30 bit_9_30 bitb_9_30 word9_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_30 q_10_30 qb_10_30 bit_10_30 bitb_10_30 word10_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_30 q_11_30 qb_11_30 bit_11_30 bitb_11_30 word11_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_30 q_12_30 qb_12_30 bit_12_30 bitb_12_30 word12_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_30 q_13_30 qb_13_30 bit_13_30 bitb_13_30 word13_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_30 q_14_30 qb_14_30 bit_14_30 bitb_14_30 word14_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_30 q_15_30 qb_15_30 bit_15_30 bitb_15_30 word15_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_30 q_16_30 qb_16_30 bit_16_30 bitb_16_30 word16_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_30 q_17_30 qb_17_30 bit_17_30 bitb_17_30 word17_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_30 q_18_30 qb_18_30 bit_18_30 bitb_18_30 word18_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_30 q_19_30 qb_19_30 bit_19_30 bitb_19_30 word19_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_30 q_20_30 qb_20_30 bit_20_30 bitb_20_30 word20_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_30 q_21_30 qb_21_30 bit_21_30 bitb_21_30 word21_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_30 q_22_30 qb_22_30 bit_22_30 bitb_22_30 word22_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_30 q_23_30 qb_23_30 bit_23_30 bitb_23_30 word23_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_30 q_24_30 qb_24_30 bit_24_30 bitb_24_30 word24_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_30 q_25_30 qb_25_30 bit_25_30 bitb_25_30 word25_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_30 q_26_30 qb_26_30 bit_26_30 bitb_26_30 word26_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_30 q_27_30 qb_27_30 bit_27_30 bitb_27_30 word27_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_30 q_28_30 qb_28_30 bit_28_30 bitb_28_30 word28_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_30 q_29_30 qb_29_30 bit_29_30 bitb_29_30 word29_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_30 q_30_30 qb_30_30 bit_30_30 bitb_30_30 word30_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_30 q_31_30 qb_31_30 bit_31_30 bitb_31_30 word31_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_30 q_32_30 qb_32_30 bit_32_30 bitb_32_30 word32_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_30 q_33_30 qb_33_30 bit_33_30 bitb_33_30 word33_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_30 q_34_30 qb_34_30 bit_34_30 bitb_34_30 word34_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_30 q_35_30 qb_35_30 bit_35_30 bitb_35_30 word35_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_30 q_36_30 qb_36_30 bit_36_30 bitb_36_30 word36_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_30 q_37_30 qb_37_30 bit_37_30 bitb_37_30 word37_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_30 q_38_30 qb_38_30 bit_38_30 bitb_38_30 word38_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_30 q_39_30 qb_39_30 bit_39_30 bitb_39_30 word39_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_30 q_40_30 qb_40_30 bit_40_30 bitb_40_30 word40_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_30 q_41_30 qb_41_30 bit_41_30 bitb_41_30 word41_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_30 q_42_30 qb_42_30 bit_42_30 bitb_42_30 word42_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_30 q_43_30 qb_43_30 bit_43_30 bitb_43_30 word43_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_30 q_44_30 qb_44_30 bit_44_30 bitb_44_30 word44_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_30 q_45_30 qb_45_30 bit_45_30 bitb_45_30 word45_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_30 q_46_30 qb_46_30 bit_46_30 bitb_46_30 word46_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_30 q_47_30 qb_47_30 bit_47_30 bitb_47_30 word47_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_30 q_48_30 qb_48_30 bit_48_30 bitb_48_30 word48_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_30 q_49_30 qb_49_30 bit_49_30 bitb_49_30 word49_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_30 q_50_30 qb_50_30 bit_50_30 bitb_50_30 word50_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_30 q_51_30 qb_51_30 bit_51_30 bitb_51_30 word51_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_30 q_52_30 qb_52_30 bit_52_30 bitb_52_30 word52_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_30 q_53_30 qb_53_30 bit_53_30 bitb_53_30 word53_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_30 q_54_30 qb_54_30 bit_54_30 bitb_54_30 word54_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_30 q_55_30 qb_55_30 bit_55_30 bitb_55_30 word55_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_30 q_56_30 qb_56_30 bit_56_30 bitb_56_30 word56_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_30 q_57_30 qb_57_30 bit_57_30 bitb_57_30 word57_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_30 q_58_30 qb_58_30 bit_58_30 bitb_58_30 word58_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_30 q_59_30 qb_59_30 bit_59_30 bitb_59_30 word59_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_30 q_60_30 qb_60_30 bit_60_30 bitb_60_30 word60_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_30 q_61_30 qb_61_30 bit_61_30 bitb_61_30 word61_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_30 q_62_30 qb_62_30 bit_62_30 bitb_62_30 word62_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_30 q_63_30 qb_63_30 bit_63_30 bitb_63_30 word63_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_30 q_64_30 qb_64_30 bit_64_30 bitb_64_30 word64_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_30 q_65_30 qb_65_30 bit_65_30 bitb_65_30 word65_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_30 q_66_30 qb_66_30 bit_66_30 bitb_66_30 word66_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_30 q_67_30 qb_67_30 bit_67_30 bitb_67_30 word67_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_30 q_68_30 qb_68_30 bit_68_30 bitb_68_30 word68_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_30 q_69_30 qb_69_30 bit_69_30 bitb_69_30 word69_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_30 q_70_30 qb_70_30 bit_70_30 bitb_70_30 word70_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_30 q_71_30 qb_71_30 bit_71_30 bitb_71_30 word71_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_30 q_72_30 qb_72_30 bit_72_30 bitb_72_30 word72_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_30 q_73_30 qb_73_30 bit_73_30 bitb_73_30 word73_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_30 q_74_30 qb_74_30 bit_74_30 bitb_74_30 word74_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_30 q_75_30 qb_75_30 bit_75_30 bitb_75_30 word75_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_30 q_76_30 qb_76_30 bit_76_30 bitb_76_30 word76_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_30 q_77_30 qb_77_30 bit_77_30 bitb_77_30 word77_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_30 q_78_30 qb_78_30 bit_78_30 bitb_78_30 word78_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_30 q_79_30 qb_79_30 bit_79_30 bitb_79_30 word79_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_30 q_80_30 qb_80_30 bit_80_30 bitb_80_30 word80_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_30 q_81_30 qb_81_30 bit_81_30 bitb_81_30 word81_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_30 q_82_30 qb_82_30 bit_82_30 bitb_82_30 word82_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_30 q_83_30 qb_83_30 bit_83_30 bitb_83_30 word83_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_30 q_84_30 qb_84_30 bit_84_30 bitb_84_30 word84_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_30 q_85_30 qb_85_30 bit_85_30 bitb_85_30 word85_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_30 q_86_30 qb_86_30 bit_86_30 bitb_86_30 word86_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_30 q_87_30 qb_87_30 bit_87_30 bitb_87_30 word87_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_30 q_88_30 qb_88_30 bit_88_30 bitb_88_30 word88_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_30 q_89_30 qb_89_30 bit_89_30 bitb_89_30 word89_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_30 q_90_30 qb_90_30 bit_90_30 bitb_90_30 word90_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_30 q_91_30 qb_91_30 bit_91_30 bitb_91_30 word91_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_30 q_92_30 qb_92_30 bit_92_30 bitb_92_30 word92_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_30 q_93_30 qb_93_30 bit_93_30 bitb_93_30 word93_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_30 q_94_30 qb_94_30 bit_94_30 bitb_94_30 word94_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_30 q_95_30 qb_95_30 bit_95_30 bitb_95_30 word95_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_30 q_96_30 qb_96_30 bit_96_30 bitb_96_30 word96_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_30 q_97_30 qb_97_30 bit_97_30 bitb_97_30 word97_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_30 q_98_30 qb_98_30 bit_98_30 bitb_98_30 word98_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_30 q_99_30 qb_99_30 bit_99_30 bitb_99_30 word99_30 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_31 q_0_31 qb_0_31 bit_0_31 bitb_0_31 word0_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_31 q_1_31 qb_1_31 bit_1_31 bitb_1_31 word1_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_31 q_2_31 qb_2_31 bit_2_31 bitb_2_31 word2_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_31 q_3_31 qb_3_31 bit_3_31 bitb_3_31 word3_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_31 q_4_31 qb_4_31 bit_4_31 bitb_4_31 word4_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_31 q_5_31 qb_5_31 bit_5_31 bitb_5_31 word5_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_31 q_6_31 qb_6_31 bit_6_31 bitb_6_31 word6_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_31 q_7_31 qb_7_31 bit_7_31 bitb_7_31 word7_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_31 q_8_31 qb_8_31 bit_8_31 bitb_8_31 word8_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_31 q_9_31 qb_9_31 bit_9_31 bitb_9_31 word9_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_31 q_10_31 qb_10_31 bit_10_31 bitb_10_31 word10_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_31 q_11_31 qb_11_31 bit_11_31 bitb_11_31 word11_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_31 q_12_31 qb_12_31 bit_12_31 bitb_12_31 word12_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_31 q_13_31 qb_13_31 bit_13_31 bitb_13_31 word13_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_31 q_14_31 qb_14_31 bit_14_31 bitb_14_31 word14_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_31 q_15_31 qb_15_31 bit_15_31 bitb_15_31 word15_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_31 q_16_31 qb_16_31 bit_16_31 bitb_16_31 word16_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_31 q_17_31 qb_17_31 bit_17_31 bitb_17_31 word17_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_31 q_18_31 qb_18_31 bit_18_31 bitb_18_31 word18_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_31 q_19_31 qb_19_31 bit_19_31 bitb_19_31 word19_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_31 q_20_31 qb_20_31 bit_20_31 bitb_20_31 word20_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_31 q_21_31 qb_21_31 bit_21_31 bitb_21_31 word21_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_31 q_22_31 qb_22_31 bit_22_31 bitb_22_31 word22_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_31 q_23_31 qb_23_31 bit_23_31 bitb_23_31 word23_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_31 q_24_31 qb_24_31 bit_24_31 bitb_24_31 word24_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_31 q_25_31 qb_25_31 bit_25_31 bitb_25_31 word25_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_31 q_26_31 qb_26_31 bit_26_31 bitb_26_31 word26_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_31 q_27_31 qb_27_31 bit_27_31 bitb_27_31 word27_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_31 q_28_31 qb_28_31 bit_28_31 bitb_28_31 word28_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_31 q_29_31 qb_29_31 bit_29_31 bitb_29_31 word29_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_31 q_30_31 qb_30_31 bit_30_31 bitb_30_31 word30_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_31 q_31_31 qb_31_31 bit_31_31 bitb_31_31 word31_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_31 q_32_31 qb_32_31 bit_32_31 bitb_32_31 word32_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_31 q_33_31 qb_33_31 bit_33_31 bitb_33_31 word33_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_31 q_34_31 qb_34_31 bit_34_31 bitb_34_31 word34_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_31 q_35_31 qb_35_31 bit_35_31 bitb_35_31 word35_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_31 q_36_31 qb_36_31 bit_36_31 bitb_36_31 word36_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_31 q_37_31 qb_37_31 bit_37_31 bitb_37_31 word37_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_31 q_38_31 qb_38_31 bit_38_31 bitb_38_31 word38_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_31 q_39_31 qb_39_31 bit_39_31 bitb_39_31 word39_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_31 q_40_31 qb_40_31 bit_40_31 bitb_40_31 word40_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_31 q_41_31 qb_41_31 bit_41_31 bitb_41_31 word41_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_31 q_42_31 qb_42_31 bit_42_31 bitb_42_31 word42_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_31 q_43_31 qb_43_31 bit_43_31 bitb_43_31 word43_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_31 q_44_31 qb_44_31 bit_44_31 bitb_44_31 word44_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_31 q_45_31 qb_45_31 bit_45_31 bitb_45_31 word45_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_31 q_46_31 qb_46_31 bit_46_31 bitb_46_31 word46_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_31 q_47_31 qb_47_31 bit_47_31 bitb_47_31 word47_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_31 q_48_31 qb_48_31 bit_48_31 bitb_48_31 word48_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_31 q_49_31 qb_49_31 bit_49_31 bitb_49_31 word49_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_31 q_50_31 qb_50_31 bit_50_31 bitb_50_31 word50_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_31 q_51_31 qb_51_31 bit_51_31 bitb_51_31 word51_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_31 q_52_31 qb_52_31 bit_52_31 bitb_52_31 word52_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_31 q_53_31 qb_53_31 bit_53_31 bitb_53_31 word53_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_31 q_54_31 qb_54_31 bit_54_31 bitb_54_31 word54_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_31 q_55_31 qb_55_31 bit_55_31 bitb_55_31 word55_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_31 q_56_31 qb_56_31 bit_56_31 bitb_56_31 word56_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_31 q_57_31 qb_57_31 bit_57_31 bitb_57_31 word57_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_31 q_58_31 qb_58_31 bit_58_31 bitb_58_31 word58_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_31 q_59_31 qb_59_31 bit_59_31 bitb_59_31 word59_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_31 q_60_31 qb_60_31 bit_60_31 bitb_60_31 word60_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_31 q_61_31 qb_61_31 bit_61_31 bitb_61_31 word61_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_31 q_62_31 qb_62_31 bit_62_31 bitb_62_31 word62_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_31 q_63_31 qb_63_31 bit_63_31 bitb_63_31 word63_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_31 q_64_31 qb_64_31 bit_64_31 bitb_64_31 word64_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_31 q_65_31 qb_65_31 bit_65_31 bitb_65_31 word65_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_31 q_66_31 qb_66_31 bit_66_31 bitb_66_31 word66_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_31 q_67_31 qb_67_31 bit_67_31 bitb_67_31 word67_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_31 q_68_31 qb_68_31 bit_68_31 bitb_68_31 word68_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_31 q_69_31 qb_69_31 bit_69_31 bitb_69_31 word69_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_31 q_70_31 qb_70_31 bit_70_31 bitb_70_31 word70_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_31 q_71_31 qb_71_31 bit_71_31 bitb_71_31 word71_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_31 q_72_31 qb_72_31 bit_72_31 bitb_72_31 word72_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_31 q_73_31 qb_73_31 bit_73_31 bitb_73_31 word73_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_31 q_74_31 qb_74_31 bit_74_31 bitb_74_31 word74_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_31 q_75_31 qb_75_31 bit_75_31 bitb_75_31 word75_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_31 q_76_31 qb_76_31 bit_76_31 bitb_76_31 word76_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_31 q_77_31 qb_77_31 bit_77_31 bitb_77_31 word77_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_31 q_78_31 qb_78_31 bit_78_31 bitb_78_31 word78_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_31 q_79_31 qb_79_31 bit_79_31 bitb_79_31 word79_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_31 q_80_31 qb_80_31 bit_80_31 bitb_80_31 word80_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_31 q_81_31 qb_81_31 bit_81_31 bitb_81_31 word81_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_31 q_82_31 qb_82_31 bit_82_31 bitb_82_31 word82_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_31 q_83_31 qb_83_31 bit_83_31 bitb_83_31 word83_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_31 q_84_31 qb_84_31 bit_84_31 bitb_84_31 word84_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_31 q_85_31 qb_85_31 bit_85_31 bitb_85_31 word85_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_31 q_86_31 qb_86_31 bit_86_31 bitb_86_31 word86_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_31 q_87_31 qb_87_31 bit_87_31 bitb_87_31 word87_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_31 q_88_31 qb_88_31 bit_88_31 bitb_88_31 word88_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_31 q_89_31 qb_89_31 bit_89_31 bitb_89_31 word89_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_31 q_90_31 qb_90_31 bit_90_31 bitb_90_31 word90_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_31 q_91_31 qb_91_31 bit_91_31 bitb_91_31 word91_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_31 q_92_31 qb_92_31 bit_92_31 bitb_92_31 word92_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_31 q_93_31 qb_93_31 bit_93_31 bitb_93_31 word93_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_31 q_94_31 qb_94_31 bit_94_31 bitb_94_31 word94_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_31 q_95_31 qb_95_31 bit_95_31 bitb_95_31 word95_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_31 q_96_31 qb_96_31 bit_96_31 bitb_96_31 word96_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_31 q_97_31 qb_97_31 bit_97_31 bitb_97_31 word97_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_31 q_98_31 qb_98_31 bit_98_31 bitb_98_31 word98_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_31 q_99_31 qb_99_31 bit_99_31 bitb_99_31 word99_31 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_32 q_0_32 qb_0_32 bit_0_32 bitb_0_32 word0_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_32 q_1_32 qb_1_32 bit_1_32 bitb_1_32 word1_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_32 q_2_32 qb_2_32 bit_2_32 bitb_2_32 word2_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_32 q_3_32 qb_3_32 bit_3_32 bitb_3_32 word3_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_32 q_4_32 qb_4_32 bit_4_32 bitb_4_32 word4_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_32 q_5_32 qb_5_32 bit_5_32 bitb_5_32 word5_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_32 q_6_32 qb_6_32 bit_6_32 bitb_6_32 word6_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_32 q_7_32 qb_7_32 bit_7_32 bitb_7_32 word7_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_32 q_8_32 qb_8_32 bit_8_32 bitb_8_32 word8_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_32 q_9_32 qb_9_32 bit_9_32 bitb_9_32 word9_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_32 q_10_32 qb_10_32 bit_10_32 bitb_10_32 word10_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_32 q_11_32 qb_11_32 bit_11_32 bitb_11_32 word11_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_32 q_12_32 qb_12_32 bit_12_32 bitb_12_32 word12_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_32 q_13_32 qb_13_32 bit_13_32 bitb_13_32 word13_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_32 q_14_32 qb_14_32 bit_14_32 bitb_14_32 word14_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_32 q_15_32 qb_15_32 bit_15_32 bitb_15_32 word15_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_32 q_16_32 qb_16_32 bit_16_32 bitb_16_32 word16_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_32 q_17_32 qb_17_32 bit_17_32 bitb_17_32 word17_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_32 q_18_32 qb_18_32 bit_18_32 bitb_18_32 word18_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_32 q_19_32 qb_19_32 bit_19_32 bitb_19_32 word19_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_32 q_20_32 qb_20_32 bit_20_32 bitb_20_32 word20_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_32 q_21_32 qb_21_32 bit_21_32 bitb_21_32 word21_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_32 q_22_32 qb_22_32 bit_22_32 bitb_22_32 word22_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_32 q_23_32 qb_23_32 bit_23_32 bitb_23_32 word23_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_32 q_24_32 qb_24_32 bit_24_32 bitb_24_32 word24_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_32 q_25_32 qb_25_32 bit_25_32 bitb_25_32 word25_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_32 q_26_32 qb_26_32 bit_26_32 bitb_26_32 word26_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_32 q_27_32 qb_27_32 bit_27_32 bitb_27_32 word27_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_32 q_28_32 qb_28_32 bit_28_32 bitb_28_32 word28_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_32 q_29_32 qb_29_32 bit_29_32 bitb_29_32 word29_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_32 q_30_32 qb_30_32 bit_30_32 bitb_30_32 word30_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_32 q_31_32 qb_31_32 bit_31_32 bitb_31_32 word31_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_32 q_32_32 qb_32_32 bit_32_32 bitb_32_32 word32_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_32 q_33_32 qb_33_32 bit_33_32 bitb_33_32 word33_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_32 q_34_32 qb_34_32 bit_34_32 bitb_34_32 word34_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_32 q_35_32 qb_35_32 bit_35_32 bitb_35_32 word35_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_32 q_36_32 qb_36_32 bit_36_32 bitb_36_32 word36_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_32 q_37_32 qb_37_32 bit_37_32 bitb_37_32 word37_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_32 q_38_32 qb_38_32 bit_38_32 bitb_38_32 word38_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_32 q_39_32 qb_39_32 bit_39_32 bitb_39_32 word39_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_32 q_40_32 qb_40_32 bit_40_32 bitb_40_32 word40_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_32 q_41_32 qb_41_32 bit_41_32 bitb_41_32 word41_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_32 q_42_32 qb_42_32 bit_42_32 bitb_42_32 word42_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_32 q_43_32 qb_43_32 bit_43_32 bitb_43_32 word43_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_32 q_44_32 qb_44_32 bit_44_32 bitb_44_32 word44_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_32 q_45_32 qb_45_32 bit_45_32 bitb_45_32 word45_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_32 q_46_32 qb_46_32 bit_46_32 bitb_46_32 word46_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_32 q_47_32 qb_47_32 bit_47_32 bitb_47_32 word47_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_32 q_48_32 qb_48_32 bit_48_32 bitb_48_32 word48_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_32 q_49_32 qb_49_32 bit_49_32 bitb_49_32 word49_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_32 q_50_32 qb_50_32 bit_50_32 bitb_50_32 word50_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_32 q_51_32 qb_51_32 bit_51_32 bitb_51_32 word51_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_32 q_52_32 qb_52_32 bit_52_32 bitb_52_32 word52_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_32 q_53_32 qb_53_32 bit_53_32 bitb_53_32 word53_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_32 q_54_32 qb_54_32 bit_54_32 bitb_54_32 word54_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_32 q_55_32 qb_55_32 bit_55_32 bitb_55_32 word55_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_32 q_56_32 qb_56_32 bit_56_32 bitb_56_32 word56_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_32 q_57_32 qb_57_32 bit_57_32 bitb_57_32 word57_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_32 q_58_32 qb_58_32 bit_58_32 bitb_58_32 word58_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_32 q_59_32 qb_59_32 bit_59_32 bitb_59_32 word59_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_32 q_60_32 qb_60_32 bit_60_32 bitb_60_32 word60_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_32 q_61_32 qb_61_32 bit_61_32 bitb_61_32 word61_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_32 q_62_32 qb_62_32 bit_62_32 bitb_62_32 word62_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_32 q_63_32 qb_63_32 bit_63_32 bitb_63_32 word63_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_32 q_64_32 qb_64_32 bit_64_32 bitb_64_32 word64_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_32 q_65_32 qb_65_32 bit_65_32 bitb_65_32 word65_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_32 q_66_32 qb_66_32 bit_66_32 bitb_66_32 word66_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_32 q_67_32 qb_67_32 bit_67_32 bitb_67_32 word67_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_32 q_68_32 qb_68_32 bit_68_32 bitb_68_32 word68_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_32 q_69_32 qb_69_32 bit_69_32 bitb_69_32 word69_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_32 q_70_32 qb_70_32 bit_70_32 bitb_70_32 word70_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_32 q_71_32 qb_71_32 bit_71_32 bitb_71_32 word71_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_32 q_72_32 qb_72_32 bit_72_32 bitb_72_32 word72_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_32 q_73_32 qb_73_32 bit_73_32 bitb_73_32 word73_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_32 q_74_32 qb_74_32 bit_74_32 bitb_74_32 word74_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_32 q_75_32 qb_75_32 bit_75_32 bitb_75_32 word75_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_32 q_76_32 qb_76_32 bit_76_32 bitb_76_32 word76_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_32 q_77_32 qb_77_32 bit_77_32 bitb_77_32 word77_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_32 q_78_32 qb_78_32 bit_78_32 bitb_78_32 word78_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_32 q_79_32 qb_79_32 bit_79_32 bitb_79_32 word79_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_32 q_80_32 qb_80_32 bit_80_32 bitb_80_32 word80_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_32 q_81_32 qb_81_32 bit_81_32 bitb_81_32 word81_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_32 q_82_32 qb_82_32 bit_82_32 bitb_82_32 word82_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_32 q_83_32 qb_83_32 bit_83_32 bitb_83_32 word83_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_32 q_84_32 qb_84_32 bit_84_32 bitb_84_32 word84_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_32 q_85_32 qb_85_32 bit_85_32 bitb_85_32 word85_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_32 q_86_32 qb_86_32 bit_86_32 bitb_86_32 word86_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_32 q_87_32 qb_87_32 bit_87_32 bitb_87_32 word87_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_32 q_88_32 qb_88_32 bit_88_32 bitb_88_32 word88_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_32 q_89_32 qb_89_32 bit_89_32 bitb_89_32 word89_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_32 q_90_32 qb_90_32 bit_90_32 bitb_90_32 word90_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_32 q_91_32 qb_91_32 bit_91_32 bitb_91_32 word91_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_32 q_92_32 qb_92_32 bit_92_32 bitb_92_32 word92_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_32 q_93_32 qb_93_32 bit_93_32 bitb_93_32 word93_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_32 q_94_32 qb_94_32 bit_94_32 bitb_94_32 word94_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_32 q_95_32 qb_95_32 bit_95_32 bitb_95_32 word95_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_32 q_96_32 qb_96_32 bit_96_32 bitb_96_32 word96_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_32 q_97_32 qb_97_32 bit_97_32 bitb_97_32 word97_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_32 q_98_32 qb_98_32 bit_98_32 bitb_98_32 word98_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_32 q_99_32 qb_99_32 bit_99_32 bitb_99_32 word99_32 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_33 q_0_33 qb_0_33 bit_0_33 bitb_0_33 word0_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_33 q_1_33 qb_1_33 bit_1_33 bitb_1_33 word1_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_33 q_2_33 qb_2_33 bit_2_33 bitb_2_33 word2_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_33 q_3_33 qb_3_33 bit_3_33 bitb_3_33 word3_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_33 q_4_33 qb_4_33 bit_4_33 bitb_4_33 word4_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_33 q_5_33 qb_5_33 bit_5_33 bitb_5_33 word5_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_33 q_6_33 qb_6_33 bit_6_33 bitb_6_33 word6_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_33 q_7_33 qb_7_33 bit_7_33 bitb_7_33 word7_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_33 q_8_33 qb_8_33 bit_8_33 bitb_8_33 word8_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_33 q_9_33 qb_9_33 bit_9_33 bitb_9_33 word9_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_33 q_10_33 qb_10_33 bit_10_33 bitb_10_33 word10_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_33 q_11_33 qb_11_33 bit_11_33 bitb_11_33 word11_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_33 q_12_33 qb_12_33 bit_12_33 bitb_12_33 word12_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_33 q_13_33 qb_13_33 bit_13_33 bitb_13_33 word13_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_33 q_14_33 qb_14_33 bit_14_33 bitb_14_33 word14_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_33 q_15_33 qb_15_33 bit_15_33 bitb_15_33 word15_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_33 q_16_33 qb_16_33 bit_16_33 bitb_16_33 word16_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_33 q_17_33 qb_17_33 bit_17_33 bitb_17_33 word17_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_33 q_18_33 qb_18_33 bit_18_33 bitb_18_33 word18_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_33 q_19_33 qb_19_33 bit_19_33 bitb_19_33 word19_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_33 q_20_33 qb_20_33 bit_20_33 bitb_20_33 word20_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_33 q_21_33 qb_21_33 bit_21_33 bitb_21_33 word21_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_33 q_22_33 qb_22_33 bit_22_33 bitb_22_33 word22_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_33 q_23_33 qb_23_33 bit_23_33 bitb_23_33 word23_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_33 q_24_33 qb_24_33 bit_24_33 bitb_24_33 word24_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_33 q_25_33 qb_25_33 bit_25_33 bitb_25_33 word25_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_33 q_26_33 qb_26_33 bit_26_33 bitb_26_33 word26_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_33 q_27_33 qb_27_33 bit_27_33 bitb_27_33 word27_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_33 q_28_33 qb_28_33 bit_28_33 bitb_28_33 word28_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_33 q_29_33 qb_29_33 bit_29_33 bitb_29_33 word29_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_33 q_30_33 qb_30_33 bit_30_33 bitb_30_33 word30_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_33 q_31_33 qb_31_33 bit_31_33 bitb_31_33 word31_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_33 q_32_33 qb_32_33 bit_32_33 bitb_32_33 word32_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_33 q_33_33 qb_33_33 bit_33_33 bitb_33_33 word33_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_33 q_34_33 qb_34_33 bit_34_33 bitb_34_33 word34_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_33 q_35_33 qb_35_33 bit_35_33 bitb_35_33 word35_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_33 q_36_33 qb_36_33 bit_36_33 bitb_36_33 word36_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_33 q_37_33 qb_37_33 bit_37_33 bitb_37_33 word37_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_33 q_38_33 qb_38_33 bit_38_33 bitb_38_33 word38_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_33 q_39_33 qb_39_33 bit_39_33 bitb_39_33 word39_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_33 q_40_33 qb_40_33 bit_40_33 bitb_40_33 word40_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_33 q_41_33 qb_41_33 bit_41_33 bitb_41_33 word41_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_33 q_42_33 qb_42_33 bit_42_33 bitb_42_33 word42_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_33 q_43_33 qb_43_33 bit_43_33 bitb_43_33 word43_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_33 q_44_33 qb_44_33 bit_44_33 bitb_44_33 word44_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_33 q_45_33 qb_45_33 bit_45_33 bitb_45_33 word45_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_33 q_46_33 qb_46_33 bit_46_33 bitb_46_33 word46_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_33 q_47_33 qb_47_33 bit_47_33 bitb_47_33 word47_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_33 q_48_33 qb_48_33 bit_48_33 bitb_48_33 word48_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_33 q_49_33 qb_49_33 bit_49_33 bitb_49_33 word49_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_33 q_50_33 qb_50_33 bit_50_33 bitb_50_33 word50_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_33 q_51_33 qb_51_33 bit_51_33 bitb_51_33 word51_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_33 q_52_33 qb_52_33 bit_52_33 bitb_52_33 word52_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_33 q_53_33 qb_53_33 bit_53_33 bitb_53_33 word53_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_33 q_54_33 qb_54_33 bit_54_33 bitb_54_33 word54_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_33 q_55_33 qb_55_33 bit_55_33 bitb_55_33 word55_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_33 q_56_33 qb_56_33 bit_56_33 bitb_56_33 word56_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_33 q_57_33 qb_57_33 bit_57_33 bitb_57_33 word57_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_33 q_58_33 qb_58_33 bit_58_33 bitb_58_33 word58_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_33 q_59_33 qb_59_33 bit_59_33 bitb_59_33 word59_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_33 q_60_33 qb_60_33 bit_60_33 bitb_60_33 word60_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_33 q_61_33 qb_61_33 bit_61_33 bitb_61_33 word61_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_33 q_62_33 qb_62_33 bit_62_33 bitb_62_33 word62_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_33 q_63_33 qb_63_33 bit_63_33 bitb_63_33 word63_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_33 q_64_33 qb_64_33 bit_64_33 bitb_64_33 word64_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_33 q_65_33 qb_65_33 bit_65_33 bitb_65_33 word65_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_33 q_66_33 qb_66_33 bit_66_33 bitb_66_33 word66_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_33 q_67_33 qb_67_33 bit_67_33 bitb_67_33 word67_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_33 q_68_33 qb_68_33 bit_68_33 bitb_68_33 word68_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_33 q_69_33 qb_69_33 bit_69_33 bitb_69_33 word69_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_33 q_70_33 qb_70_33 bit_70_33 bitb_70_33 word70_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_33 q_71_33 qb_71_33 bit_71_33 bitb_71_33 word71_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_33 q_72_33 qb_72_33 bit_72_33 bitb_72_33 word72_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_33 q_73_33 qb_73_33 bit_73_33 bitb_73_33 word73_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_33 q_74_33 qb_74_33 bit_74_33 bitb_74_33 word74_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_33 q_75_33 qb_75_33 bit_75_33 bitb_75_33 word75_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_33 q_76_33 qb_76_33 bit_76_33 bitb_76_33 word76_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_33 q_77_33 qb_77_33 bit_77_33 bitb_77_33 word77_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_33 q_78_33 qb_78_33 bit_78_33 bitb_78_33 word78_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_33 q_79_33 qb_79_33 bit_79_33 bitb_79_33 word79_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_33 q_80_33 qb_80_33 bit_80_33 bitb_80_33 word80_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_33 q_81_33 qb_81_33 bit_81_33 bitb_81_33 word81_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_33 q_82_33 qb_82_33 bit_82_33 bitb_82_33 word82_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_33 q_83_33 qb_83_33 bit_83_33 bitb_83_33 word83_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_33 q_84_33 qb_84_33 bit_84_33 bitb_84_33 word84_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_33 q_85_33 qb_85_33 bit_85_33 bitb_85_33 word85_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_33 q_86_33 qb_86_33 bit_86_33 bitb_86_33 word86_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_33 q_87_33 qb_87_33 bit_87_33 bitb_87_33 word87_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_33 q_88_33 qb_88_33 bit_88_33 bitb_88_33 word88_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_33 q_89_33 qb_89_33 bit_89_33 bitb_89_33 word89_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_33 q_90_33 qb_90_33 bit_90_33 bitb_90_33 word90_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_33 q_91_33 qb_91_33 bit_91_33 bitb_91_33 word91_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_33 q_92_33 qb_92_33 bit_92_33 bitb_92_33 word92_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_33 q_93_33 qb_93_33 bit_93_33 bitb_93_33 word93_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_33 q_94_33 qb_94_33 bit_94_33 bitb_94_33 word94_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_33 q_95_33 qb_95_33 bit_95_33 bitb_95_33 word95_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_33 q_96_33 qb_96_33 bit_96_33 bitb_96_33 word96_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_33 q_97_33 qb_97_33 bit_97_33 bitb_97_33 word97_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_33 q_98_33 qb_98_33 bit_98_33 bitb_98_33 word98_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_33 q_99_33 qb_99_33 bit_99_33 bitb_99_33 word99_33 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_34 q_0_34 qb_0_34 bit_0_34 bitb_0_34 word0_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_34 q_1_34 qb_1_34 bit_1_34 bitb_1_34 word1_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_34 q_2_34 qb_2_34 bit_2_34 bitb_2_34 word2_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_34 q_3_34 qb_3_34 bit_3_34 bitb_3_34 word3_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_34 q_4_34 qb_4_34 bit_4_34 bitb_4_34 word4_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_34 q_5_34 qb_5_34 bit_5_34 bitb_5_34 word5_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_34 q_6_34 qb_6_34 bit_6_34 bitb_6_34 word6_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_34 q_7_34 qb_7_34 bit_7_34 bitb_7_34 word7_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_34 q_8_34 qb_8_34 bit_8_34 bitb_8_34 word8_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_34 q_9_34 qb_9_34 bit_9_34 bitb_9_34 word9_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_34 q_10_34 qb_10_34 bit_10_34 bitb_10_34 word10_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_34 q_11_34 qb_11_34 bit_11_34 bitb_11_34 word11_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_34 q_12_34 qb_12_34 bit_12_34 bitb_12_34 word12_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_34 q_13_34 qb_13_34 bit_13_34 bitb_13_34 word13_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_34 q_14_34 qb_14_34 bit_14_34 bitb_14_34 word14_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_34 q_15_34 qb_15_34 bit_15_34 bitb_15_34 word15_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_34 q_16_34 qb_16_34 bit_16_34 bitb_16_34 word16_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_34 q_17_34 qb_17_34 bit_17_34 bitb_17_34 word17_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_34 q_18_34 qb_18_34 bit_18_34 bitb_18_34 word18_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_34 q_19_34 qb_19_34 bit_19_34 bitb_19_34 word19_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_34 q_20_34 qb_20_34 bit_20_34 bitb_20_34 word20_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_34 q_21_34 qb_21_34 bit_21_34 bitb_21_34 word21_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_34 q_22_34 qb_22_34 bit_22_34 bitb_22_34 word22_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_34 q_23_34 qb_23_34 bit_23_34 bitb_23_34 word23_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_34 q_24_34 qb_24_34 bit_24_34 bitb_24_34 word24_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_34 q_25_34 qb_25_34 bit_25_34 bitb_25_34 word25_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_34 q_26_34 qb_26_34 bit_26_34 bitb_26_34 word26_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_34 q_27_34 qb_27_34 bit_27_34 bitb_27_34 word27_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_34 q_28_34 qb_28_34 bit_28_34 bitb_28_34 word28_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_34 q_29_34 qb_29_34 bit_29_34 bitb_29_34 word29_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_34 q_30_34 qb_30_34 bit_30_34 bitb_30_34 word30_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_34 q_31_34 qb_31_34 bit_31_34 bitb_31_34 word31_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_34 q_32_34 qb_32_34 bit_32_34 bitb_32_34 word32_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_34 q_33_34 qb_33_34 bit_33_34 bitb_33_34 word33_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_34 q_34_34 qb_34_34 bit_34_34 bitb_34_34 word34_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_34 q_35_34 qb_35_34 bit_35_34 bitb_35_34 word35_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_34 q_36_34 qb_36_34 bit_36_34 bitb_36_34 word36_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_34 q_37_34 qb_37_34 bit_37_34 bitb_37_34 word37_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_34 q_38_34 qb_38_34 bit_38_34 bitb_38_34 word38_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_34 q_39_34 qb_39_34 bit_39_34 bitb_39_34 word39_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_34 q_40_34 qb_40_34 bit_40_34 bitb_40_34 word40_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_34 q_41_34 qb_41_34 bit_41_34 bitb_41_34 word41_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_34 q_42_34 qb_42_34 bit_42_34 bitb_42_34 word42_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_34 q_43_34 qb_43_34 bit_43_34 bitb_43_34 word43_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_34 q_44_34 qb_44_34 bit_44_34 bitb_44_34 word44_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_34 q_45_34 qb_45_34 bit_45_34 bitb_45_34 word45_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_34 q_46_34 qb_46_34 bit_46_34 bitb_46_34 word46_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_34 q_47_34 qb_47_34 bit_47_34 bitb_47_34 word47_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_34 q_48_34 qb_48_34 bit_48_34 bitb_48_34 word48_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_34 q_49_34 qb_49_34 bit_49_34 bitb_49_34 word49_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_34 q_50_34 qb_50_34 bit_50_34 bitb_50_34 word50_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_34 q_51_34 qb_51_34 bit_51_34 bitb_51_34 word51_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_34 q_52_34 qb_52_34 bit_52_34 bitb_52_34 word52_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_34 q_53_34 qb_53_34 bit_53_34 bitb_53_34 word53_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_34 q_54_34 qb_54_34 bit_54_34 bitb_54_34 word54_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_34 q_55_34 qb_55_34 bit_55_34 bitb_55_34 word55_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_34 q_56_34 qb_56_34 bit_56_34 bitb_56_34 word56_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_34 q_57_34 qb_57_34 bit_57_34 bitb_57_34 word57_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_34 q_58_34 qb_58_34 bit_58_34 bitb_58_34 word58_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_34 q_59_34 qb_59_34 bit_59_34 bitb_59_34 word59_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_34 q_60_34 qb_60_34 bit_60_34 bitb_60_34 word60_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_34 q_61_34 qb_61_34 bit_61_34 bitb_61_34 word61_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_34 q_62_34 qb_62_34 bit_62_34 bitb_62_34 word62_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_34 q_63_34 qb_63_34 bit_63_34 bitb_63_34 word63_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_34 q_64_34 qb_64_34 bit_64_34 bitb_64_34 word64_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_34 q_65_34 qb_65_34 bit_65_34 bitb_65_34 word65_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_34 q_66_34 qb_66_34 bit_66_34 bitb_66_34 word66_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_34 q_67_34 qb_67_34 bit_67_34 bitb_67_34 word67_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_34 q_68_34 qb_68_34 bit_68_34 bitb_68_34 word68_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_34 q_69_34 qb_69_34 bit_69_34 bitb_69_34 word69_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_34 q_70_34 qb_70_34 bit_70_34 bitb_70_34 word70_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_34 q_71_34 qb_71_34 bit_71_34 bitb_71_34 word71_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_34 q_72_34 qb_72_34 bit_72_34 bitb_72_34 word72_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_34 q_73_34 qb_73_34 bit_73_34 bitb_73_34 word73_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_34 q_74_34 qb_74_34 bit_74_34 bitb_74_34 word74_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_34 q_75_34 qb_75_34 bit_75_34 bitb_75_34 word75_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_34 q_76_34 qb_76_34 bit_76_34 bitb_76_34 word76_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_34 q_77_34 qb_77_34 bit_77_34 bitb_77_34 word77_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_34 q_78_34 qb_78_34 bit_78_34 bitb_78_34 word78_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_34 q_79_34 qb_79_34 bit_79_34 bitb_79_34 word79_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_34 q_80_34 qb_80_34 bit_80_34 bitb_80_34 word80_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_34 q_81_34 qb_81_34 bit_81_34 bitb_81_34 word81_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_34 q_82_34 qb_82_34 bit_82_34 bitb_82_34 word82_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_34 q_83_34 qb_83_34 bit_83_34 bitb_83_34 word83_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_34 q_84_34 qb_84_34 bit_84_34 bitb_84_34 word84_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_34 q_85_34 qb_85_34 bit_85_34 bitb_85_34 word85_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_34 q_86_34 qb_86_34 bit_86_34 bitb_86_34 word86_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_34 q_87_34 qb_87_34 bit_87_34 bitb_87_34 word87_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_34 q_88_34 qb_88_34 bit_88_34 bitb_88_34 word88_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_34 q_89_34 qb_89_34 bit_89_34 bitb_89_34 word89_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_34 q_90_34 qb_90_34 bit_90_34 bitb_90_34 word90_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_34 q_91_34 qb_91_34 bit_91_34 bitb_91_34 word91_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_34 q_92_34 qb_92_34 bit_92_34 bitb_92_34 word92_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_34 q_93_34 qb_93_34 bit_93_34 bitb_93_34 word93_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_34 q_94_34 qb_94_34 bit_94_34 bitb_94_34 word94_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_34 q_95_34 qb_95_34 bit_95_34 bitb_95_34 word95_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_34 q_96_34 qb_96_34 bit_96_34 bitb_96_34 word96_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_34 q_97_34 qb_97_34 bit_97_34 bitb_97_34 word97_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_34 q_98_34 qb_98_34 bit_98_34 bitb_98_34 word98_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_34 q_99_34 qb_99_34 bit_99_34 bitb_99_34 word99_34 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_35 q_0_35 qb_0_35 bit_0_35 bitb_0_35 word0_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_35 q_1_35 qb_1_35 bit_1_35 bitb_1_35 word1_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_35 q_2_35 qb_2_35 bit_2_35 bitb_2_35 word2_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_35 q_3_35 qb_3_35 bit_3_35 bitb_3_35 word3_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_35 q_4_35 qb_4_35 bit_4_35 bitb_4_35 word4_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_35 q_5_35 qb_5_35 bit_5_35 bitb_5_35 word5_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_35 q_6_35 qb_6_35 bit_6_35 bitb_6_35 word6_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_35 q_7_35 qb_7_35 bit_7_35 bitb_7_35 word7_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_35 q_8_35 qb_8_35 bit_8_35 bitb_8_35 word8_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_35 q_9_35 qb_9_35 bit_9_35 bitb_9_35 word9_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_35 q_10_35 qb_10_35 bit_10_35 bitb_10_35 word10_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_35 q_11_35 qb_11_35 bit_11_35 bitb_11_35 word11_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_35 q_12_35 qb_12_35 bit_12_35 bitb_12_35 word12_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_35 q_13_35 qb_13_35 bit_13_35 bitb_13_35 word13_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_35 q_14_35 qb_14_35 bit_14_35 bitb_14_35 word14_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_35 q_15_35 qb_15_35 bit_15_35 bitb_15_35 word15_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_35 q_16_35 qb_16_35 bit_16_35 bitb_16_35 word16_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_35 q_17_35 qb_17_35 bit_17_35 bitb_17_35 word17_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_35 q_18_35 qb_18_35 bit_18_35 bitb_18_35 word18_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_35 q_19_35 qb_19_35 bit_19_35 bitb_19_35 word19_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_35 q_20_35 qb_20_35 bit_20_35 bitb_20_35 word20_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_35 q_21_35 qb_21_35 bit_21_35 bitb_21_35 word21_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_35 q_22_35 qb_22_35 bit_22_35 bitb_22_35 word22_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_35 q_23_35 qb_23_35 bit_23_35 bitb_23_35 word23_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_35 q_24_35 qb_24_35 bit_24_35 bitb_24_35 word24_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_35 q_25_35 qb_25_35 bit_25_35 bitb_25_35 word25_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_35 q_26_35 qb_26_35 bit_26_35 bitb_26_35 word26_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_35 q_27_35 qb_27_35 bit_27_35 bitb_27_35 word27_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_35 q_28_35 qb_28_35 bit_28_35 bitb_28_35 word28_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_35 q_29_35 qb_29_35 bit_29_35 bitb_29_35 word29_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_35 q_30_35 qb_30_35 bit_30_35 bitb_30_35 word30_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_35 q_31_35 qb_31_35 bit_31_35 bitb_31_35 word31_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_35 q_32_35 qb_32_35 bit_32_35 bitb_32_35 word32_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_35 q_33_35 qb_33_35 bit_33_35 bitb_33_35 word33_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_35 q_34_35 qb_34_35 bit_34_35 bitb_34_35 word34_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_35 q_35_35 qb_35_35 bit_35_35 bitb_35_35 word35_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_35 q_36_35 qb_36_35 bit_36_35 bitb_36_35 word36_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_35 q_37_35 qb_37_35 bit_37_35 bitb_37_35 word37_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_35 q_38_35 qb_38_35 bit_38_35 bitb_38_35 word38_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_35 q_39_35 qb_39_35 bit_39_35 bitb_39_35 word39_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_35 q_40_35 qb_40_35 bit_40_35 bitb_40_35 word40_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_35 q_41_35 qb_41_35 bit_41_35 bitb_41_35 word41_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_35 q_42_35 qb_42_35 bit_42_35 bitb_42_35 word42_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_35 q_43_35 qb_43_35 bit_43_35 bitb_43_35 word43_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_35 q_44_35 qb_44_35 bit_44_35 bitb_44_35 word44_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_35 q_45_35 qb_45_35 bit_45_35 bitb_45_35 word45_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_35 q_46_35 qb_46_35 bit_46_35 bitb_46_35 word46_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_35 q_47_35 qb_47_35 bit_47_35 bitb_47_35 word47_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_35 q_48_35 qb_48_35 bit_48_35 bitb_48_35 word48_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_35 q_49_35 qb_49_35 bit_49_35 bitb_49_35 word49_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_35 q_50_35 qb_50_35 bit_50_35 bitb_50_35 word50_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_35 q_51_35 qb_51_35 bit_51_35 bitb_51_35 word51_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_35 q_52_35 qb_52_35 bit_52_35 bitb_52_35 word52_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_35 q_53_35 qb_53_35 bit_53_35 bitb_53_35 word53_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_35 q_54_35 qb_54_35 bit_54_35 bitb_54_35 word54_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_35 q_55_35 qb_55_35 bit_55_35 bitb_55_35 word55_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_35 q_56_35 qb_56_35 bit_56_35 bitb_56_35 word56_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_35 q_57_35 qb_57_35 bit_57_35 bitb_57_35 word57_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_35 q_58_35 qb_58_35 bit_58_35 bitb_58_35 word58_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_35 q_59_35 qb_59_35 bit_59_35 bitb_59_35 word59_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_35 q_60_35 qb_60_35 bit_60_35 bitb_60_35 word60_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_35 q_61_35 qb_61_35 bit_61_35 bitb_61_35 word61_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_35 q_62_35 qb_62_35 bit_62_35 bitb_62_35 word62_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_35 q_63_35 qb_63_35 bit_63_35 bitb_63_35 word63_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_35 q_64_35 qb_64_35 bit_64_35 bitb_64_35 word64_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_35 q_65_35 qb_65_35 bit_65_35 bitb_65_35 word65_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_35 q_66_35 qb_66_35 bit_66_35 bitb_66_35 word66_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_35 q_67_35 qb_67_35 bit_67_35 bitb_67_35 word67_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_35 q_68_35 qb_68_35 bit_68_35 bitb_68_35 word68_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_35 q_69_35 qb_69_35 bit_69_35 bitb_69_35 word69_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_35 q_70_35 qb_70_35 bit_70_35 bitb_70_35 word70_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_35 q_71_35 qb_71_35 bit_71_35 bitb_71_35 word71_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_35 q_72_35 qb_72_35 bit_72_35 bitb_72_35 word72_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_35 q_73_35 qb_73_35 bit_73_35 bitb_73_35 word73_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_35 q_74_35 qb_74_35 bit_74_35 bitb_74_35 word74_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_35 q_75_35 qb_75_35 bit_75_35 bitb_75_35 word75_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_35 q_76_35 qb_76_35 bit_76_35 bitb_76_35 word76_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_35 q_77_35 qb_77_35 bit_77_35 bitb_77_35 word77_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_35 q_78_35 qb_78_35 bit_78_35 bitb_78_35 word78_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_35 q_79_35 qb_79_35 bit_79_35 bitb_79_35 word79_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_35 q_80_35 qb_80_35 bit_80_35 bitb_80_35 word80_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_35 q_81_35 qb_81_35 bit_81_35 bitb_81_35 word81_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_35 q_82_35 qb_82_35 bit_82_35 bitb_82_35 word82_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_35 q_83_35 qb_83_35 bit_83_35 bitb_83_35 word83_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_35 q_84_35 qb_84_35 bit_84_35 bitb_84_35 word84_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_35 q_85_35 qb_85_35 bit_85_35 bitb_85_35 word85_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_35 q_86_35 qb_86_35 bit_86_35 bitb_86_35 word86_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_35 q_87_35 qb_87_35 bit_87_35 bitb_87_35 word87_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_35 q_88_35 qb_88_35 bit_88_35 bitb_88_35 word88_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_35 q_89_35 qb_89_35 bit_89_35 bitb_89_35 word89_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_35 q_90_35 qb_90_35 bit_90_35 bitb_90_35 word90_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_35 q_91_35 qb_91_35 bit_91_35 bitb_91_35 word91_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_35 q_92_35 qb_92_35 bit_92_35 bitb_92_35 word92_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_35 q_93_35 qb_93_35 bit_93_35 bitb_93_35 word93_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_35 q_94_35 qb_94_35 bit_94_35 bitb_94_35 word94_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_35 q_95_35 qb_95_35 bit_95_35 bitb_95_35 word95_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_35 q_96_35 qb_96_35 bit_96_35 bitb_96_35 word96_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_35 q_97_35 qb_97_35 bit_97_35 bitb_97_35 word97_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_35 q_98_35 qb_98_35 bit_98_35 bitb_98_35 word98_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_35 q_99_35 qb_99_35 bit_99_35 bitb_99_35 word99_35 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_36 q_0_36 qb_0_36 bit_0_36 bitb_0_36 word0_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_36 q_1_36 qb_1_36 bit_1_36 bitb_1_36 word1_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_36 q_2_36 qb_2_36 bit_2_36 bitb_2_36 word2_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_36 q_3_36 qb_3_36 bit_3_36 bitb_3_36 word3_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_36 q_4_36 qb_4_36 bit_4_36 bitb_4_36 word4_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_36 q_5_36 qb_5_36 bit_5_36 bitb_5_36 word5_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_36 q_6_36 qb_6_36 bit_6_36 bitb_6_36 word6_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_36 q_7_36 qb_7_36 bit_7_36 bitb_7_36 word7_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_36 q_8_36 qb_8_36 bit_8_36 bitb_8_36 word8_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_36 q_9_36 qb_9_36 bit_9_36 bitb_9_36 word9_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_36 q_10_36 qb_10_36 bit_10_36 bitb_10_36 word10_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_36 q_11_36 qb_11_36 bit_11_36 bitb_11_36 word11_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_36 q_12_36 qb_12_36 bit_12_36 bitb_12_36 word12_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_36 q_13_36 qb_13_36 bit_13_36 bitb_13_36 word13_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_36 q_14_36 qb_14_36 bit_14_36 bitb_14_36 word14_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_36 q_15_36 qb_15_36 bit_15_36 bitb_15_36 word15_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_36 q_16_36 qb_16_36 bit_16_36 bitb_16_36 word16_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_36 q_17_36 qb_17_36 bit_17_36 bitb_17_36 word17_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_36 q_18_36 qb_18_36 bit_18_36 bitb_18_36 word18_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_36 q_19_36 qb_19_36 bit_19_36 bitb_19_36 word19_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_36 q_20_36 qb_20_36 bit_20_36 bitb_20_36 word20_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_36 q_21_36 qb_21_36 bit_21_36 bitb_21_36 word21_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_36 q_22_36 qb_22_36 bit_22_36 bitb_22_36 word22_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_36 q_23_36 qb_23_36 bit_23_36 bitb_23_36 word23_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_36 q_24_36 qb_24_36 bit_24_36 bitb_24_36 word24_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_36 q_25_36 qb_25_36 bit_25_36 bitb_25_36 word25_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_36 q_26_36 qb_26_36 bit_26_36 bitb_26_36 word26_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_36 q_27_36 qb_27_36 bit_27_36 bitb_27_36 word27_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_36 q_28_36 qb_28_36 bit_28_36 bitb_28_36 word28_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_36 q_29_36 qb_29_36 bit_29_36 bitb_29_36 word29_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_36 q_30_36 qb_30_36 bit_30_36 bitb_30_36 word30_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_36 q_31_36 qb_31_36 bit_31_36 bitb_31_36 word31_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_36 q_32_36 qb_32_36 bit_32_36 bitb_32_36 word32_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_36 q_33_36 qb_33_36 bit_33_36 bitb_33_36 word33_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_36 q_34_36 qb_34_36 bit_34_36 bitb_34_36 word34_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_36 q_35_36 qb_35_36 bit_35_36 bitb_35_36 word35_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_36 q_36_36 qb_36_36 bit_36_36 bitb_36_36 word36_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_36 q_37_36 qb_37_36 bit_37_36 bitb_37_36 word37_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_36 q_38_36 qb_38_36 bit_38_36 bitb_38_36 word38_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_36 q_39_36 qb_39_36 bit_39_36 bitb_39_36 word39_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_36 q_40_36 qb_40_36 bit_40_36 bitb_40_36 word40_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_36 q_41_36 qb_41_36 bit_41_36 bitb_41_36 word41_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_36 q_42_36 qb_42_36 bit_42_36 bitb_42_36 word42_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_36 q_43_36 qb_43_36 bit_43_36 bitb_43_36 word43_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_36 q_44_36 qb_44_36 bit_44_36 bitb_44_36 word44_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_36 q_45_36 qb_45_36 bit_45_36 bitb_45_36 word45_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_36 q_46_36 qb_46_36 bit_46_36 bitb_46_36 word46_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_36 q_47_36 qb_47_36 bit_47_36 bitb_47_36 word47_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_36 q_48_36 qb_48_36 bit_48_36 bitb_48_36 word48_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_36 q_49_36 qb_49_36 bit_49_36 bitb_49_36 word49_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_36 q_50_36 qb_50_36 bit_50_36 bitb_50_36 word50_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_36 q_51_36 qb_51_36 bit_51_36 bitb_51_36 word51_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_36 q_52_36 qb_52_36 bit_52_36 bitb_52_36 word52_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_36 q_53_36 qb_53_36 bit_53_36 bitb_53_36 word53_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_36 q_54_36 qb_54_36 bit_54_36 bitb_54_36 word54_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_36 q_55_36 qb_55_36 bit_55_36 bitb_55_36 word55_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_36 q_56_36 qb_56_36 bit_56_36 bitb_56_36 word56_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_36 q_57_36 qb_57_36 bit_57_36 bitb_57_36 word57_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_36 q_58_36 qb_58_36 bit_58_36 bitb_58_36 word58_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_36 q_59_36 qb_59_36 bit_59_36 bitb_59_36 word59_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_36 q_60_36 qb_60_36 bit_60_36 bitb_60_36 word60_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_36 q_61_36 qb_61_36 bit_61_36 bitb_61_36 word61_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_36 q_62_36 qb_62_36 bit_62_36 bitb_62_36 word62_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_36 q_63_36 qb_63_36 bit_63_36 bitb_63_36 word63_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_36 q_64_36 qb_64_36 bit_64_36 bitb_64_36 word64_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_36 q_65_36 qb_65_36 bit_65_36 bitb_65_36 word65_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_36 q_66_36 qb_66_36 bit_66_36 bitb_66_36 word66_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_36 q_67_36 qb_67_36 bit_67_36 bitb_67_36 word67_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_36 q_68_36 qb_68_36 bit_68_36 bitb_68_36 word68_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_36 q_69_36 qb_69_36 bit_69_36 bitb_69_36 word69_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_36 q_70_36 qb_70_36 bit_70_36 bitb_70_36 word70_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_36 q_71_36 qb_71_36 bit_71_36 bitb_71_36 word71_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_36 q_72_36 qb_72_36 bit_72_36 bitb_72_36 word72_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_36 q_73_36 qb_73_36 bit_73_36 bitb_73_36 word73_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_36 q_74_36 qb_74_36 bit_74_36 bitb_74_36 word74_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_36 q_75_36 qb_75_36 bit_75_36 bitb_75_36 word75_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_36 q_76_36 qb_76_36 bit_76_36 bitb_76_36 word76_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_36 q_77_36 qb_77_36 bit_77_36 bitb_77_36 word77_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_36 q_78_36 qb_78_36 bit_78_36 bitb_78_36 word78_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_36 q_79_36 qb_79_36 bit_79_36 bitb_79_36 word79_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_36 q_80_36 qb_80_36 bit_80_36 bitb_80_36 word80_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_36 q_81_36 qb_81_36 bit_81_36 bitb_81_36 word81_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_36 q_82_36 qb_82_36 bit_82_36 bitb_82_36 word82_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_36 q_83_36 qb_83_36 bit_83_36 bitb_83_36 word83_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_36 q_84_36 qb_84_36 bit_84_36 bitb_84_36 word84_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_36 q_85_36 qb_85_36 bit_85_36 bitb_85_36 word85_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_36 q_86_36 qb_86_36 bit_86_36 bitb_86_36 word86_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_36 q_87_36 qb_87_36 bit_87_36 bitb_87_36 word87_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_36 q_88_36 qb_88_36 bit_88_36 bitb_88_36 word88_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_36 q_89_36 qb_89_36 bit_89_36 bitb_89_36 word89_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_36 q_90_36 qb_90_36 bit_90_36 bitb_90_36 word90_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_36 q_91_36 qb_91_36 bit_91_36 bitb_91_36 word91_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_36 q_92_36 qb_92_36 bit_92_36 bitb_92_36 word92_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_36 q_93_36 qb_93_36 bit_93_36 bitb_93_36 word93_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_36 q_94_36 qb_94_36 bit_94_36 bitb_94_36 word94_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_36 q_95_36 qb_95_36 bit_95_36 bitb_95_36 word95_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_36 q_96_36 qb_96_36 bit_96_36 bitb_96_36 word96_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_36 q_97_36 qb_97_36 bit_97_36 bitb_97_36 word97_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_36 q_98_36 qb_98_36 bit_98_36 bitb_98_36 word98_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_36 q_99_36 qb_99_36 bit_99_36 bitb_99_36 word99_36 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_37 q_0_37 qb_0_37 bit_0_37 bitb_0_37 word0_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_37 q_1_37 qb_1_37 bit_1_37 bitb_1_37 word1_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_37 q_2_37 qb_2_37 bit_2_37 bitb_2_37 word2_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_37 q_3_37 qb_3_37 bit_3_37 bitb_3_37 word3_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_37 q_4_37 qb_4_37 bit_4_37 bitb_4_37 word4_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_37 q_5_37 qb_5_37 bit_5_37 bitb_5_37 word5_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_37 q_6_37 qb_6_37 bit_6_37 bitb_6_37 word6_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_37 q_7_37 qb_7_37 bit_7_37 bitb_7_37 word7_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_37 q_8_37 qb_8_37 bit_8_37 bitb_8_37 word8_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_37 q_9_37 qb_9_37 bit_9_37 bitb_9_37 word9_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_37 q_10_37 qb_10_37 bit_10_37 bitb_10_37 word10_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_37 q_11_37 qb_11_37 bit_11_37 bitb_11_37 word11_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_37 q_12_37 qb_12_37 bit_12_37 bitb_12_37 word12_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_37 q_13_37 qb_13_37 bit_13_37 bitb_13_37 word13_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_37 q_14_37 qb_14_37 bit_14_37 bitb_14_37 word14_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_37 q_15_37 qb_15_37 bit_15_37 bitb_15_37 word15_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_37 q_16_37 qb_16_37 bit_16_37 bitb_16_37 word16_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_37 q_17_37 qb_17_37 bit_17_37 bitb_17_37 word17_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_37 q_18_37 qb_18_37 bit_18_37 bitb_18_37 word18_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_37 q_19_37 qb_19_37 bit_19_37 bitb_19_37 word19_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_37 q_20_37 qb_20_37 bit_20_37 bitb_20_37 word20_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_37 q_21_37 qb_21_37 bit_21_37 bitb_21_37 word21_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_37 q_22_37 qb_22_37 bit_22_37 bitb_22_37 word22_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_37 q_23_37 qb_23_37 bit_23_37 bitb_23_37 word23_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_37 q_24_37 qb_24_37 bit_24_37 bitb_24_37 word24_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_37 q_25_37 qb_25_37 bit_25_37 bitb_25_37 word25_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_37 q_26_37 qb_26_37 bit_26_37 bitb_26_37 word26_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_37 q_27_37 qb_27_37 bit_27_37 bitb_27_37 word27_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_37 q_28_37 qb_28_37 bit_28_37 bitb_28_37 word28_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_37 q_29_37 qb_29_37 bit_29_37 bitb_29_37 word29_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_37 q_30_37 qb_30_37 bit_30_37 bitb_30_37 word30_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_37 q_31_37 qb_31_37 bit_31_37 bitb_31_37 word31_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_37 q_32_37 qb_32_37 bit_32_37 bitb_32_37 word32_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_37 q_33_37 qb_33_37 bit_33_37 bitb_33_37 word33_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_37 q_34_37 qb_34_37 bit_34_37 bitb_34_37 word34_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_37 q_35_37 qb_35_37 bit_35_37 bitb_35_37 word35_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_37 q_36_37 qb_36_37 bit_36_37 bitb_36_37 word36_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_37 q_37_37 qb_37_37 bit_37_37 bitb_37_37 word37_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_37 q_38_37 qb_38_37 bit_38_37 bitb_38_37 word38_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_37 q_39_37 qb_39_37 bit_39_37 bitb_39_37 word39_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_37 q_40_37 qb_40_37 bit_40_37 bitb_40_37 word40_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_37 q_41_37 qb_41_37 bit_41_37 bitb_41_37 word41_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_37 q_42_37 qb_42_37 bit_42_37 bitb_42_37 word42_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_37 q_43_37 qb_43_37 bit_43_37 bitb_43_37 word43_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_37 q_44_37 qb_44_37 bit_44_37 bitb_44_37 word44_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_37 q_45_37 qb_45_37 bit_45_37 bitb_45_37 word45_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_37 q_46_37 qb_46_37 bit_46_37 bitb_46_37 word46_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_37 q_47_37 qb_47_37 bit_47_37 bitb_47_37 word47_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_37 q_48_37 qb_48_37 bit_48_37 bitb_48_37 word48_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_37 q_49_37 qb_49_37 bit_49_37 bitb_49_37 word49_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_37 q_50_37 qb_50_37 bit_50_37 bitb_50_37 word50_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_37 q_51_37 qb_51_37 bit_51_37 bitb_51_37 word51_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_37 q_52_37 qb_52_37 bit_52_37 bitb_52_37 word52_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_37 q_53_37 qb_53_37 bit_53_37 bitb_53_37 word53_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_37 q_54_37 qb_54_37 bit_54_37 bitb_54_37 word54_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_37 q_55_37 qb_55_37 bit_55_37 bitb_55_37 word55_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_37 q_56_37 qb_56_37 bit_56_37 bitb_56_37 word56_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_37 q_57_37 qb_57_37 bit_57_37 bitb_57_37 word57_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_37 q_58_37 qb_58_37 bit_58_37 bitb_58_37 word58_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_37 q_59_37 qb_59_37 bit_59_37 bitb_59_37 word59_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_37 q_60_37 qb_60_37 bit_60_37 bitb_60_37 word60_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_37 q_61_37 qb_61_37 bit_61_37 bitb_61_37 word61_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_37 q_62_37 qb_62_37 bit_62_37 bitb_62_37 word62_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_37 q_63_37 qb_63_37 bit_63_37 bitb_63_37 word63_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_37 q_64_37 qb_64_37 bit_64_37 bitb_64_37 word64_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_37 q_65_37 qb_65_37 bit_65_37 bitb_65_37 word65_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_37 q_66_37 qb_66_37 bit_66_37 bitb_66_37 word66_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_37 q_67_37 qb_67_37 bit_67_37 bitb_67_37 word67_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_37 q_68_37 qb_68_37 bit_68_37 bitb_68_37 word68_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_37 q_69_37 qb_69_37 bit_69_37 bitb_69_37 word69_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_37 q_70_37 qb_70_37 bit_70_37 bitb_70_37 word70_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_37 q_71_37 qb_71_37 bit_71_37 bitb_71_37 word71_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_37 q_72_37 qb_72_37 bit_72_37 bitb_72_37 word72_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_37 q_73_37 qb_73_37 bit_73_37 bitb_73_37 word73_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_37 q_74_37 qb_74_37 bit_74_37 bitb_74_37 word74_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_37 q_75_37 qb_75_37 bit_75_37 bitb_75_37 word75_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_37 q_76_37 qb_76_37 bit_76_37 bitb_76_37 word76_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_37 q_77_37 qb_77_37 bit_77_37 bitb_77_37 word77_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_37 q_78_37 qb_78_37 bit_78_37 bitb_78_37 word78_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_37 q_79_37 qb_79_37 bit_79_37 bitb_79_37 word79_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_37 q_80_37 qb_80_37 bit_80_37 bitb_80_37 word80_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_37 q_81_37 qb_81_37 bit_81_37 bitb_81_37 word81_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_37 q_82_37 qb_82_37 bit_82_37 bitb_82_37 word82_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_37 q_83_37 qb_83_37 bit_83_37 bitb_83_37 word83_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_37 q_84_37 qb_84_37 bit_84_37 bitb_84_37 word84_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_37 q_85_37 qb_85_37 bit_85_37 bitb_85_37 word85_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_37 q_86_37 qb_86_37 bit_86_37 bitb_86_37 word86_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_37 q_87_37 qb_87_37 bit_87_37 bitb_87_37 word87_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_37 q_88_37 qb_88_37 bit_88_37 bitb_88_37 word88_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_37 q_89_37 qb_89_37 bit_89_37 bitb_89_37 word89_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_37 q_90_37 qb_90_37 bit_90_37 bitb_90_37 word90_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_37 q_91_37 qb_91_37 bit_91_37 bitb_91_37 word91_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_37 q_92_37 qb_92_37 bit_92_37 bitb_92_37 word92_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_37 q_93_37 qb_93_37 bit_93_37 bitb_93_37 word93_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_37 q_94_37 qb_94_37 bit_94_37 bitb_94_37 word94_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_37 q_95_37 qb_95_37 bit_95_37 bitb_95_37 word95_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_37 q_96_37 qb_96_37 bit_96_37 bitb_96_37 word96_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_37 q_97_37 qb_97_37 bit_97_37 bitb_97_37 word97_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_37 q_98_37 qb_98_37 bit_98_37 bitb_98_37 word98_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_37 q_99_37 qb_99_37 bit_99_37 bitb_99_37 word99_37 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_38 q_0_38 qb_0_38 bit_0_38 bitb_0_38 word0_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_38 q_1_38 qb_1_38 bit_1_38 bitb_1_38 word1_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_38 q_2_38 qb_2_38 bit_2_38 bitb_2_38 word2_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_38 q_3_38 qb_3_38 bit_3_38 bitb_3_38 word3_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_38 q_4_38 qb_4_38 bit_4_38 bitb_4_38 word4_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_38 q_5_38 qb_5_38 bit_5_38 bitb_5_38 word5_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_38 q_6_38 qb_6_38 bit_6_38 bitb_6_38 word6_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_38 q_7_38 qb_7_38 bit_7_38 bitb_7_38 word7_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_38 q_8_38 qb_8_38 bit_8_38 bitb_8_38 word8_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_38 q_9_38 qb_9_38 bit_9_38 bitb_9_38 word9_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_38 q_10_38 qb_10_38 bit_10_38 bitb_10_38 word10_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_38 q_11_38 qb_11_38 bit_11_38 bitb_11_38 word11_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_38 q_12_38 qb_12_38 bit_12_38 bitb_12_38 word12_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_38 q_13_38 qb_13_38 bit_13_38 bitb_13_38 word13_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_38 q_14_38 qb_14_38 bit_14_38 bitb_14_38 word14_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_38 q_15_38 qb_15_38 bit_15_38 bitb_15_38 word15_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_38 q_16_38 qb_16_38 bit_16_38 bitb_16_38 word16_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_38 q_17_38 qb_17_38 bit_17_38 bitb_17_38 word17_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_38 q_18_38 qb_18_38 bit_18_38 bitb_18_38 word18_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_38 q_19_38 qb_19_38 bit_19_38 bitb_19_38 word19_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_38 q_20_38 qb_20_38 bit_20_38 bitb_20_38 word20_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_38 q_21_38 qb_21_38 bit_21_38 bitb_21_38 word21_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_38 q_22_38 qb_22_38 bit_22_38 bitb_22_38 word22_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_38 q_23_38 qb_23_38 bit_23_38 bitb_23_38 word23_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_38 q_24_38 qb_24_38 bit_24_38 bitb_24_38 word24_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_38 q_25_38 qb_25_38 bit_25_38 bitb_25_38 word25_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_38 q_26_38 qb_26_38 bit_26_38 bitb_26_38 word26_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_38 q_27_38 qb_27_38 bit_27_38 bitb_27_38 word27_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_38 q_28_38 qb_28_38 bit_28_38 bitb_28_38 word28_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_38 q_29_38 qb_29_38 bit_29_38 bitb_29_38 word29_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_38 q_30_38 qb_30_38 bit_30_38 bitb_30_38 word30_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_38 q_31_38 qb_31_38 bit_31_38 bitb_31_38 word31_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_38 q_32_38 qb_32_38 bit_32_38 bitb_32_38 word32_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_38 q_33_38 qb_33_38 bit_33_38 bitb_33_38 word33_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_38 q_34_38 qb_34_38 bit_34_38 bitb_34_38 word34_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_38 q_35_38 qb_35_38 bit_35_38 bitb_35_38 word35_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_38 q_36_38 qb_36_38 bit_36_38 bitb_36_38 word36_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_38 q_37_38 qb_37_38 bit_37_38 bitb_37_38 word37_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_38 q_38_38 qb_38_38 bit_38_38 bitb_38_38 word38_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_38 q_39_38 qb_39_38 bit_39_38 bitb_39_38 word39_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_38 q_40_38 qb_40_38 bit_40_38 bitb_40_38 word40_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_38 q_41_38 qb_41_38 bit_41_38 bitb_41_38 word41_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_38 q_42_38 qb_42_38 bit_42_38 bitb_42_38 word42_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_38 q_43_38 qb_43_38 bit_43_38 bitb_43_38 word43_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_38 q_44_38 qb_44_38 bit_44_38 bitb_44_38 word44_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_38 q_45_38 qb_45_38 bit_45_38 bitb_45_38 word45_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_38 q_46_38 qb_46_38 bit_46_38 bitb_46_38 word46_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_38 q_47_38 qb_47_38 bit_47_38 bitb_47_38 word47_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_38 q_48_38 qb_48_38 bit_48_38 bitb_48_38 word48_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_38 q_49_38 qb_49_38 bit_49_38 bitb_49_38 word49_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_38 q_50_38 qb_50_38 bit_50_38 bitb_50_38 word50_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_38 q_51_38 qb_51_38 bit_51_38 bitb_51_38 word51_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_38 q_52_38 qb_52_38 bit_52_38 bitb_52_38 word52_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_38 q_53_38 qb_53_38 bit_53_38 bitb_53_38 word53_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_38 q_54_38 qb_54_38 bit_54_38 bitb_54_38 word54_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_38 q_55_38 qb_55_38 bit_55_38 bitb_55_38 word55_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_38 q_56_38 qb_56_38 bit_56_38 bitb_56_38 word56_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_38 q_57_38 qb_57_38 bit_57_38 bitb_57_38 word57_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_38 q_58_38 qb_58_38 bit_58_38 bitb_58_38 word58_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_38 q_59_38 qb_59_38 bit_59_38 bitb_59_38 word59_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_38 q_60_38 qb_60_38 bit_60_38 bitb_60_38 word60_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_38 q_61_38 qb_61_38 bit_61_38 bitb_61_38 word61_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_38 q_62_38 qb_62_38 bit_62_38 bitb_62_38 word62_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_38 q_63_38 qb_63_38 bit_63_38 bitb_63_38 word63_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_38 q_64_38 qb_64_38 bit_64_38 bitb_64_38 word64_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_38 q_65_38 qb_65_38 bit_65_38 bitb_65_38 word65_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_38 q_66_38 qb_66_38 bit_66_38 bitb_66_38 word66_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_38 q_67_38 qb_67_38 bit_67_38 bitb_67_38 word67_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_38 q_68_38 qb_68_38 bit_68_38 bitb_68_38 word68_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_38 q_69_38 qb_69_38 bit_69_38 bitb_69_38 word69_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_38 q_70_38 qb_70_38 bit_70_38 bitb_70_38 word70_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_38 q_71_38 qb_71_38 bit_71_38 bitb_71_38 word71_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_38 q_72_38 qb_72_38 bit_72_38 bitb_72_38 word72_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_38 q_73_38 qb_73_38 bit_73_38 bitb_73_38 word73_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_38 q_74_38 qb_74_38 bit_74_38 bitb_74_38 word74_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_38 q_75_38 qb_75_38 bit_75_38 bitb_75_38 word75_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_38 q_76_38 qb_76_38 bit_76_38 bitb_76_38 word76_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_38 q_77_38 qb_77_38 bit_77_38 bitb_77_38 word77_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_38 q_78_38 qb_78_38 bit_78_38 bitb_78_38 word78_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_38 q_79_38 qb_79_38 bit_79_38 bitb_79_38 word79_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_38 q_80_38 qb_80_38 bit_80_38 bitb_80_38 word80_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_38 q_81_38 qb_81_38 bit_81_38 bitb_81_38 word81_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_38 q_82_38 qb_82_38 bit_82_38 bitb_82_38 word82_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_38 q_83_38 qb_83_38 bit_83_38 bitb_83_38 word83_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_38 q_84_38 qb_84_38 bit_84_38 bitb_84_38 word84_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_38 q_85_38 qb_85_38 bit_85_38 bitb_85_38 word85_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_38 q_86_38 qb_86_38 bit_86_38 bitb_86_38 word86_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_38 q_87_38 qb_87_38 bit_87_38 bitb_87_38 word87_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_38 q_88_38 qb_88_38 bit_88_38 bitb_88_38 word88_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_38 q_89_38 qb_89_38 bit_89_38 bitb_89_38 word89_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_38 q_90_38 qb_90_38 bit_90_38 bitb_90_38 word90_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_38 q_91_38 qb_91_38 bit_91_38 bitb_91_38 word91_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_38 q_92_38 qb_92_38 bit_92_38 bitb_92_38 word92_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_38 q_93_38 qb_93_38 bit_93_38 bitb_93_38 word93_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_38 q_94_38 qb_94_38 bit_94_38 bitb_94_38 word94_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_38 q_95_38 qb_95_38 bit_95_38 bitb_95_38 word95_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_38 q_96_38 qb_96_38 bit_96_38 bitb_96_38 word96_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_38 q_97_38 qb_97_38 bit_97_38 bitb_97_38 word97_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_38 q_98_38 qb_98_38 bit_98_38 bitb_98_38 word98_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_38 q_99_38 qb_99_38 bit_99_38 bitb_99_38 word99_38 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_39 q_0_39 qb_0_39 bit_0_39 bitb_0_39 word0_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_39 q_1_39 qb_1_39 bit_1_39 bitb_1_39 word1_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_39 q_2_39 qb_2_39 bit_2_39 bitb_2_39 word2_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_39 q_3_39 qb_3_39 bit_3_39 bitb_3_39 word3_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_39 q_4_39 qb_4_39 bit_4_39 bitb_4_39 word4_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_39 q_5_39 qb_5_39 bit_5_39 bitb_5_39 word5_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_39 q_6_39 qb_6_39 bit_6_39 bitb_6_39 word6_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_39 q_7_39 qb_7_39 bit_7_39 bitb_7_39 word7_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_39 q_8_39 qb_8_39 bit_8_39 bitb_8_39 word8_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_39 q_9_39 qb_9_39 bit_9_39 bitb_9_39 word9_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_39 q_10_39 qb_10_39 bit_10_39 bitb_10_39 word10_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_39 q_11_39 qb_11_39 bit_11_39 bitb_11_39 word11_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_39 q_12_39 qb_12_39 bit_12_39 bitb_12_39 word12_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_39 q_13_39 qb_13_39 bit_13_39 bitb_13_39 word13_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_39 q_14_39 qb_14_39 bit_14_39 bitb_14_39 word14_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_39 q_15_39 qb_15_39 bit_15_39 bitb_15_39 word15_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_39 q_16_39 qb_16_39 bit_16_39 bitb_16_39 word16_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_39 q_17_39 qb_17_39 bit_17_39 bitb_17_39 word17_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_39 q_18_39 qb_18_39 bit_18_39 bitb_18_39 word18_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_39 q_19_39 qb_19_39 bit_19_39 bitb_19_39 word19_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_39 q_20_39 qb_20_39 bit_20_39 bitb_20_39 word20_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_39 q_21_39 qb_21_39 bit_21_39 bitb_21_39 word21_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_39 q_22_39 qb_22_39 bit_22_39 bitb_22_39 word22_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_39 q_23_39 qb_23_39 bit_23_39 bitb_23_39 word23_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_39 q_24_39 qb_24_39 bit_24_39 bitb_24_39 word24_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_39 q_25_39 qb_25_39 bit_25_39 bitb_25_39 word25_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_39 q_26_39 qb_26_39 bit_26_39 bitb_26_39 word26_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_39 q_27_39 qb_27_39 bit_27_39 bitb_27_39 word27_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_39 q_28_39 qb_28_39 bit_28_39 bitb_28_39 word28_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_39 q_29_39 qb_29_39 bit_29_39 bitb_29_39 word29_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_39 q_30_39 qb_30_39 bit_30_39 bitb_30_39 word30_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_39 q_31_39 qb_31_39 bit_31_39 bitb_31_39 word31_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_39 q_32_39 qb_32_39 bit_32_39 bitb_32_39 word32_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_39 q_33_39 qb_33_39 bit_33_39 bitb_33_39 word33_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_39 q_34_39 qb_34_39 bit_34_39 bitb_34_39 word34_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_39 q_35_39 qb_35_39 bit_35_39 bitb_35_39 word35_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_39 q_36_39 qb_36_39 bit_36_39 bitb_36_39 word36_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_39 q_37_39 qb_37_39 bit_37_39 bitb_37_39 word37_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_39 q_38_39 qb_38_39 bit_38_39 bitb_38_39 word38_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_39 q_39_39 qb_39_39 bit_39_39 bitb_39_39 word39_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_39 q_40_39 qb_40_39 bit_40_39 bitb_40_39 word40_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_39 q_41_39 qb_41_39 bit_41_39 bitb_41_39 word41_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_39 q_42_39 qb_42_39 bit_42_39 bitb_42_39 word42_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_39 q_43_39 qb_43_39 bit_43_39 bitb_43_39 word43_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_39 q_44_39 qb_44_39 bit_44_39 bitb_44_39 word44_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_39 q_45_39 qb_45_39 bit_45_39 bitb_45_39 word45_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_39 q_46_39 qb_46_39 bit_46_39 bitb_46_39 word46_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_39 q_47_39 qb_47_39 bit_47_39 bitb_47_39 word47_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_39 q_48_39 qb_48_39 bit_48_39 bitb_48_39 word48_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_39 q_49_39 qb_49_39 bit_49_39 bitb_49_39 word49_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_39 q_50_39 qb_50_39 bit_50_39 bitb_50_39 word50_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_39 q_51_39 qb_51_39 bit_51_39 bitb_51_39 word51_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_39 q_52_39 qb_52_39 bit_52_39 bitb_52_39 word52_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_39 q_53_39 qb_53_39 bit_53_39 bitb_53_39 word53_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_39 q_54_39 qb_54_39 bit_54_39 bitb_54_39 word54_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_39 q_55_39 qb_55_39 bit_55_39 bitb_55_39 word55_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_39 q_56_39 qb_56_39 bit_56_39 bitb_56_39 word56_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_39 q_57_39 qb_57_39 bit_57_39 bitb_57_39 word57_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_39 q_58_39 qb_58_39 bit_58_39 bitb_58_39 word58_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_39 q_59_39 qb_59_39 bit_59_39 bitb_59_39 word59_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_39 q_60_39 qb_60_39 bit_60_39 bitb_60_39 word60_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_39 q_61_39 qb_61_39 bit_61_39 bitb_61_39 word61_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_39 q_62_39 qb_62_39 bit_62_39 bitb_62_39 word62_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_39 q_63_39 qb_63_39 bit_63_39 bitb_63_39 word63_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_39 q_64_39 qb_64_39 bit_64_39 bitb_64_39 word64_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_39 q_65_39 qb_65_39 bit_65_39 bitb_65_39 word65_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_39 q_66_39 qb_66_39 bit_66_39 bitb_66_39 word66_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_39 q_67_39 qb_67_39 bit_67_39 bitb_67_39 word67_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_39 q_68_39 qb_68_39 bit_68_39 bitb_68_39 word68_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_39 q_69_39 qb_69_39 bit_69_39 bitb_69_39 word69_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_39 q_70_39 qb_70_39 bit_70_39 bitb_70_39 word70_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_39 q_71_39 qb_71_39 bit_71_39 bitb_71_39 word71_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_39 q_72_39 qb_72_39 bit_72_39 bitb_72_39 word72_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_39 q_73_39 qb_73_39 bit_73_39 bitb_73_39 word73_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_39 q_74_39 qb_74_39 bit_74_39 bitb_74_39 word74_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_39 q_75_39 qb_75_39 bit_75_39 bitb_75_39 word75_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_39 q_76_39 qb_76_39 bit_76_39 bitb_76_39 word76_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_39 q_77_39 qb_77_39 bit_77_39 bitb_77_39 word77_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_39 q_78_39 qb_78_39 bit_78_39 bitb_78_39 word78_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_39 q_79_39 qb_79_39 bit_79_39 bitb_79_39 word79_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_39 q_80_39 qb_80_39 bit_80_39 bitb_80_39 word80_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_39 q_81_39 qb_81_39 bit_81_39 bitb_81_39 word81_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_39 q_82_39 qb_82_39 bit_82_39 bitb_82_39 word82_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_39 q_83_39 qb_83_39 bit_83_39 bitb_83_39 word83_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_39 q_84_39 qb_84_39 bit_84_39 bitb_84_39 word84_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_39 q_85_39 qb_85_39 bit_85_39 bitb_85_39 word85_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_39 q_86_39 qb_86_39 bit_86_39 bitb_86_39 word86_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_39 q_87_39 qb_87_39 bit_87_39 bitb_87_39 word87_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_39 q_88_39 qb_88_39 bit_88_39 bitb_88_39 word88_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_39 q_89_39 qb_89_39 bit_89_39 bitb_89_39 word89_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_39 q_90_39 qb_90_39 bit_90_39 bitb_90_39 word90_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_39 q_91_39 qb_91_39 bit_91_39 bitb_91_39 word91_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_39 q_92_39 qb_92_39 bit_92_39 bitb_92_39 word92_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_39 q_93_39 qb_93_39 bit_93_39 bitb_93_39 word93_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_39 q_94_39 qb_94_39 bit_94_39 bitb_94_39 word94_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_39 q_95_39 qb_95_39 bit_95_39 bitb_95_39 word95_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_39 q_96_39 qb_96_39 bit_96_39 bitb_96_39 word96_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_39 q_97_39 qb_97_39 bit_97_39 bitb_97_39 word97_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_39 q_98_39 qb_98_39 bit_98_39 bitb_98_39 word98_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_39 q_99_39 qb_99_39 bit_99_39 bitb_99_39 word99_39 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_40 q_0_40 qb_0_40 bit_0_40 bitb_0_40 word0_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_40 q_1_40 qb_1_40 bit_1_40 bitb_1_40 word1_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_40 q_2_40 qb_2_40 bit_2_40 bitb_2_40 word2_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_40 q_3_40 qb_3_40 bit_3_40 bitb_3_40 word3_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_40 q_4_40 qb_4_40 bit_4_40 bitb_4_40 word4_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_40 q_5_40 qb_5_40 bit_5_40 bitb_5_40 word5_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_40 q_6_40 qb_6_40 bit_6_40 bitb_6_40 word6_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_40 q_7_40 qb_7_40 bit_7_40 bitb_7_40 word7_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_40 q_8_40 qb_8_40 bit_8_40 bitb_8_40 word8_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_40 q_9_40 qb_9_40 bit_9_40 bitb_9_40 word9_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_40 q_10_40 qb_10_40 bit_10_40 bitb_10_40 word10_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_40 q_11_40 qb_11_40 bit_11_40 bitb_11_40 word11_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_40 q_12_40 qb_12_40 bit_12_40 bitb_12_40 word12_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_40 q_13_40 qb_13_40 bit_13_40 bitb_13_40 word13_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_40 q_14_40 qb_14_40 bit_14_40 bitb_14_40 word14_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_40 q_15_40 qb_15_40 bit_15_40 bitb_15_40 word15_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_40 q_16_40 qb_16_40 bit_16_40 bitb_16_40 word16_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_40 q_17_40 qb_17_40 bit_17_40 bitb_17_40 word17_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_40 q_18_40 qb_18_40 bit_18_40 bitb_18_40 word18_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_40 q_19_40 qb_19_40 bit_19_40 bitb_19_40 word19_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_40 q_20_40 qb_20_40 bit_20_40 bitb_20_40 word20_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_40 q_21_40 qb_21_40 bit_21_40 bitb_21_40 word21_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_40 q_22_40 qb_22_40 bit_22_40 bitb_22_40 word22_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_40 q_23_40 qb_23_40 bit_23_40 bitb_23_40 word23_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_40 q_24_40 qb_24_40 bit_24_40 bitb_24_40 word24_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_40 q_25_40 qb_25_40 bit_25_40 bitb_25_40 word25_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_40 q_26_40 qb_26_40 bit_26_40 bitb_26_40 word26_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_40 q_27_40 qb_27_40 bit_27_40 bitb_27_40 word27_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_40 q_28_40 qb_28_40 bit_28_40 bitb_28_40 word28_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_40 q_29_40 qb_29_40 bit_29_40 bitb_29_40 word29_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_40 q_30_40 qb_30_40 bit_30_40 bitb_30_40 word30_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_40 q_31_40 qb_31_40 bit_31_40 bitb_31_40 word31_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_40 q_32_40 qb_32_40 bit_32_40 bitb_32_40 word32_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_40 q_33_40 qb_33_40 bit_33_40 bitb_33_40 word33_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_40 q_34_40 qb_34_40 bit_34_40 bitb_34_40 word34_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_40 q_35_40 qb_35_40 bit_35_40 bitb_35_40 word35_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_40 q_36_40 qb_36_40 bit_36_40 bitb_36_40 word36_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_40 q_37_40 qb_37_40 bit_37_40 bitb_37_40 word37_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_40 q_38_40 qb_38_40 bit_38_40 bitb_38_40 word38_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_40 q_39_40 qb_39_40 bit_39_40 bitb_39_40 word39_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_40 q_40_40 qb_40_40 bit_40_40 bitb_40_40 word40_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_40 q_41_40 qb_41_40 bit_41_40 bitb_41_40 word41_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_40 q_42_40 qb_42_40 bit_42_40 bitb_42_40 word42_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_40 q_43_40 qb_43_40 bit_43_40 bitb_43_40 word43_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_40 q_44_40 qb_44_40 bit_44_40 bitb_44_40 word44_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_40 q_45_40 qb_45_40 bit_45_40 bitb_45_40 word45_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_40 q_46_40 qb_46_40 bit_46_40 bitb_46_40 word46_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_40 q_47_40 qb_47_40 bit_47_40 bitb_47_40 word47_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_40 q_48_40 qb_48_40 bit_48_40 bitb_48_40 word48_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_40 q_49_40 qb_49_40 bit_49_40 bitb_49_40 word49_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_40 q_50_40 qb_50_40 bit_50_40 bitb_50_40 word50_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_40 q_51_40 qb_51_40 bit_51_40 bitb_51_40 word51_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_40 q_52_40 qb_52_40 bit_52_40 bitb_52_40 word52_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_40 q_53_40 qb_53_40 bit_53_40 bitb_53_40 word53_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_40 q_54_40 qb_54_40 bit_54_40 bitb_54_40 word54_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_40 q_55_40 qb_55_40 bit_55_40 bitb_55_40 word55_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_40 q_56_40 qb_56_40 bit_56_40 bitb_56_40 word56_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_40 q_57_40 qb_57_40 bit_57_40 bitb_57_40 word57_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_40 q_58_40 qb_58_40 bit_58_40 bitb_58_40 word58_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_40 q_59_40 qb_59_40 bit_59_40 bitb_59_40 word59_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_40 q_60_40 qb_60_40 bit_60_40 bitb_60_40 word60_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_40 q_61_40 qb_61_40 bit_61_40 bitb_61_40 word61_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_40 q_62_40 qb_62_40 bit_62_40 bitb_62_40 word62_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_40 q_63_40 qb_63_40 bit_63_40 bitb_63_40 word63_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_40 q_64_40 qb_64_40 bit_64_40 bitb_64_40 word64_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_40 q_65_40 qb_65_40 bit_65_40 bitb_65_40 word65_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_40 q_66_40 qb_66_40 bit_66_40 bitb_66_40 word66_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_40 q_67_40 qb_67_40 bit_67_40 bitb_67_40 word67_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_40 q_68_40 qb_68_40 bit_68_40 bitb_68_40 word68_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_40 q_69_40 qb_69_40 bit_69_40 bitb_69_40 word69_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_40 q_70_40 qb_70_40 bit_70_40 bitb_70_40 word70_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_40 q_71_40 qb_71_40 bit_71_40 bitb_71_40 word71_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_40 q_72_40 qb_72_40 bit_72_40 bitb_72_40 word72_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_40 q_73_40 qb_73_40 bit_73_40 bitb_73_40 word73_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_40 q_74_40 qb_74_40 bit_74_40 bitb_74_40 word74_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_40 q_75_40 qb_75_40 bit_75_40 bitb_75_40 word75_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_40 q_76_40 qb_76_40 bit_76_40 bitb_76_40 word76_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_40 q_77_40 qb_77_40 bit_77_40 bitb_77_40 word77_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_40 q_78_40 qb_78_40 bit_78_40 bitb_78_40 word78_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_40 q_79_40 qb_79_40 bit_79_40 bitb_79_40 word79_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_40 q_80_40 qb_80_40 bit_80_40 bitb_80_40 word80_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_40 q_81_40 qb_81_40 bit_81_40 bitb_81_40 word81_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_40 q_82_40 qb_82_40 bit_82_40 bitb_82_40 word82_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_40 q_83_40 qb_83_40 bit_83_40 bitb_83_40 word83_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_40 q_84_40 qb_84_40 bit_84_40 bitb_84_40 word84_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_40 q_85_40 qb_85_40 bit_85_40 bitb_85_40 word85_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_40 q_86_40 qb_86_40 bit_86_40 bitb_86_40 word86_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_40 q_87_40 qb_87_40 bit_87_40 bitb_87_40 word87_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_40 q_88_40 qb_88_40 bit_88_40 bitb_88_40 word88_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_40 q_89_40 qb_89_40 bit_89_40 bitb_89_40 word89_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_40 q_90_40 qb_90_40 bit_90_40 bitb_90_40 word90_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_40 q_91_40 qb_91_40 bit_91_40 bitb_91_40 word91_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_40 q_92_40 qb_92_40 bit_92_40 bitb_92_40 word92_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_40 q_93_40 qb_93_40 bit_93_40 bitb_93_40 word93_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_40 q_94_40 qb_94_40 bit_94_40 bitb_94_40 word94_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_40 q_95_40 qb_95_40 bit_95_40 bitb_95_40 word95_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_40 q_96_40 qb_96_40 bit_96_40 bitb_96_40 word96_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_40 q_97_40 qb_97_40 bit_97_40 bitb_97_40 word97_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_40 q_98_40 qb_98_40 bit_98_40 bitb_98_40 word98_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_40 q_99_40 qb_99_40 bit_99_40 bitb_99_40 word99_40 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_41 q_0_41 qb_0_41 bit_0_41 bitb_0_41 word0_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_41 q_1_41 qb_1_41 bit_1_41 bitb_1_41 word1_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_41 q_2_41 qb_2_41 bit_2_41 bitb_2_41 word2_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_41 q_3_41 qb_3_41 bit_3_41 bitb_3_41 word3_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_41 q_4_41 qb_4_41 bit_4_41 bitb_4_41 word4_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_41 q_5_41 qb_5_41 bit_5_41 bitb_5_41 word5_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_41 q_6_41 qb_6_41 bit_6_41 bitb_6_41 word6_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_41 q_7_41 qb_7_41 bit_7_41 bitb_7_41 word7_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_41 q_8_41 qb_8_41 bit_8_41 bitb_8_41 word8_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_41 q_9_41 qb_9_41 bit_9_41 bitb_9_41 word9_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_41 q_10_41 qb_10_41 bit_10_41 bitb_10_41 word10_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_41 q_11_41 qb_11_41 bit_11_41 bitb_11_41 word11_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_41 q_12_41 qb_12_41 bit_12_41 bitb_12_41 word12_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_41 q_13_41 qb_13_41 bit_13_41 bitb_13_41 word13_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_41 q_14_41 qb_14_41 bit_14_41 bitb_14_41 word14_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_41 q_15_41 qb_15_41 bit_15_41 bitb_15_41 word15_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_41 q_16_41 qb_16_41 bit_16_41 bitb_16_41 word16_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_41 q_17_41 qb_17_41 bit_17_41 bitb_17_41 word17_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_41 q_18_41 qb_18_41 bit_18_41 bitb_18_41 word18_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_41 q_19_41 qb_19_41 bit_19_41 bitb_19_41 word19_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_41 q_20_41 qb_20_41 bit_20_41 bitb_20_41 word20_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_41 q_21_41 qb_21_41 bit_21_41 bitb_21_41 word21_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_41 q_22_41 qb_22_41 bit_22_41 bitb_22_41 word22_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_41 q_23_41 qb_23_41 bit_23_41 bitb_23_41 word23_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_41 q_24_41 qb_24_41 bit_24_41 bitb_24_41 word24_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_41 q_25_41 qb_25_41 bit_25_41 bitb_25_41 word25_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_41 q_26_41 qb_26_41 bit_26_41 bitb_26_41 word26_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_41 q_27_41 qb_27_41 bit_27_41 bitb_27_41 word27_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_41 q_28_41 qb_28_41 bit_28_41 bitb_28_41 word28_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_41 q_29_41 qb_29_41 bit_29_41 bitb_29_41 word29_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_41 q_30_41 qb_30_41 bit_30_41 bitb_30_41 word30_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_41 q_31_41 qb_31_41 bit_31_41 bitb_31_41 word31_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_41 q_32_41 qb_32_41 bit_32_41 bitb_32_41 word32_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_41 q_33_41 qb_33_41 bit_33_41 bitb_33_41 word33_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_41 q_34_41 qb_34_41 bit_34_41 bitb_34_41 word34_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_41 q_35_41 qb_35_41 bit_35_41 bitb_35_41 word35_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_41 q_36_41 qb_36_41 bit_36_41 bitb_36_41 word36_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_41 q_37_41 qb_37_41 bit_37_41 bitb_37_41 word37_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_41 q_38_41 qb_38_41 bit_38_41 bitb_38_41 word38_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_41 q_39_41 qb_39_41 bit_39_41 bitb_39_41 word39_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_41 q_40_41 qb_40_41 bit_40_41 bitb_40_41 word40_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_41 q_41_41 qb_41_41 bit_41_41 bitb_41_41 word41_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_41 q_42_41 qb_42_41 bit_42_41 bitb_42_41 word42_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_41 q_43_41 qb_43_41 bit_43_41 bitb_43_41 word43_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_41 q_44_41 qb_44_41 bit_44_41 bitb_44_41 word44_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_41 q_45_41 qb_45_41 bit_45_41 bitb_45_41 word45_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_41 q_46_41 qb_46_41 bit_46_41 bitb_46_41 word46_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_41 q_47_41 qb_47_41 bit_47_41 bitb_47_41 word47_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_41 q_48_41 qb_48_41 bit_48_41 bitb_48_41 word48_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_41 q_49_41 qb_49_41 bit_49_41 bitb_49_41 word49_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_41 q_50_41 qb_50_41 bit_50_41 bitb_50_41 word50_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_41 q_51_41 qb_51_41 bit_51_41 bitb_51_41 word51_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_41 q_52_41 qb_52_41 bit_52_41 bitb_52_41 word52_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_41 q_53_41 qb_53_41 bit_53_41 bitb_53_41 word53_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_41 q_54_41 qb_54_41 bit_54_41 bitb_54_41 word54_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_41 q_55_41 qb_55_41 bit_55_41 bitb_55_41 word55_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_41 q_56_41 qb_56_41 bit_56_41 bitb_56_41 word56_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_41 q_57_41 qb_57_41 bit_57_41 bitb_57_41 word57_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_41 q_58_41 qb_58_41 bit_58_41 bitb_58_41 word58_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_41 q_59_41 qb_59_41 bit_59_41 bitb_59_41 word59_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_41 q_60_41 qb_60_41 bit_60_41 bitb_60_41 word60_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_41 q_61_41 qb_61_41 bit_61_41 bitb_61_41 word61_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_41 q_62_41 qb_62_41 bit_62_41 bitb_62_41 word62_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_41 q_63_41 qb_63_41 bit_63_41 bitb_63_41 word63_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_41 q_64_41 qb_64_41 bit_64_41 bitb_64_41 word64_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_41 q_65_41 qb_65_41 bit_65_41 bitb_65_41 word65_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_41 q_66_41 qb_66_41 bit_66_41 bitb_66_41 word66_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_41 q_67_41 qb_67_41 bit_67_41 bitb_67_41 word67_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_41 q_68_41 qb_68_41 bit_68_41 bitb_68_41 word68_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_41 q_69_41 qb_69_41 bit_69_41 bitb_69_41 word69_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_41 q_70_41 qb_70_41 bit_70_41 bitb_70_41 word70_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_41 q_71_41 qb_71_41 bit_71_41 bitb_71_41 word71_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_41 q_72_41 qb_72_41 bit_72_41 bitb_72_41 word72_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_41 q_73_41 qb_73_41 bit_73_41 bitb_73_41 word73_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_41 q_74_41 qb_74_41 bit_74_41 bitb_74_41 word74_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_41 q_75_41 qb_75_41 bit_75_41 bitb_75_41 word75_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_41 q_76_41 qb_76_41 bit_76_41 bitb_76_41 word76_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_41 q_77_41 qb_77_41 bit_77_41 bitb_77_41 word77_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_41 q_78_41 qb_78_41 bit_78_41 bitb_78_41 word78_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_41 q_79_41 qb_79_41 bit_79_41 bitb_79_41 word79_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_41 q_80_41 qb_80_41 bit_80_41 bitb_80_41 word80_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_41 q_81_41 qb_81_41 bit_81_41 bitb_81_41 word81_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_41 q_82_41 qb_82_41 bit_82_41 bitb_82_41 word82_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_41 q_83_41 qb_83_41 bit_83_41 bitb_83_41 word83_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_41 q_84_41 qb_84_41 bit_84_41 bitb_84_41 word84_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_41 q_85_41 qb_85_41 bit_85_41 bitb_85_41 word85_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_41 q_86_41 qb_86_41 bit_86_41 bitb_86_41 word86_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_41 q_87_41 qb_87_41 bit_87_41 bitb_87_41 word87_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_41 q_88_41 qb_88_41 bit_88_41 bitb_88_41 word88_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_41 q_89_41 qb_89_41 bit_89_41 bitb_89_41 word89_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_41 q_90_41 qb_90_41 bit_90_41 bitb_90_41 word90_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_41 q_91_41 qb_91_41 bit_91_41 bitb_91_41 word91_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_41 q_92_41 qb_92_41 bit_92_41 bitb_92_41 word92_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_41 q_93_41 qb_93_41 bit_93_41 bitb_93_41 word93_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_41 q_94_41 qb_94_41 bit_94_41 bitb_94_41 word94_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_41 q_95_41 qb_95_41 bit_95_41 bitb_95_41 word95_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_41 q_96_41 qb_96_41 bit_96_41 bitb_96_41 word96_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_41 q_97_41 qb_97_41 bit_97_41 bitb_97_41 word97_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_41 q_98_41 qb_98_41 bit_98_41 bitb_98_41 word98_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_41 q_99_41 qb_99_41 bit_99_41 bitb_99_41 word99_41 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_42 q_0_42 qb_0_42 bit_0_42 bitb_0_42 word0_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_42 q_1_42 qb_1_42 bit_1_42 bitb_1_42 word1_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_42 q_2_42 qb_2_42 bit_2_42 bitb_2_42 word2_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_42 q_3_42 qb_3_42 bit_3_42 bitb_3_42 word3_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_42 q_4_42 qb_4_42 bit_4_42 bitb_4_42 word4_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_42 q_5_42 qb_5_42 bit_5_42 bitb_5_42 word5_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_42 q_6_42 qb_6_42 bit_6_42 bitb_6_42 word6_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_42 q_7_42 qb_7_42 bit_7_42 bitb_7_42 word7_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_42 q_8_42 qb_8_42 bit_8_42 bitb_8_42 word8_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_42 q_9_42 qb_9_42 bit_9_42 bitb_9_42 word9_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_42 q_10_42 qb_10_42 bit_10_42 bitb_10_42 word10_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_42 q_11_42 qb_11_42 bit_11_42 bitb_11_42 word11_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_42 q_12_42 qb_12_42 bit_12_42 bitb_12_42 word12_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_42 q_13_42 qb_13_42 bit_13_42 bitb_13_42 word13_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_42 q_14_42 qb_14_42 bit_14_42 bitb_14_42 word14_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_42 q_15_42 qb_15_42 bit_15_42 bitb_15_42 word15_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_42 q_16_42 qb_16_42 bit_16_42 bitb_16_42 word16_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_42 q_17_42 qb_17_42 bit_17_42 bitb_17_42 word17_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_42 q_18_42 qb_18_42 bit_18_42 bitb_18_42 word18_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_42 q_19_42 qb_19_42 bit_19_42 bitb_19_42 word19_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_42 q_20_42 qb_20_42 bit_20_42 bitb_20_42 word20_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_42 q_21_42 qb_21_42 bit_21_42 bitb_21_42 word21_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_42 q_22_42 qb_22_42 bit_22_42 bitb_22_42 word22_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_42 q_23_42 qb_23_42 bit_23_42 bitb_23_42 word23_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_42 q_24_42 qb_24_42 bit_24_42 bitb_24_42 word24_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_42 q_25_42 qb_25_42 bit_25_42 bitb_25_42 word25_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_42 q_26_42 qb_26_42 bit_26_42 bitb_26_42 word26_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_42 q_27_42 qb_27_42 bit_27_42 bitb_27_42 word27_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_42 q_28_42 qb_28_42 bit_28_42 bitb_28_42 word28_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_42 q_29_42 qb_29_42 bit_29_42 bitb_29_42 word29_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_42 q_30_42 qb_30_42 bit_30_42 bitb_30_42 word30_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_42 q_31_42 qb_31_42 bit_31_42 bitb_31_42 word31_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_42 q_32_42 qb_32_42 bit_32_42 bitb_32_42 word32_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_42 q_33_42 qb_33_42 bit_33_42 bitb_33_42 word33_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_42 q_34_42 qb_34_42 bit_34_42 bitb_34_42 word34_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_42 q_35_42 qb_35_42 bit_35_42 bitb_35_42 word35_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_42 q_36_42 qb_36_42 bit_36_42 bitb_36_42 word36_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_42 q_37_42 qb_37_42 bit_37_42 bitb_37_42 word37_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_42 q_38_42 qb_38_42 bit_38_42 bitb_38_42 word38_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_42 q_39_42 qb_39_42 bit_39_42 bitb_39_42 word39_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_42 q_40_42 qb_40_42 bit_40_42 bitb_40_42 word40_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_42 q_41_42 qb_41_42 bit_41_42 bitb_41_42 word41_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_42 q_42_42 qb_42_42 bit_42_42 bitb_42_42 word42_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_42 q_43_42 qb_43_42 bit_43_42 bitb_43_42 word43_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_42 q_44_42 qb_44_42 bit_44_42 bitb_44_42 word44_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_42 q_45_42 qb_45_42 bit_45_42 bitb_45_42 word45_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_42 q_46_42 qb_46_42 bit_46_42 bitb_46_42 word46_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_42 q_47_42 qb_47_42 bit_47_42 bitb_47_42 word47_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_42 q_48_42 qb_48_42 bit_48_42 bitb_48_42 word48_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_42 q_49_42 qb_49_42 bit_49_42 bitb_49_42 word49_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_42 q_50_42 qb_50_42 bit_50_42 bitb_50_42 word50_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_42 q_51_42 qb_51_42 bit_51_42 bitb_51_42 word51_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_42 q_52_42 qb_52_42 bit_52_42 bitb_52_42 word52_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_42 q_53_42 qb_53_42 bit_53_42 bitb_53_42 word53_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_42 q_54_42 qb_54_42 bit_54_42 bitb_54_42 word54_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_42 q_55_42 qb_55_42 bit_55_42 bitb_55_42 word55_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_42 q_56_42 qb_56_42 bit_56_42 bitb_56_42 word56_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_42 q_57_42 qb_57_42 bit_57_42 bitb_57_42 word57_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_42 q_58_42 qb_58_42 bit_58_42 bitb_58_42 word58_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_42 q_59_42 qb_59_42 bit_59_42 bitb_59_42 word59_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_42 q_60_42 qb_60_42 bit_60_42 bitb_60_42 word60_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_42 q_61_42 qb_61_42 bit_61_42 bitb_61_42 word61_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_42 q_62_42 qb_62_42 bit_62_42 bitb_62_42 word62_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_42 q_63_42 qb_63_42 bit_63_42 bitb_63_42 word63_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_42 q_64_42 qb_64_42 bit_64_42 bitb_64_42 word64_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_42 q_65_42 qb_65_42 bit_65_42 bitb_65_42 word65_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_42 q_66_42 qb_66_42 bit_66_42 bitb_66_42 word66_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_42 q_67_42 qb_67_42 bit_67_42 bitb_67_42 word67_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_42 q_68_42 qb_68_42 bit_68_42 bitb_68_42 word68_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_42 q_69_42 qb_69_42 bit_69_42 bitb_69_42 word69_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_42 q_70_42 qb_70_42 bit_70_42 bitb_70_42 word70_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_42 q_71_42 qb_71_42 bit_71_42 bitb_71_42 word71_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_42 q_72_42 qb_72_42 bit_72_42 bitb_72_42 word72_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_42 q_73_42 qb_73_42 bit_73_42 bitb_73_42 word73_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_42 q_74_42 qb_74_42 bit_74_42 bitb_74_42 word74_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_42 q_75_42 qb_75_42 bit_75_42 bitb_75_42 word75_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_42 q_76_42 qb_76_42 bit_76_42 bitb_76_42 word76_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_42 q_77_42 qb_77_42 bit_77_42 bitb_77_42 word77_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_42 q_78_42 qb_78_42 bit_78_42 bitb_78_42 word78_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_42 q_79_42 qb_79_42 bit_79_42 bitb_79_42 word79_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_42 q_80_42 qb_80_42 bit_80_42 bitb_80_42 word80_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_42 q_81_42 qb_81_42 bit_81_42 bitb_81_42 word81_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_42 q_82_42 qb_82_42 bit_82_42 bitb_82_42 word82_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_42 q_83_42 qb_83_42 bit_83_42 bitb_83_42 word83_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_42 q_84_42 qb_84_42 bit_84_42 bitb_84_42 word84_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_42 q_85_42 qb_85_42 bit_85_42 bitb_85_42 word85_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_42 q_86_42 qb_86_42 bit_86_42 bitb_86_42 word86_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_42 q_87_42 qb_87_42 bit_87_42 bitb_87_42 word87_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_42 q_88_42 qb_88_42 bit_88_42 bitb_88_42 word88_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_42 q_89_42 qb_89_42 bit_89_42 bitb_89_42 word89_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_42 q_90_42 qb_90_42 bit_90_42 bitb_90_42 word90_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_42 q_91_42 qb_91_42 bit_91_42 bitb_91_42 word91_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_42 q_92_42 qb_92_42 bit_92_42 bitb_92_42 word92_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_42 q_93_42 qb_93_42 bit_93_42 bitb_93_42 word93_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_42 q_94_42 qb_94_42 bit_94_42 bitb_94_42 word94_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_42 q_95_42 qb_95_42 bit_95_42 bitb_95_42 word95_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_42 q_96_42 qb_96_42 bit_96_42 bitb_96_42 word96_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_42 q_97_42 qb_97_42 bit_97_42 bitb_97_42 word97_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_42 q_98_42 qb_98_42 bit_98_42 bitb_98_42 word98_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_42 q_99_42 qb_99_42 bit_99_42 bitb_99_42 word99_42 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_43 q_0_43 qb_0_43 bit_0_43 bitb_0_43 word0_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_43 q_1_43 qb_1_43 bit_1_43 bitb_1_43 word1_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_43 q_2_43 qb_2_43 bit_2_43 bitb_2_43 word2_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_43 q_3_43 qb_3_43 bit_3_43 bitb_3_43 word3_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_43 q_4_43 qb_4_43 bit_4_43 bitb_4_43 word4_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_43 q_5_43 qb_5_43 bit_5_43 bitb_5_43 word5_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_43 q_6_43 qb_6_43 bit_6_43 bitb_6_43 word6_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_43 q_7_43 qb_7_43 bit_7_43 bitb_7_43 word7_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_43 q_8_43 qb_8_43 bit_8_43 bitb_8_43 word8_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_43 q_9_43 qb_9_43 bit_9_43 bitb_9_43 word9_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_43 q_10_43 qb_10_43 bit_10_43 bitb_10_43 word10_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_43 q_11_43 qb_11_43 bit_11_43 bitb_11_43 word11_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_43 q_12_43 qb_12_43 bit_12_43 bitb_12_43 word12_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_43 q_13_43 qb_13_43 bit_13_43 bitb_13_43 word13_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_43 q_14_43 qb_14_43 bit_14_43 bitb_14_43 word14_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_43 q_15_43 qb_15_43 bit_15_43 bitb_15_43 word15_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_43 q_16_43 qb_16_43 bit_16_43 bitb_16_43 word16_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_43 q_17_43 qb_17_43 bit_17_43 bitb_17_43 word17_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_43 q_18_43 qb_18_43 bit_18_43 bitb_18_43 word18_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_43 q_19_43 qb_19_43 bit_19_43 bitb_19_43 word19_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_43 q_20_43 qb_20_43 bit_20_43 bitb_20_43 word20_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_43 q_21_43 qb_21_43 bit_21_43 bitb_21_43 word21_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_43 q_22_43 qb_22_43 bit_22_43 bitb_22_43 word22_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_43 q_23_43 qb_23_43 bit_23_43 bitb_23_43 word23_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_43 q_24_43 qb_24_43 bit_24_43 bitb_24_43 word24_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_43 q_25_43 qb_25_43 bit_25_43 bitb_25_43 word25_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_43 q_26_43 qb_26_43 bit_26_43 bitb_26_43 word26_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_43 q_27_43 qb_27_43 bit_27_43 bitb_27_43 word27_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_43 q_28_43 qb_28_43 bit_28_43 bitb_28_43 word28_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_43 q_29_43 qb_29_43 bit_29_43 bitb_29_43 word29_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_43 q_30_43 qb_30_43 bit_30_43 bitb_30_43 word30_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_43 q_31_43 qb_31_43 bit_31_43 bitb_31_43 word31_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_43 q_32_43 qb_32_43 bit_32_43 bitb_32_43 word32_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_43 q_33_43 qb_33_43 bit_33_43 bitb_33_43 word33_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_43 q_34_43 qb_34_43 bit_34_43 bitb_34_43 word34_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_43 q_35_43 qb_35_43 bit_35_43 bitb_35_43 word35_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_43 q_36_43 qb_36_43 bit_36_43 bitb_36_43 word36_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_43 q_37_43 qb_37_43 bit_37_43 bitb_37_43 word37_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_43 q_38_43 qb_38_43 bit_38_43 bitb_38_43 word38_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_43 q_39_43 qb_39_43 bit_39_43 bitb_39_43 word39_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_43 q_40_43 qb_40_43 bit_40_43 bitb_40_43 word40_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_43 q_41_43 qb_41_43 bit_41_43 bitb_41_43 word41_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_43 q_42_43 qb_42_43 bit_42_43 bitb_42_43 word42_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_43 q_43_43 qb_43_43 bit_43_43 bitb_43_43 word43_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_43 q_44_43 qb_44_43 bit_44_43 bitb_44_43 word44_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_43 q_45_43 qb_45_43 bit_45_43 bitb_45_43 word45_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_43 q_46_43 qb_46_43 bit_46_43 bitb_46_43 word46_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_43 q_47_43 qb_47_43 bit_47_43 bitb_47_43 word47_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_43 q_48_43 qb_48_43 bit_48_43 bitb_48_43 word48_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_43 q_49_43 qb_49_43 bit_49_43 bitb_49_43 word49_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_43 q_50_43 qb_50_43 bit_50_43 bitb_50_43 word50_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_43 q_51_43 qb_51_43 bit_51_43 bitb_51_43 word51_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_43 q_52_43 qb_52_43 bit_52_43 bitb_52_43 word52_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_43 q_53_43 qb_53_43 bit_53_43 bitb_53_43 word53_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_43 q_54_43 qb_54_43 bit_54_43 bitb_54_43 word54_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_43 q_55_43 qb_55_43 bit_55_43 bitb_55_43 word55_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_43 q_56_43 qb_56_43 bit_56_43 bitb_56_43 word56_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_43 q_57_43 qb_57_43 bit_57_43 bitb_57_43 word57_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_43 q_58_43 qb_58_43 bit_58_43 bitb_58_43 word58_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_43 q_59_43 qb_59_43 bit_59_43 bitb_59_43 word59_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_43 q_60_43 qb_60_43 bit_60_43 bitb_60_43 word60_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_43 q_61_43 qb_61_43 bit_61_43 bitb_61_43 word61_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_43 q_62_43 qb_62_43 bit_62_43 bitb_62_43 word62_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_43 q_63_43 qb_63_43 bit_63_43 bitb_63_43 word63_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_43 q_64_43 qb_64_43 bit_64_43 bitb_64_43 word64_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_43 q_65_43 qb_65_43 bit_65_43 bitb_65_43 word65_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_43 q_66_43 qb_66_43 bit_66_43 bitb_66_43 word66_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_43 q_67_43 qb_67_43 bit_67_43 bitb_67_43 word67_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_43 q_68_43 qb_68_43 bit_68_43 bitb_68_43 word68_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_43 q_69_43 qb_69_43 bit_69_43 bitb_69_43 word69_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_43 q_70_43 qb_70_43 bit_70_43 bitb_70_43 word70_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_43 q_71_43 qb_71_43 bit_71_43 bitb_71_43 word71_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_43 q_72_43 qb_72_43 bit_72_43 bitb_72_43 word72_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_43 q_73_43 qb_73_43 bit_73_43 bitb_73_43 word73_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_43 q_74_43 qb_74_43 bit_74_43 bitb_74_43 word74_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_43 q_75_43 qb_75_43 bit_75_43 bitb_75_43 word75_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_43 q_76_43 qb_76_43 bit_76_43 bitb_76_43 word76_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_43 q_77_43 qb_77_43 bit_77_43 bitb_77_43 word77_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_43 q_78_43 qb_78_43 bit_78_43 bitb_78_43 word78_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_43 q_79_43 qb_79_43 bit_79_43 bitb_79_43 word79_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_43 q_80_43 qb_80_43 bit_80_43 bitb_80_43 word80_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_43 q_81_43 qb_81_43 bit_81_43 bitb_81_43 word81_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_43 q_82_43 qb_82_43 bit_82_43 bitb_82_43 word82_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_43 q_83_43 qb_83_43 bit_83_43 bitb_83_43 word83_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_43 q_84_43 qb_84_43 bit_84_43 bitb_84_43 word84_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_43 q_85_43 qb_85_43 bit_85_43 bitb_85_43 word85_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_43 q_86_43 qb_86_43 bit_86_43 bitb_86_43 word86_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_43 q_87_43 qb_87_43 bit_87_43 bitb_87_43 word87_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_43 q_88_43 qb_88_43 bit_88_43 bitb_88_43 word88_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_43 q_89_43 qb_89_43 bit_89_43 bitb_89_43 word89_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_43 q_90_43 qb_90_43 bit_90_43 bitb_90_43 word90_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_43 q_91_43 qb_91_43 bit_91_43 bitb_91_43 word91_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_43 q_92_43 qb_92_43 bit_92_43 bitb_92_43 word92_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_43 q_93_43 qb_93_43 bit_93_43 bitb_93_43 word93_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_43 q_94_43 qb_94_43 bit_94_43 bitb_94_43 word94_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_43 q_95_43 qb_95_43 bit_95_43 bitb_95_43 word95_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_43 q_96_43 qb_96_43 bit_96_43 bitb_96_43 word96_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_43 q_97_43 qb_97_43 bit_97_43 bitb_97_43 word97_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_43 q_98_43 qb_98_43 bit_98_43 bitb_98_43 word98_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_43 q_99_43 qb_99_43 bit_99_43 bitb_99_43 word99_43 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_44 q_0_44 qb_0_44 bit_0_44 bitb_0_44 word0_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_44 q_1_44 qb_1_44 bit_1_44 bitb_1_44 word1_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_44 q_2_44 qb_2_44 bit_2_44 bitb_2_44 word2_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_44 q_3_44 qb_3_44 bit_3_44 bitb_3_44 word3_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_44 q_4_44 qb_4_44 bit_4_44 bitb_4_44 word4_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_44 q_5_44 qb_5_44 bit_5_44 bitb_5_44 word5_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_44 q_6_44 qb_6_44 bit_6_44 bitb_6_44 word6_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_44 q_7_44 qb_7_44 bit_7_44 bitb_7_44 word7_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_44 q_8_44 qb_8_44 bit_8_44 bitb_8_44 word8_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_44 q_9_44 qb_9_44 bit_9_44 bitb_9_44 word9_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_44 q_10_44 qb_10_44 bit_10_44 bitb_10_44 word10_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_44 q_11_44 qb_11_44 bit_11_44 bitb_11_44 word11_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_44 q_12_44 qb_12_44 bit_12_44 bitb_12_44 word12_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_44 q_13_44 qb_13_44 bit_13_44 bitb_13_44 word13_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_44 q_14_44 qb_14_44 bit_14_44 bitb_14_44 word14_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_44 q_15_44 qb_15_44 bit_15_44 bitb_15_44 word15_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_44 q_16_44 qb_16_44 bit_16_44 bitb_16_44 word16_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_44 q_17_44 qb_17_44 bit_17_44 bitb_17_44 word17_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_44 q_18_44 qb_18_44 bit_18_44 bitb_18_44 word18_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_44 q_19_44 qb_19_44 bit_19_44 bitb_19_44 word19_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_44 q_20_44 qb_20_44 bit_20_44 bitb_20_44 word20_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_44 q_21_44 qb_21_44 bit_21_44 bitb_21_44 word21_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_44 q_22_44 qb_22_44 bit_22_44 bitb_22_44 word22_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_44 q_23_44 qb_23_44 bit_23_44 bitb_23_44 word23_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_44 q_24_44 qb_24_44 bit_24_44 bitb_24_44 word24_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_44 q_25_44 qb_25_44 bit_25_44 bitb_25_44 word25_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_44 q_26_44 qb_26_44 bit_26_44 bitb_26_44 word26_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_44 q_27_44 qb_27_44 bit_27_44 bitb_27_44 word27_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_44 q_28_44 qb_28_44 bit_28_44 bitb_28_44 word28_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_44 q_29_44 qb_29_44 bit_29_44 bitb_29_44 word29_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_44 q_30_44 qb_30_44 bit_30_44 bitb_30_44 word30_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_44 q_31_44 qb_31_44 bit_31_44 bitb_31_44 word31_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_44 q_32_44 qb_32_44 bit_32_44 bitb_32_44 word32_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_44 q_33_44 qb_33_44 bit_33_44 bitb_33_44 word33_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_44 q_34_44 qb_34_44 bit_34_44 bitb_34_44 word34_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_44 q_35_44 qb_35_44 bit_35_44 bitb_35_44 word35_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_44 q_36_44 qb_36_44 bit_36_44 bitb_36_44 word36_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_44 q_37_44 qb_37_44 bit_37_44 bitb_37_44 word37_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_44 q_38_44 qb_38_44 bit_38_44 bitb_38_44 word38_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_44 q_39_44 qb_39_44 bit_39_44 bitb_39_44 word39_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_44 q_40_44 qb_40_44 bit_40_44 bitb_40_44 word40_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_44 q_41_44 qb_41_44 bit_41_44 bitb_41_44 word41_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_44 q_42_44 qb_42_44 bit_42_44 bitb_42_44 word42_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_44 q_43_44 qb_43_44 bit_43_44 bitb_43_44 word43_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_44 q_44_44 qb_44_44 bit_44_44 bitb_44_44 word44_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_44 q_45_44 qb_45_44 bit_45_44 bitb_45_44 word45_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_44 q_46_44 qb_46_44 bit_46_44 bitb_46_44 word46_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_44 q_47_44 qb_47_44 bit_47_44 bitb_47_44 word47_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_44 q_48_44 qb_48_44 bit_48_44 bitb_48_44 word48_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_44 q_49_44 qb_49_44 bit_49_44 bitb_49_44 word49_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_44 q_50_44 qb_50_44 bit_50_44 bitb_50_44 word50_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_44 q_51_44 qb_51_44 bit_51_44 bitb_51_44 word51_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_44 q_52_44 qb_52_44 bit_52_44 bitb_52_44 word52_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_44 q_53_44 qb_53_44 bit_53_44 bitb_53_44 word53_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_44 q_54_44 qb_54_44 bit_54_44 bitb_54_44 word54_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_44 q_55_44 qb_55_44 bit_55_44 bitb_55_44 word55_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_44 q_56_44 qb_56_44 bit_56_44 bitb_56_44 word56_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_44 q_57_44 qb_57_44 bit_57_44 bitb_57_44 word57_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_44 q_58_44 qb_58_44 bit_58_44 bitb_58_44 word58_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_44 q_59_44 qb_59_44 bit_59_44 bitb_59_44 word59_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_44 q_60_44 qb_60_44 bit_60_44 bitb_60_44 word60_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_44 q_61_44 qb_61_44 bit_61_44 bitb_61_44 word61_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_44 q_62_44 qb_62_44 bit_62_44 bitb_62_44 word62_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_44 q_63_44 qb_63_44 bit_63_44 bitb_63_44 word63_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_44 q_64_44 qb_64_44 bit_64_44 bitb_64_44 word64_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_44 q_65_44 qb_65_44 bit_65_44 bitb_65_44 word65_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_44 q_66_44 qb_66_44 bit_66_44 bitb_66_44 word66_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_44 q_67_44 qb_67_44 bit_67_44 bitb_67_44 word67_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_44 q_68_44 qb_68_44 bit_68_44 bitb_68_44 word68_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_44 q_69_44 qb_69_44 bit_69_44 bitb_69_44 word69_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_44 q_70_44 qb_70_44 bit_70_44 bitb_70_44 word70_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_44 q_71_44 qb_71_44 bit_71_44 bitb_71_44 word71_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_44 q_72_44 qb_72_44 bit_72_44 bitb_72_44 word72_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_44 q_73_44 qb_73_44 bit_73_44 bitb_73_44 word73_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_44 q_74_44 qb_74_44 bit_74_44 bitb_74_44 word74_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_44 q_75_44 qb_75_44 bit_75_44 bitb_75_44 word75_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_44 q_76_44 qb_76_44 bit_76_44 bitb_76_44 word76_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_44 q_77_44 qb_77_44 bit_77_44 bitb_77_44 word77_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_44 q_78_44 qb_78_44 bit_78_44 bitb_78_44 word78_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_44 q_79_44 qb_79_44 bit_79_44 bitb_79_44 word79_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_44 q_80_44 qb_80_44 bit_80_44 bitb_80_44 word80_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_44 q_81_44 qb_81_44 bit_81_44 bitb_81_44 word81_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_44 q_82_44 qb_82_44 bit_82_44 bitb_82_44 word82_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_44 q_83_44 qb_83_44 bit_83_44 bitb_83_44 word83_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_44 q_84_44 qb_84_44 bit_84_44 bitb_84_44 word84_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_44 q_85_44 qb_85_44 bit_85_44 bitb_85_44 word85_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_44 q_86_44 qb_86_44 bit_86_44 bitb_86_44 word86_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_44 q_87_44 qb_87_44 bit_87_44 bitb_87_44 word87_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_44 q_88_44 qb_88_44 bit_88_44 bitb_88_44 word88_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_44 q_89_44 qb_89_44 bit_89_44 bitb_89_44 word89_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_44 q_90_44 qb_90_44 bit_90_44 bitb_90_44 word90_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_44 q_91_44 qb_91_44 bit_91_44 bitb_91_44 word91_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_44 q_92_44 qb_92_44 bit_92_44 bitb_92_44 word92_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_44 q_93_44 qb_93_44 bit_93_44 bitb_93_44 word93_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_44 q_94_44 qb_94_44 bit_94_44 bitb_94_44 word94_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_44 q_95_44 qb_95_44 bit_95_44 bitb_95_44 word95_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_44 q_96_44 qb_96_44 bit_96_44 bitb_96_44 word96_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_44 q_97_44 qb_97_44 bit_97_44 bitb_97_44 word97_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_44 q_98_44 qb_98_44 bit_98_44 bitb_98_44 word98_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_44 q_99_44 qb_99_44 bit_99_44 bitb_99_44 word99_44 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_45 q_0_45 qb_0_45 bit_0_45 bitb_0_45 word0_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_45 q_1_45 qb_1_45 bit_1_45 bitb_1_45 word1_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_45 q_2_45 qb_2_45 bit_2_45 bitb_2_45 word2_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_45 q_3_45 qb_3_45 bit_3_45 bitb_3_45 word3_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_45 q_4_45 qb_4_45 bit_4_45 bitb_4_45 word4_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_45 q_5_45 qb_5_45 bit_5_45 bitb_5_45 word5_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_45 q_6_45 qb_6_45 bit_6_45 bitb_6_45 word6_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_45 q_7_45 qb_7_45 bit_7_45 bitb_7_45 word7_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_45 q_8_45 qb_8_45 bit_8_45 bitb_8_45 word8_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_45 q_9_45 qb_9_45 bit_9_45 bitb_9_45 word9_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_45 q_10_45 qb_10_45 bit_10_45 bitb_10_45 word10_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_45 q_11_45 qb_11_45 bit_11_45 bitb_11_45 word11_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_45 q_12_45 qb_12_45 bit_12_45 bitb_12_45 word12_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_45 q_13_45 qb_13_45 bit_13_45 bitb_13_45 word13_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_45 q_14_45 qb_14_45 bit_14_45 bitb_14_45 word14_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_45 q_15_45 qb_15_45 bit_15_45 bitb_15_45 word15_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_45 q_16_45 qb_16_45 bit_16_45 bitb_16_45 word16_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_45 q_17_45 qb_17_45 bit_17_45 bitb_17_45 word17_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_45 q_18_45 qb_18_45 bit_18_45 bitb_18_45 word18_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_45 q_19_45 qb_19_45 bit_19_45 bitb_19_45 word19_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_45 q_20_45 qb_20_45 bit_20_45 bitb_20_45 word20_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_45 q_21_45 qb_21_45 bit_21_45 bitb_21_45 word21_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_45 q_22_45 qb_22_45 bit_22_45 bitb_22_45 word22_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_45 q_23_45 qb_23_45 bit_23_45 bitb_23_45 word23_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_45 q_24_45 qb_24_45 bit_24_45 bitb_24_45 word24_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_45 q_25_45 qb_25_45 bit_25_45 bitb_25_45 word25_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_45 q_26_45 qb_26_45 bit_26_45 bitb_26_45 word26_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_45 q_27_45 qb_27_45 bit_27_45 bitb_27_45 word27_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_45 q_28_45 qb_28_45 bit_28_45 bitb_28_45 word28_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_45 q_29_45 qb_29_45 bit_29_45 bitb_29_45 word29_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_45 q_30_45 qb_30_45 bit_30_45 bitb_30_45 word30_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_45 q_31_45 qb_31_45 bit_31_45 bitb_31_45 word31_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_45 q_32_45 qb_32_45 bit_32_45 bitb_32_45 word32_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_45 q_33_45 qb_33_45 bit_33_45 bitb_33_45 word33_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_45 q_34_45 qb_34_45 bit_34_45 bitb_34_45 word34_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_45 q_35_45 qb_35_45 bit_35_45 bitb_35_45 word35_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_45 q_36_45 qb_36_45 bit_36_45 bitb_36_45 word36_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_45 q_37_45 qb_37_45 bit_37_45 bitb_37_45 word37_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_45 q_38_45 qb_38_45 bit_38_45 bitb_38_45 word38_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_45 q_39_45 qb_39_45 bit_39_45 bitb_39_45 word39_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_45 q_40_45 qb_40_45 bit_40_45 bitb_40_45 word40_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_45 q_41_45 qb_41_45 bit_41_45 bitb_41_45 word41_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_45 q_42_45 qb_42_45 bit_42_45 bitb_42_45 word42_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_45 q_43_45 qb_43_45 bit_43_45 bitb_43_45 word43_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_45 q_44_45 qb_44_45 bit_44_45 bitb_44_45 word44_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_45 q_45_45 qb_45_45 bit_45_45 bitb_45_45 word45_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_45 q_46_45 qb_46_45 bit_46_45 bitb_46_45 word46_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_45 q_47_45 qb_47_45 bit_47_45 bitb_47_45 word47_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_45 q_48_45 qb_48_45 bit_48_45 bitb_48_45 word48_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_45 q_49_45 qb_49_45 bit_49_45 bitb_49_45 word49_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_45 q_50_45 qb_50_45 bit_50_45 bitb_50_45 word50_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_45 q_51_45 qb_51_45 bit_51_45 bitb_51_45 word51_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_45 q_52_45 qb_52_45 bit_52_45 bitb_52_45 word52_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_45 q_53_45 qb_53_45 bit_53_45 bitb_53_45 word53_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_45 q_54_45 qb_54_45 bit_54_45 bitb_54_45 word54_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_45 q_55_45 qb_55_45 bit_55_45 bitb_55_45 word55_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_45 q_56_45 qb_56_45 bit_56_45 bitb_56_45 word56_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_45 q_57_45 qb_57_45 bit_57_45 bitb_57_45 word57_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_45 q_58_45 qb_58_45 bit_58_45 bitb_58_45 word58_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_45 q_59_45 qb_59_45 bit_59_45 bitb_59_45 word59_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_45 q_60_45 qb_60_45 bit_60_45 bitb_60_45 word60_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_45 q_61_45 qb_61_45 bit_61_45 bitb_61_45 word61_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_45 q_62_45 qb_62_45 bit_62_45 bitb_62_45 word62_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_45 q_63_45 qb_63_45 bit_63_45 bitb_63_45 word63_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_45 q_64_45 qb_64_45 bit_64_45 bitb_64_45 word64_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_45 q_65_45 qb_65_45 bit_65_45 bitb_65_45 word65_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_45 q_66_45 qb_66_45 bit_66_45 bitb_66_45 word66_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_45 q_67_45 qb_67_45 bit_67_45 bitb_67_45 word67_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_45 q_68_45 qb_68_45 bit_68_45 bitb_68_45 word68_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_45 q_69_45 qb_69_45 bit_69_45 bitb_69_45 word69_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_45 q_70_45 qb_70_45 bit_70_45 bitb_70_45 word70_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_45 q_71_45 qb_71_45 bit_71_45 bitb_71_45 word71_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_45 q_72_45 qb_72_45 bit_72_45 bitb_72_45 word72_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_45 q_73_45 qb_73_45 bit_73_45 bitb_73_45 word73_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_45 q_74_45 qb_74_45 bit_74_45 bitb_74_45 word74_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_45 q_75_45 qb_75_45 bit_75_45 bitb_75_45 word75_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_45 q_76_45 qb_76_45 bit_76_45 bitb_76_45 word76_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_45 q_77_45 qb_77_45 bit_77_45 bitb_77_45 word77_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_45 q_78_45 qb_78_45 bit_78_45 bitb_78_45 word78_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_45 q_79_45 qb_79_45 bit_79_45 bitb_79_45 word79_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_45 q_80_45 qb_80_45 bit_80_45 bitb_80_45 word80_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_45 q_81_45 qb_81_45 bit_81_45 bitb_81_45 word81_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_45 q_82_45 qb_82_45 bit_82_45 bitb_82_45 word82_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_45 q_83_45 qb_83_45 bit_83_45 bitb_83_45 word83_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_45 q_84_45 qb_84_45 bit_84_45 bitb_84_45 word84_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_45 q_85_45 qb_85_45 bit_85_45 bitb_85_45 word85_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_45 q_86_45 qb_86_45 bit_86_45 bitb_86_45 word86_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_45 q_87_45 qb_87_45 bit_87_45 bitb_87_45 word87_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_45 q_88_45 qb_88_45 bit_88_45 bitb_88_45 word88_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_45 q_89_45 qb_89_45 bit_89_45 bitb_89_45 word89_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_45 q_90_45 qb_90_45 bit_90_45 bitb_90_45 word90_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_45 q_91_45 qb_91_45 bit_91_45 bitb_91_45 word91_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_45 q_92_45 qb_92_45 bit_92_45 bitb_92_45 word92_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_45 q_93_45 qb_93_45 bit_93_45 bitb_93_45 word93_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_45 q_94_45 qb_94_45 bit_94_45 bitb_94_45 word94_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_45 q_95_45 qb_95_45 bit_95_45 bitb_95_45 word95_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_45 q_96_45 qb_96_45 bit_96_45 bitb_96_45 word96_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_45 q_97_45 qb_97_45 bit_97_45 bitb_97_45 word97_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_45 q_98_45 qb_98_45 bit_98_45 bitb_98_45 word98_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_45 q_99_45 qb_99_45 bit_99_45 bitb_99_45 word99_45 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_46 q_0_46 qb_0_46 bit_0_46 bitb_0_46 word0_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_46 q_1_46 qb_1_46 bit_1_46 bitb_1_46 word1_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_46 q_2_46 qb_2_46 bit_2_46 bitb_2_46 word2_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_46 q_3_46 qb_3_46 bit_3_46 bitb_3_46 word3_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_46 q_4_46 qb_4_46 bit_4_46 bitb_4_46 word4_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_46 q_5_46 qb_5_46 bit_5_46 bitb_5_46 word5_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_46 q_6_46 qb_6_46 bit_6_46 bitb_6_46 word6_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_46 q_7_46 qb_7_46 bit_7_46 bitb_7_46 word7_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_46 q_8_46 qb_8_46 bit_8_46 bitb_8_46 word8_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_46 q_9_46 qb_9_46 bit_9_46 bitb_9_46 word9_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_46 q_10_46 qb_10_46 bit_10_46 bitb_10_46 word10_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_46 q_11_46 qb_11_46 bit_11_46 bitb_11_46 word11_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_46 q_12_46 qb_12_46 bit_12_46 bitb_12_46 word12_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_46 q_13_46 qb_13_46 bit_13_46 bitb_13_46 word13_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_46 q_14_46 qb_14_46 bit_14_46 bitb_14_46 word14_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_46 q_15_46 qb_15_46 bit_15_46 bitb_15_46 word15_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_46 q_16_46 qb_16_46 bit_16_46 bitb_16_46 word16_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_46 q_17_46 qb_17_46 bit_17_46 bitb_17_46 word17_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_46 q_18_46 qb_18_46 bit_18_46 bitb_18_46 word18_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_46 q_19_46 qb_19_46 bit_19_46 bitb_19_46 word19_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_46 q_20_46 qb_20_46 bit_20_46 bitb_20_46 word20_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_46 q_21_46 qb_21_46 bit_21_46 bitb_21_46 word21_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_46 q_22_46 qb_22_46 bit_22_46 bitb_22_46 word22_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_46 q_23_46 qb_23_46 bit_23_46 bitb_23_46 word23_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_46 q_24_46 qb_24_46 bit_24_46 bitb_24_46 word24_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_46 q_25_46 qb_25_46 bit_25_46 bitb_25_46 word25_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_46 q_26_46 qb_26_46 bit_26_46 bitb_26_46 word26_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_46 q_27_46 qb_27_46 bit_27_46 bitb_27_46 word27_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_46 q_28_46 qb_28_46 bit_28_46 bitb_28_46 word28_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_46 q_29_46 qb_29_46 bit_29_46 bitb_29_46 word29_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_46 q_30_46 qb_30_46 bit_30_46 bitb_30_46 word30_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_46 q_31_46 qb_31_46 bit_31_46 bitb_31_46 word31_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_46 q_32_46 qb_32_46 bit_32_46 bitb_32_46 word32_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_46 q_33_46 qb_33_46 bit_33_46 bitb_33_46 word33_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_46 q_34_46 qb_34_46 bit_34_46 bitb_34_46 word34_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_46 q_35_46 qb_35_46 bit_35_46 bitb_35_46 word35_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_46 q_36_46 qb_36_46 bit_36_46 bitb_36_46 word36_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_46 q_37_46 qb_37_46 bit_37_46 bitb_37_46 word37_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_46 q_38_46 qb_38_46 bit_38_46 bitb_38_46 word38_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_46 q_39_46 qb_39_46 bit_39_46 bitb_39_46 word39_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_46 q_40_46 qb_40_46 bit_40_46 bitb_40_46 word40_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_46 q_41_46 qb_41_46 bit_41_46 bitb_41_46 word41_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_46 q_42_46 qb_42_46 bit_42_46 bitb_42_46 word42_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_46 q_43_46 qb_43_46 bit_43_46 bitb_43_46 word43_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_46 q_44_46 qb_44_46 bit_44_46 bitb_44_46 word44_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_46 q_45_46 qb_45_46 bit_45_46 bitb_45_46 word45_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_46 q_46_46 qb_46_46 bit_46_46 bitb_46_46 word46_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_46 q_47_46 qb_47_46 bit_47_46 bitb_47_46 word47_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_46 q_48_46 qb_48_46 bit_48_46 bitb_48_46 word48_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_46 q_49_46 qb_49_46 bit_49_46 bitb_49_46 word49_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_46 q_50_46 qb_50_46 bit_50_46 bitb_50_46 word50_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_46 q_51_46 qb_51_46 bit_51_46 bitb_51_46 word51_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_46 q_52_46 qb_52_46 bit_52_46 bitb_52_46 word52_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_46 q_53_46 qb_53_46 bit_53_46 bitb_53_46 word53_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_46 q_54_46 qb_54_46 bit_54_46 bitb_54_46 word54_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_46 q_55_46 qb_55_46 bit_55_46 bitb_55_46 word55_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_46 q_56_46 qb_56_46 bit_56_46 bitb_56_46 word56_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_46 q_57_46 qb_57_46 bit_57_46 bitb_57_46 word57_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_46 q_58_46 qb_58_46 bit_58_46 bitb_58_46 word58_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_46 q_59_46 qb_59_46 bit_59_46 bitb_59_46 word59_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_46 q_60_46 qb_60_46 bit_60_46 bitb_60_46 word60_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_46 q_61_46 qb_61_46 bit_61_46 bitb_61_46 word61_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_46 q_62_46 qb_62_46 bit_62_46 bitb_62_46 word62_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_46 q_63_46 qb_63_46 bit_63_46 bitb_63_46 word63_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_46 q_64_46 qb_64_46 bit_64_46 bitb_64_46 word64_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_46 q_65_46 qb_65_46 bit_65_46 bitb_65_46 word65_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_46 q_66_46 qb_66_46 bit_66_46 bitb_66_46 word66_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_46 q_67_46 qb_67_46 bit_67_46 bitb_67_46 word67_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_46 q_68_46 qb_68_46 bit_68_46 bitb_68_46 word68_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_46 q_69_46 qb_69_46 bit_69_46 bitb_69_46 word69_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_46 q_70_46 qb_70_46 bit_70_46 bitb_70_46 word70_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_46 q_71_46 qb_71_46 bit_71_46 bitb_71_46 word71_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_46 q_72_46 qb_72_46 bit_72_46 bitb_72_46 word72_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_46 q_73_46 qb_73_46 bit_73_46 bitb_73_46 word73_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_46 q_74_46 qb_74_46 bit_74_46 bitb_74_46 word74_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_46 q_75_46 qb_75_46 bit_75_46 bitb_75_46 word75_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_46 q_76_46 qb_76_46 bit_76_46 bitb_76_46 word76_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_46 q_77_46 qb_77_46 bit_77_46 bitb_77_46 word77_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_46 q_78_46 qb_78_46 bit_78_46 bitb_78_46 word78_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_46 q_79_46 qb_79_46 bit_79_46 bitb_79_46 word79_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_46 q_80_46 qb_80_46 bit_80_46 bitb_80_46 word80_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_46 q_81_46 qb_81_46 bit_81_46 bitb_81_46 word81_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_46 q_82_46 qb_82_46 bit_82_46 bitb_82_46 word82_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_46 q_83_46 qb_83_46 bit_83_46 bitb_83_46 word83_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_46 q_84_46 qb_84_46 bit_84_46 bitb_84_46 word84_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_46 q_85_46 qb_85_46 bit_85_46 bitb_85_46 word85_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_46 q_86_46 qb_86_46 bit_86_46 bitb_86_46 word86_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_46 q_87_46 qb_87_46 bit_87_46 bitb_87_46 word87_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_46 q_88_46 qb_88_46 bit_88_46 bitb_88_46 word88_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_46 q_89_46 qb_89_46 bit_89_46 bitb_89_46 word89_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_46 q_90_46 qb_90_46 bit_90_46 bitb_90_46 word90_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_46 q_91_46 qb_91_46 bit_91_46 bitb_91_46 word91_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_46 q_92_46 qb_92_46 bit_92_46 bitb_92_46 word92_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_46 q_93_46 qb_93_46 bit_93_46 bitb_93_46 word93_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_46 q_94_46 qb_94_46 bit_94_46 bitb_94_46 word94_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_46 q_95_46 qb_95_46 bit_95_46 bitb_95_46 word95_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_46 q_96_46 qb_96_46 bit_96_46 bitb_96_46 word96_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_46 q_97_46 qb_97_46 bit_97_46 bitb_97_46 word97_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_46 q_98_46 qb_98_46 bit_98_46 bitb_98_46 word98_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_46 q_99_46 qb_99_46 bit_99_46 bitb_99_46 word99_46 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_47 q_0_47 qb_0_47 bit_0_47 bitb_0_47 word0_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_47 q_1_47 qb_1_47 bit_1_47 bitb_1_47 word1_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_47 q_2_47 qb_2_47 bit_2_47 bitb_2_47 word2_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_47 q_3_47 qb_3_47 bit_3_47 bitb_3_47 word3_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_47 q_4_47 qb_4_47 bit_4_47 bitb_4_47 word4_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_47 q_5_47 qb_5_47 bit_5_47 bitb_5_47 word5_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_47 q_6_47 qb_6_47 bit_6_47 bitb_6_47 word6_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_47 q_7_47 qb_7_47 bit_7_47 bitb_7_47 word7_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_47 q_8_47 qb_8_47 bit_8_47 bitb_8_47 word8_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_47 q_9_47 qb_9_47 bit_9_47 bitb_9_47 word9_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_47 q_10_47 qb_10_47 bit_10_47 bitb_10_47 word10_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_47 q_11_47 qb_11_47 bit_11_47 bitb_11_47 word11_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_47 q_12_47 qb_12_47 bit_12_47 bitb_12_47 word12_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_47 q_13_47 qb_13_47 bit_13_47 bitb_13_47 word13_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_47 q_14_47 qb_14_47 bit_14_47 bitb_14_47 word14_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_47 q_15_47 qb_15_47 bit_15_47 bitb_15_47 word15_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_47 q_16_47 qb_16_47 bit_16_47 bitb_16_47 word16_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_47 q_17_47 qb_17_47 bit_17_47 bitb_17_47 word17_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_47 q_18_47 qb_18_47 bit_18_47 bitb_18_47 word18_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_47 q_19_47 qb_19_47 bit_19_47 bitb_19_47 word19_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_47 q_20_47 qb_20_47 bit_20_47 bitb_20_47 word20_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_47 q_21_47 qb_21_47 bit_21_47 bitb_21_47 word21_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_47 q_22_47 qb_22_47 bit_22_47 bitb_22_47 word22_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_47 q_23_47 qb_23_47 bit_23_47 bitb_23_47 word23_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_47 q_24_47 qb_24_47 bit_24_47 bitb_24_47 word24_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_47 q_25_47 qb_25_47 bit_25_47 bitb_25_47 word25_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_47 q_26_47 qb_26_47 bit_26_47 bitb_26_47 word26_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_47 q_27_47 qb_27_47 bit_27_47 bitb_27_47 word27_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_47 q_28_47 qb_28_47 bit_28_47 bitb_28_47 word28_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_47 q_29_47 qb_29_47 bit_29_47 bitb_29_47 word29_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_47 q_30_47 qb_30_47 bit_30_47 bitb_30_47 word30_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_47 q_31_47 qb_31_47 bit_31_47 bitb_31_47 word31_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_47 q_32_47 qb_32_47 bit_32_47 bitb_32_47 word32_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_47 q_33_47 qb_33_47 bit_33_47 bitb_33_47 word33_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_47 q_34_47 qb_34_47 bit_34_47 bitb_34_47 word34_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_47 q_35_47 qb_35_47 bit_35_47 bitb_35_47 word35_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_47 q_36_47 qb_36_47 bit_36_47 bitb_36_47 word36_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_47 q_37_47 qb_37_47 bit_37_47 bitb_37_47 word37_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_47 q_38_47 qb_38_47 bit_38_47 bitb_38_47 word38_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_47 q_39_47 qb_39_47 bit_39_47 bitb_39_47 word39_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_47 q_40_47 qb_40_47 bit_40_47 bitb_40_47 word40_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_47 q_41_47 qb_41_47 bit_41_47 bitb_41_47 word41_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_47 q_42_47 qb_42_47 bit_42_47 bitb_42_47 word42_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_47 q_43_47 qb_43_47 bit_43_47 bitb_43_47 word43_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_47 q_44_47 qb_44_47 bit_44_47 bitb_44_47 word44_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_47 q_45_47 qb_45_47 bit_45_47 bitb_45_47 word45_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_47 q_46_47 qb_46_47 bit_46_47 bitb_46_47 word46_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_47 q_47_47 qb_47_47 bit_47_47 bitb_47_47 word47_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_47 q_48_47 qb_48_47 bit_48_47 bitb_48_47 word48_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_47 q_49_47 qb_49_47 bit_49_47 bitb_49_47 word49_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_47 q_50_47 qb_50_47 bit_50_47 bitb_50_47 word50_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_47 q_51_47 qb_51_47 bit_51_47 bitb_51_47 word51_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_47 q_52_47 qb_52_47 bit_52_47 bitb_52_47 word52_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_47 q_53_47 qb_53_47 bit_53_47 bitb_53_47 word53_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_47 q_54_47 qb_54_47 bit_54_47 bitb_54_47 word54_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_47 q_55_47 qb_55_47 bit_55_47 bitb_55_47 word55_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_47 q_56_47 qb_56_47 bit_56_47 bitb_56_47 word56_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_47 q_57_47 qb_57_47 bit_57_47 bitb_57_47 word57_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_47 q_58_47 qb_58_47 bit_58_47 bitb_58_47 word58_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_47 q_59_47 qb_59_47 bit_59_47 bitb_59_47 word59_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_47 q_60_47 qb_60_47 bit_60_47 bitb_60_47 word60_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_47 q_61_47 qb_61_47 bit_61_47 bitb_61_47 word61_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_47 q_62_47 qb_62_47 bit_62_47 bitb_62_47 word62_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_47 q_63_47 qb_63_47 bit_63_47 bitb_63_47 word63_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_47 q_64_47 qb_64_47 bit_64_47 bitb_64_47 word64_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_47 q_65_47 qb_65_47 bit_65_47 bitb_65_47 word65_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_47 q_66_47 qb_66_47 bit_66_47 bitb_66_47 word66_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_47 q_67_47 qb_67_47 bit_67_47 bitb_67_47 word67_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_47 q_68_47 qb_68_47 bit_68_47 bitb_68_47 word68_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_47 q_69_47 qb_69_47 bit_69_47 bitb_69_47 word69_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_47 q_70_47 qb_70_47 bit_70_47 bitb_70_47 word70_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_47 q_71_47 qb_71_47 bit_71_47 bitb_71_47 word71_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_47 q_72_47 qb_72_47 bit_72_47 bitb_72_47 word72_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_47 q_73_47 qb_73_47 bit_73_47 bitb_73_47 word73_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_47 q_74_47 qb_74_47 bit_74_47 bitb_74_47 word74_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_47 q_75_47 qb_75_47 bit_75_47 bitb_75_47 word75_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_47 q_76_47 qb_76_47 bit_76_47 bitb_76_47 word76_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_47 q_77_47 qb_77_47 bit_77_47 bitb_77_47 word77_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_47 q_78_47 qb_78_47 bit_78_47 bitb_78_47 word78_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_47 q_79_47 qb_79_47 bit_79_47 bitb_79_47 word79_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_47 q_80_47 qb_80_47 bit_80_47 bitb_80_47 word80_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_47 q_81_47 qb_81_47 bit_81_47 bitb_81_47 word81_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_47 q_82_47 qb_82_47 bit_82_47 bitb_82_47 word82_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_47 q_83_47 qb_83_47 bit_83_47 bitb_83_47 word83_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_47 q_84_47 qb_84_47 bit_84_47 bitb_84_47 word84_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_47 q_85_47 qb_85_47 bit_85_47 bitb_85_47 word85_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_47 q_86_47 qb_86_47 bit_86_47 bitb_86_47 word86_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_47 q_87_47 qb_87_47 bit_87_47 bitb_87_47 word87_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_47 q_88_47 qb_88_47 bit_88_47 bitb_88_47 word88_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_47 q_89_47 qb_89_47 bit_89_47 bitb_89_47 word89_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_47 q_90_47 qb_90_47 bit_90_47 bitb_90_47 word90_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_47 q_91_47 qb_91_47 bit_91_47 bitb_91_47 word91_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_47 q_92_47 qb_92_47 bit_92_47 bitb_92_47 word92_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_47 q_93_47 qb_93_47 bit_93_47 bitb_93_47 word93_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_47 q_94_47 qb_94_47 bit_94_47 bitb_94_47 word94_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_47 q_95_47 qb_95_47 bit_95_47 bitb_95_47 word95_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_47 q_96_47 qb_96_47 bit_96_47 bitb_96_47 word96_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_47 q_97_47 qb_97_47 bit_97_47 bitb_97_47 word97_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_47 q_98_47 qb_98_47 bit_98_47 bitb_98_47 word98_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_47 q_99_47 qb_99_47 bit_99_47 bitb_99_47 word99_47 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_48 q_0_48 qb_0_48 bit_0_48 bitb_0_48 word0_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_48 q_1_48 qb_1_48 bit_1_48 bitb_1_48 word1_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_48 q_2_48 qb_2_48 bit_2_48 bitb_2_48 word2_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_48 q_3_48 qb_3_48 bit_3_48 bitb_3_48 word3_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_48 q_4_48 qb_4_48 bit_4_48 bitb_4_48 word4_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_48 q_5_48 qb_5_48 bit_5_48 bitb_5_48 word5_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_48 q_6_48 qb_6_48 bit_6_48 bitb_6_48 word6_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_48 q_7_48 qb_7_48 bit_7_48 bitb_7_48 word7_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_48 q_8_48 qb_8_48 bit_8_48 bitb_8_48 word8_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_48 q_9_48 qb_9_48 bit_9_48 bitb_9_48 word9_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_48 q_10_48 qb_10_48 bit_10_48 bitb_10_48 word10_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_48 q_11_48 qb_11_48 bit_11_48 bitb_11_48 word11_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_48 q_12_48 qb_12_48 bit_12_48 bitb_12_48 word12_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_48 q_13_48 qb_13_48 bit_13_48 bitb_13_48 word13_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_48 q_14_48 qb_14_48 bit_14_48 bitb_14_48 word14_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_48 q_15_48 qb_15_48 bit_15_48 bitb_15_48 word15_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_48 q_16_48 qb_16_48 bit_16_48 bitb_16_48 word16_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_48 q_17_48 qb_17_48 bit_17_48 bitb_17_48 word17_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_48 q_18_48 qb_18_48 bit_18_48 bitb_18_48 word18_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_48 q_19_48 qb_19_48 bit_19_48 bitb_19_48 word19_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_48 q_20_48 qb_20_48 bit_20_48 bitb_20_48 word20_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_48 q_21_48 qb_21_48 bit_21_48 bitb_21_48 word21_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_48 q_22_48 qb_22_48 bit_22_48 bitb_22_48 word22_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_48 q_23_48 qb_23_48 bit_23_48 bitb_23_48 word23_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_48 q_24_48 qb_24_48 bit_24_48 bitb_24_48 word24_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_48 q_25_48 qb_25_48 bit_25_48 bitb_25_48 word25_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_48 q_26_48 qb_26_48 bit_26_48 bitb_26_48 word26_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_48 q_27_48 qb_27_48 bit_27_48 bitb_27_48 word27_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_48 q_28_48 qb_28_48 bit_28_48 bitb_28_48 word28_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_48 q_29_48 qb_29_48 bit_29_48 bitb_29_48 word29_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_48 q_30_48 qb_30_48 bit_30_48 bitb_30_48 word30_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_48 q_31_48 qb_31_48 bit_31_48 bitb_31_48 word31_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_48 q_32_48 qb_32_48 bit_32_48 bitb_32_48 word32_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_48 q_33_48 qb_33_48 bit_33_48 bitb_33_48 word33_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_48 q_34_48 qb_34_48 bit_34_48 bitb_34_48 word34_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_48 q_35_48 qb_35_48 bit_35_48 bitb_35_48 word35_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_48 q_36_48 qb_36_48 bit_36_48 bitb_36_48 word36_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_48 q_37_48 qb_37_48 bit_37_48 bitb_37_48 word37_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_48 q_38_48 qb_38_48 bit_38_48 bitb_38_48 word38_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_48 q_39_48 qb_39_48 bit_39_48 bitb_39_48 word39_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_48 q_40_48 qb_40_48 bit_40_48 bitb_40_48 word40_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_48 q_41_48 qb_41_48 bit_41_48 bitb_41_48 word41_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_48 q_42_48 qb_42_48 bit_42_48 bitb_42_48 word42_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_48 q_43_48 qb_43_48 bit_43_48 bitb_43_48 word43_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_48 q_44_48 qb_44_48 bit_44_48 bitb_44_48 word44_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_48 q_45_48 qb_45_48 bit_45_48 bitb_45_48 word45_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_48 q_46_48 qb_46_48 bit_46_48 bitb_46_48 word46_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_48 q_47_48 qb_47_48 bit_47_48 bitb_47_48 word47_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_48 q_48_48 qb_48_48 bit_48_48 bitb_48_48 word48_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_48 q_49_48 qb_49_48 bit_49_48 bitb_49_48 word49_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_48 q_50_48 qb_50_48 bit_50_48 bitb_50_48 word50_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_48 q_51_48 qb_51_48 bit_51_48 bitb_51_48 word51_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_48 q_52_48 qb_52_48 bit_52_48 bitb_52_48 word52_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_48 q_53_48 qb_53_48 bit_53_48 bitb_53_48 word53_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_48 q_54_48 qb_54_48 bit_54_48 bitb_54_48 word54_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_48 q_55_48 qb_55_48 bit_55_48 bitb_55_48 word55_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_48 q_56_48 qb_56_48 bit_56_48 bitb_56_48 word56_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_48 q_57_48 qb_57_48 bit_57_48 bitb_57_48 word57_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_48 q_58_48 qb_58_48 bit_58_48 bitb_58_48 word58_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_48 q_59_48 qb_59_48 bit_59_48 bitb_59_48 word59_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_48 q_60_48 qb_60_48 bit_60_48 bitb_60_48 word60_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_48 q_61_48 qb_61_48 bit_61_48 bitb_61_48 word61_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_48 q_62_48 qb_62_48 bit_62_48 bitb_62_48 word62_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_48 q_63_48 qb_63_48 bit_63_48 bitb_63_48 word63_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_48 q_64_48 qb_64_48 bit_64_48 bitb_64_48 word64_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_48 q_65_48 qb_65_48 bit_65_48 bitb_65_48 word65_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_48 q_66_48 qb_66_48 bit_66_48 bitb_66_48 word66_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_48 q_67_48 qb_67_48 bit_67_48 bitb_67_48 word67_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_48 q_68_48 qb_68_48 bit_68_48 bitb_68_48 word68_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_48 q_69_48 qb_69_48 bit_69_48 bitb_69_48 word69_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_48 q_70_48 qb_70_48 bit_70_48 bitb_70_48 word70_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_48 q_71_48 qb_71_48 bit_71_48 bitb_71_48 word71_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_48 q_72_48 qb_72_48 bit_72_48 bitb_72_48 word72_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_48 q_73_48 qb_73_48 bit_73_48 bitb_73_48 word73_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_48 q_74_48 qb_74_48 bit_74_48 bitb_74_48 word74_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_48 q_75_48 qb_75_48 bit_75_48 bitb_75_48 word75_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_48 q_76_48 qb_76_48 bit_76_48 bitb_76_48 word76_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_48 q_77_48 qb_77_48 bit_77_48 bitb_77_48 word77_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_48 q_78_48 qb_78_48 bit_78_48 bitb_78_48 word78_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_48 q_79_48 qb_79_48 bit_79_48 bitb_79_48 word79_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_48 q_80_48 qb_80_48 bit_80_48 bitb_80_48 word80_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_48 q_81_48 qb_81_48 bit_81_48 bitb_81_48 word81_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_48 q_82_48 qb_82_48 bit_82_48 bitb_82_48 word82_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_48 q_83_48 qb_83_48 bit_83_48 bitb_83_48 word83_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_48 q_84_48 qb_84_48 bit_84_48 bitb_84_48 word84_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_48 q_85_48 qb_85_48 bit_85_48 bitb_85_48 word85_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_48 q_86_48 qb_86_48 bit_86_48 bitb_86_48 word86_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_48 q_87_48 qb_87_48 bit_87_48 bitb_87_48 word87_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_48 q_88_48 qb_88_48 bit_88_48 bitb_88_48 word88_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_48 q_89_48 qb_89_48 bit_89_48 bitb_89_48 word89_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_48 q_90_48 qb_90_48 bit_90_48 bitb_90_48 word90_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_48 q_91_48 qb_91_48 bit_91_48 bitb_91_48 word91_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_48 q_92_48 qb_92_48 bit_92_48 bitb_92_48 word92_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_48 q_93_48 qb_93_48 bit_93_48 bitb_93_48 word93_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_48 q_94_48 qb_94_48 bit_94_48 bitb_94_48 word94_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_48 q_95_48 qb_95_48 bit_95_48 bitb_95_48 word95_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_48 q_96_48 qb_96_48 bit_96_48 bitb_96_48 word96_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_48 q_97_48 qb_97_48 bit_97_48 bitb_97_48 word97_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_48 q_98_48 qb_98_48 bit_98_48 bitb_98_48 word98_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_48 q_99_48 qb_99_48 bit_99_48 bitb_99_48 word99_48 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_49 q_0_49 qb_0_49 bit_0_49 bitb_0_49 word0_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_49 q_1_49 qb_1_49 bit_1_49 bitb_1_49 word1_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_49 q_2_49 qb_2_49 bit_2_49 bitb_2_49 word2_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_49 q_3_49 qb_3_49 bit_3_49 bitb_3_49 word3_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_49 q_4_49 qb_4_49 bit_4_49 bitb_4_49 word4_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_49 q_5_49 qb_5_49 bit_5_49 bitb_5_49 word5_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_49 q_6_49 qb_6_49 bit_6_49 bitb_6_49 word6_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_49 q_7_49 qb_7_49 bit_7_49 bitb_7_49 word7_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_49 q_8_49 qb_8_49 bit_8_49 bitb_8_49 word8_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_49 q_9_49 qb_9_49 bit_9_49 bitb_9_49 word9_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_49 q_10_49 qb_10_49 bit_10_49 bitb_10_49 word10_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_49 q_11_49 qb_11_49 bit_11_49 bitb_11_49 word11_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_49 q_12_49 qb_12_49 bit_12_49 bitb_12_49 word12_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_49 q_13_49 qb_13_49 bit_13_49 bitb_13_49 word13_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_49 q_14_49 qb_14_49 bit_14_49 bitb_14_49 word14_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_49 q_15_49 qb_15_49 bit_15_49 bitb_15_49 word15_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_49 q_16_49 qb_16_49 bit_16_49 bitb_16_49 word16_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_49 q_17_49 qb_17_49 bit_17_49 bitb_17_49 word17_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_49 q_18_49 qb_18_49 bit_18_49 bitb_18_49 word18_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_49 q_19_49 qb_19_49 bit_19_49 bitb_19_49 word19_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_49 q_20_49 qb_20_49 bit_20_49 bitb_20_49 word20_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_49 q_21_49 qb_21_49 bit_21_49 bitb_21_49 word21_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_49 q_22_49 qb_22_49 bit_22_49 bitb_22_49 word22_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_49 q_23_49 qb_23_49 bit_23_49 bitb_23_49 word23_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_49 q_24_49 qb_24_49 bit_24_49 bitb_24_49 word24_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_49 q_25_49 qb_25_49 bit_25_49 bitb_25_49 word25_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_49 q_26_49 qb_26_49 bit_26_49 bitb_26_49 word26_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_49 q_27_49 qb_27_49 bit_27_49 bitb_27_49 word27_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_49 q_28_49 qb_28_49 bit_28_49 bitb_28_49 word28_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_49 q_29_49 qb_29_49 bit_29_49 bitb_29_49 word29_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_49 q_30_49 qb_30_49 bit_30_49 bitb_30_49 word30_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_49 q_31_49 qb_31_49 bit_31_49 bitb_31_49 word31_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_49 q_32_49 qb_32_49 bit_32_49 bitb_32_49 word32_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_49 q_33_49 qb_33_49 bit_33_49 bitb_33_49 word33_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_49 q_34_49 qb_34_49 bit_34_49 bitb_34_49 word34_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_49 q_35_49 qb_35_49 bit_35_49 bitb_35_49 word35_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_49 q_36_49 qb_36_49 bit_36_49 bitb_36_49 word36_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_49 q_37_49 qb_37_49 bit_37_49 bitb_37_49 word37_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_49 q_38_49 qb_38_49 bit_38_49 bitb_38_49 word38_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_49 q_39_49 qb_39_49 bit_39_49 bitb_39_49 word39_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_49 q_40_49 qb_40_49 bit_40_49 bitb_40_49 word40_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_49 q_41_49 qb_41_49 bit_41_49 bitb_41_49 word41_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_49 q_42_49 qb_42_49 bit_42_49 bitb_42_49 word42_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_49 q_43_49 qb_43_49 bit_43_49 bitb_43_49 word43_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_49 q_44_49 qb_44_49 bit_44_49 bitb_44_49 word44_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_49 q_45_49 qb_45_49 bit_45_49 bitb_45_49 word45_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_49 q_46_49 qb_46_49 bit_46_49 bitb_46_49 word46_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_49 q_47_49 qb_47_49 bit_47_49 bitb_47_49 word47_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_49 q_48_49 qb_48_49 bit_48_49 bitb_48_49 word48_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_49 q_49_49 qb_49_49 bit_49_49 bitb_49_49 word49_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_49 q_50_49 qb_50_49 bit_50_49 bitb_50_49 word50_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_49 q_51_49 qb_51_49 bit_51_49 bitb_51_49 word51_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_49 q_52_49 qb_52_49 bit_52_49 bitb_52_49 word52_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_49 q_53_49 qb_53_49 bit_53_49 bitb_53_49 word53_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_49 q_54_49 qb_54_49 bit_54_49 bitb_54_49 word54_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_49 q_55_49 qb_55_49 bit_55_49 bitb_55_49 word55_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_49 q_56_49 qb_56_49 bit_56_49 bitb_56_49 word56_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_49 q_57_49 qb_57_49 bit_57_49 bitb_57_49 word57_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_49 q_58_49 qb_58_49 bit_58_49 bitb_58_49 word58_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_49 q_59_49 qb_59_49 bit_59_49 bitb_59_49 word59_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_49 q_60_49 qb_60_49 bit_60_49 bitb_60_49 word60_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_49 q_61_49 qb_61_49 bit_61_49 bitb_61_49 word61_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_49 q_62_49 qb_62_49 bit_62_49 bitb_62_49 word62_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_49 q_63_49 qb_63_49 bit_63_49 bitb_63_49 word63_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_49 q_64_49 qb_64_49 bit_64_49 bitb_64_49 word64_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_49 q_65_49 qb_65_49 bit_65_49 bitb_65_49 word65_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_49 q_66_49 qb_66_49 bit_66_49 bitb_66_49 word66_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_49 q_67_49 qb_67_49 bit_67_49 bitb_67_49 word67_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_49 q_68_49 qb_68_49 bit_68_49 bitb_68_49 word68_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_49 q_69_49 qb_69_49 bit_69_49 bitb_69_49 word69_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_49 q_70_49 qb_70_49 bit_70_49 bitb_70_49 word70_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_49 q_71_49 qb_71_49 bit_71_49 bitb_71_49 word71_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_49 q_72_49 qb_72_49 bit_72_49 bitb_72_49 word72_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_49 q_73_49 qb_73_49 bit_73_49 bitb_73_49 word73_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_49 q_74_49 qb_74_49 bit_74_49 bitb_74_49 word74_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_49 q_75_49 qb_75_49 bit_75_49 bitb_75_49 word75_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_49 q_76_49 qb_76_49 bit_76_49 bitb_76_49 word76_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_49 q_77_49 qb_77_49 bit_77_49 bitb_77_49 word77_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_49 q_78_49 qb_78_49 bit_78_49 bitb_78_49 word78_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_49 q_79_49 qb_79_49 bit_79_49 bitb_79_49 word79_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_49 q_80_49 qb_80_49 bit_80_49 bitb_80_49 word80_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_49 q_81_49 qb_81_49 bit_81_49 bitb_81_49 word81_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_49 q_82_49 qb_82_49 bit_82_49 bitb_82_49 word82_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_49 q_83_49 qb_83_49 bit_83_49 bitb_83_49 word83_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_49 q_84_49 qb_84_49 bit_84_49 bitb_84_49 word84_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_49 q_85_49 qb_85_49 bit_85_49 bitb_85_49 word85_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_49 q_86_49 qb_86_49 bit_86_49 bitb_86_49 word86_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_49 q_87_49 qb_87_49 bit_87_49 bitb_87_49 word87_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_49 q_88_49 qb_88_49 bit_88_49 bitb_88_49 word88_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_49 q_89_49 qb_89_49 bit_89_49 bitb_89_49 word89_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_49 q_90_49 qb_90_49 bit_90_49 bitb_90_49 word90_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_49 q_91_49 qb_91_49 bit_91_49 bitb_91_49 word91_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_49 q_92_49 qb_92_49 bit_92_49 bitb_92_49 word92_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_49 q_93_49 qb_93_49 bit_93_49 bitb_93_49 word93_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_49 q_94_49 qb_94_49 bit_94_49 bitb_94_49 word94_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_49 q_95_49 qb_95_49 bit_95_49 bitb_95_49 word95_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_49 q_96_49 qb_96_49 bit_96_49 bitb_96_49 word96_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_49 q_97_49 qb_97_49 bit_97_49 bitb_97_49 word97_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_49 q_98_49 qb_98_49 bit_98_49 bitb_98_49 word98_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_49 q_99_49 qb_99_49 bit_99_49 bitb_99_49 word99_49 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_50 q_0_50 qb_0_50 bit_0_50 bitb_0_50 word0_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_50 q_1_50 qb_1_50 bit_1_50 bitb_1_50 word1_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_50 q_2_50 qb_2_50 bit_2_50 bitb_2_50 word2_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_50 q_3_50 qb_3_50 bit_3_50 bitb_3_50 word3_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_50 q_4_50 qb_4_50 bit_4_50 bitb_4_50 word4_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_50 q_5_50 qb_5_50 bit_5_50 bitb_5_50 word5_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_50 q_6_50 qb_6_50 bit_6_50 bitb_6_50 word6_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_50 q_7_50 qb_7_50 bit_7_50 bitb_7_50 word7_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_50 q_8_50 qb_8_50 bit_8_50 bitb_8_50 word8_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_50 q_9_50 qb_9_50 bit_9_50 bitb_9_50 word9_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_50 q_10_50 qb_10_50 bit_10_50 bitb_10_50 word10_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_50 q_11_50 qb_11_50 bit_11_50 bitb_11_50 word11_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_50 q_12_50 qb_12_50 bit_12_50 bitb_12_50 word12_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_50 q_13_50 qb_13_50 bit_13_50 bitb_13_50 word13_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_50 q_14_50 qb_14_50 bit_14_50 bitb_14_50 word14_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_50 q_15_50 qb_15_50 bit_15_50 bitb_15_50 word15_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_50 q_16_50 qb_16_50 bit_16_50 bitb_16_50 word16_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_50 q_17_50 qb_17_50 bit_17_50 bitb_17_50 word17_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_50 q_18_50 qb_18_50 bit_18_50 bitb_18_50 word18_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_50 q_19_50 qb_19_50 bit_19_50 bitb_19_50 word19_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_50 q_20_50 qb_20_50 bit_20_50 bitb_20_50 word20_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_50 q_21_50 qb_21_50 bit_21_50 bitb_21_50 word21_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_50 q_22_50 qb_22_50 bit_22_50 bitb_22_50 word22_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_50 q_23_50 qb_23_50 bit_23_50 bitb_23_50 word23_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_50 q_24_50 qb_24_50 bit_24_50 bitb_24_50 word24_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_50 q_25_50 qb_25_50 bit_25_50 bitb_25_50 word25_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_50 q_26_50 qb_26_50 bit_26_50 bitb_26_50 word26_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_50 q_27_50 qb_27_50 bit_27_50 bitb_27_50 word27_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_50 q_28_50 qb_28_50 bit_28_50 bitb_28_50 word28_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_50 q_29_50 qb_29_50 bit_29_50 bitb_29_50 word29_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_50 q_30_50 qb_30_50 bit_30_50 bitb_30_50 word30_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_50 q_31_50 qb_31_50 bit_31_50 bitb_31_50 word31_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_50 q_32_50 qb_32_50 bit_32_50 bitb_32_50 word32_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_50 q_33_50 qb_33_50 bit_33_50 bitb_33_50 word33_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_50 q_34_50 qb_34_50 bit_34_50 bitb_34_50 word34_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_50 q_35_50 qb_35_50 bit_35_50 bitb_35_50 word35_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_50 q_36_50 qb_36_50 bit_36_50 bitb_36_50 word36_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_50 q_37_50 qb_37_50 bit_37_50 bitb_37_50 word37_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_50 q_38_50 qb_38_50 bit_38_50 bitb_38_50 word38_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_50 q_39_50 qb_39_50 bit_39_50 bitb_39_50 word39_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_50 q_40_50 qb_40_50 bit_40_50 bitb_40_50 word40_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_50 q_41_50 qb_41_50 bit_41_50 bitb_41_50 word41_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_50 q_42_50 qb_42_50 bit_42_50 bitb_42_50 word42_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_50 q_43_50 qb_43_50 bit_43_50 bitb_43_50 word43_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_50 q_44_50 qb_44_50 bit_44_50 bitb_44_50 word44_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_50 q_45_50 qb_45_50 bit_45_50 bitb_45_50 word45_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_50 q_46_50 qb_46_50 bit_46_50 bitb_46_50 word46_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_50 q_47_50 qb_47_50 bit_47_50 bitb_47_50 word47_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_50 q_48_50 qb_48_50 bit_48_50 bitb_48_50 word48_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_50 q_49_50 qb_49_50 bit_49_50 bitb_49_50 word49_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_50 q_50_50 qb_50_50 bit_50_50 bitb_50_50 word50_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_50 q_51_50 qb_51_50 bit_51_50 bitb_51_50 word51_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_50 q_52_50 qb_52_50 bit_52_50 bitb_52_50 word52_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_50 q_53_50 qb_53_50 bit_53_50 bitb_53_50 word53_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_50 q_54_50 qb_54_50 bit_54_50 bitb_54_50 word54_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_50 q_55_50 qb_55_50 bit_55_50 bitb_55_50 word55_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_50 q_56_50 qb_56_50 bit_56_50 bitb_56_50 word56_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_50 q_57_50 qb_57_50 bit_57_50 bitb_57_50 word57_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_50 q_58_50 qb_58_50 bit_58_50 bitb_58_50 word58_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_50 q_59_50 qb_59_50 bit_59_50 bitb_59_50 word59_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_50 q_60_50 qb_60_50 bit_60_50 bitb_60_50 word60_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_50 q_61_50 qb_61_50 bit_61_50 bitb_61_50 word61_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_50 q_62_50 qb_62_50 bit_62_50 bitb_62_50 word62_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_50 q_63_50 qb_63_50 bit_63_50 bitb_63_50 word63_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_50 q_64_50 qb_64_50 bit_64_50 bitb_64_50 word64_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_50 q_65_50 qb_65_50 bit_65_50 bitb_65_50 word65_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_50 q_66_50 qb_66_50 bit_66_50 bitb_66_50 word66_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_50 q_67_50 qb_67_50 bit_67_50 bitb_67_50 word67_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_50 q_68_50 qb_68_50 bit_68_50 bitb_68_50 word68_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_50 q_69_50 qb_69_50 bit_69_50 bitb_69_50 word69_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_50 q_70_50 qb_70_50 bit_70_50 bitb_70_50 word70_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_50 q_71_50 qb_71_50 bit_71_50 bitb_71_50 word71_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_50 q_72_50 qb_72_50 bit_72_50 bitb_72_50 word72_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_50 q_73_50 qb_73_50 bit_73_50 bitb_73_50 word73_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_50 q_74_50 qb_74_50 bit_74_50 bitb_74_50 word74_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_50 q_75_50 qb_75_50 bit_75_50 bitb_75_50 word75_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_50 q_76_50 qb_76_50 bit_76_50 bitb_76_50 word76_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_50 q_77_50 qb_77_50 bit_77_50 bitb_77_50 word77_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_50 q_78_50 qb_78_50 bit_78_50 bitb_78_50 word78_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_50 q_79_50 qb_79_50 bit_79_50 bitb_79_50 word79_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_50 q_80_50 qb_80_50 bit_80_50 bitb_80_50 word80_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_50 q_81_50 qb_81_50 bit_81_50 bitb_81_50 word81_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_50 q_82_50 qb_82_50 bit_82_50 bitb_82_50 word82_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_50 q_83_50 qb_83_50 bit_83_50 bitb_83_50 word83_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_50 q_84_50 qb_84_50 bit_84_50 bitb_84_50 word84_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_50 q_85_50 qb_85_50 bit_85_50 bitb_85_50 word85_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_50 q_86_50 qb_86_50 bit_86_50 bitb_86_50 word86_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_50 q_87_50 qb_87_50 bit_87_50 bitb_87_50 word87_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_50 q_88_50 qb_88_50 bit_88_50 bitb_88_50 word88_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_50 q_89_50 qb_89_50 bit_89_50 bitb_89_50 word89_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_50 q_90_50 qb_90_50 bit_90_50 bitb_90_50 word90_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_50 q_91_50 qb_91_50 bit_91_50 bitb_91_50 word91_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_50 q_92_50 qb_92_50 bit_92_50 bitb_92_50 word92_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_50 q_93_50 qb_93_50 bit_93_50 bitb_93_50 word93_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_50 q_94_50 qb_94_50 bit_94_50 bitb_94_50 word94_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_50 q_95_50 qb_95_50 bit_95_50 bitb_95_50 word95_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_50 q_96_50 qb_96_50 bit_96_50 bitb_96_50 word96_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_50 q_97_50 qb_97_50 bit_97_50 bitb_97_50 word97_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_50 q_98_50 qb_98_50 bit_98_50 bitb_98_50 word98_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_50 q_99_50 qb_99_50 bit_99_50 bitb_99_50 word99_50 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_51 q_0_51 qb_0_51 bit_0_51 bitb_0_51 word0_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_51 q_1_51 qb_1_51 bit_1_51 bitb_1_51 word1_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_51 q_2_51 qb_2_51 bit_2_51 bitb_2_51 word2_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_51 q_3_51 qb_3_51 bit_3_51 bitb_3_51 word3_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_51 q_4_51 qb_4_51 bit_4_51 bitb_4_51 word4_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_51 q_5_51 qb_5_51 bit_5_51 bitb_5_51 word5_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_51 q_6_51 qb_6_51 bit_6_51 bitb_6_51 word6_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_51 q_7_51 qb_7_51 bit_7_51 bitb_7_51 word7_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_51 q_8_51 qb_8_51 bit_8_51 bitb_8_51 word8_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_51 q_9_51 qb_9_51 bit_9_51 bitb_9_51 word9_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_51 q_10_51 qb_10_51 bit_10_51 bitb_10_51 word10_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_51 q_11_51 qb_11_51 bit_11_51 bitb_11_51 word11_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_51 q_12_51 qb_12_51 bit_12_51 bitb_12_51 word12_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_51 q_13_51 qb_13_51 bit_13_51 bitb_13_51 word13_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_51 q_14_51 qb_14_51 bit_14_51 bitb_14_51 word14_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_51 q_15_51 qb_15_51 bit_15_51 bitb_15_51 word15_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_51 q_16_51 qb_16_51 bit_16_51 bitb_16_51 word16_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_51 q_17_51 qb_17_51 bit_17_51 bitb_17_51 word17_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_51 q_18_51 qb_18_51 bit_18_51 bitb_18_51 word18_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_51 q_19_51 qb_19_51 bit_19_51 bitb_19_51 word19_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_51 q_20_51 qb_20_51 bit_20_51 bitb_20_51 word20_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_51 q_21_51 qb_21_51 bit_21_51 bitb_21_51 word21_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_51 q_22_51 qb_22_51 bit_22_51 bitb_22_51 word22_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_51 q_23_51 qb_23_51 bit_23_51 bitb_23_51 word23_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_51 q_24_51 qb_24_51 bit_24_51 bitb_24_51 word24_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_51 q_25_51 qb_25_51 bit_25_51 bitb_25_51 word25_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_51 q_26_51 qb_26_51 bit_26_51 bitb_26_51 word26_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_51 q_27_51 qb_27_51 bit_27_51 bitb_27_51 word27_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_51 q_28_51 qb_28_51 bit_28_51 bitb_28_51 word28_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_51 q_29_51 qb_29_51 bit_29_51 bitb_29_51 word29_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_51 q_30_51 qb_30_51 bit_30_51 bitb_30_51 word30_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_51 q_31_51 qb_31_51 bit_31_51 bitb_31_51 word31_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_51 q_32_51 qb_32_51 bit_32_51 bitb_32_51 word32_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_51 q_33_51 qb_33_51 bit_33_51 bitb_33_51 word33_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_51 q_34_51 qb_34_51 bit_34_51 bitb_34_51 word34_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_51 q_35_51 qb_35_51 bit_35_51 bitb_35_51 word35_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_51 q_36_51 qb_36_51 bit_36_51 bitb_36_51 word36_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_51 q_37_51 qb_37_51 bit_37_51 bitb_37_51 word37_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_51 q_38_51 qb_38_51 bit_38_51 bitb_38_51 word38_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_51 q_39_51 qb_39_51 bit_39_51 bitb_39_51 word39_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_51 q_40_51 qb_40_51 bit_40_51 bitb_40_51 word40_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_51 q_41_51 qb_41_51 bit_41_51 bitb_41_51 word41_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_51 q_42_51 qb_42_51 bit_42_51 bitb_42_51 word42_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_51 q_43_51 qb_43_51 bit_43_51 bitb_43_51 word43_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_51 q_44_51 qb_44_51 bit_44_51 bitb_44_51 word44_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_51 q_45_51 qb_45_51 bit_45_51 bitb_45_51 word45_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_51 q_46_51 qb_46_51 bit_46_51 bitb_46_51 word46_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_51 q_47_51 qb_47_51 bit_47_51 bitb_47_51 word47_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_51 q_48_51 qb_48_51 bit_48_51 bitb_48_51 word48_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_51 q_49_51 qb_49_51 bit_49_51 bitb_49_51 word49_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_51 q_50_51 qb_50_51 bit_50_51 bitb_50_51 word50_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_51 q_51_51 qb_51_51 bit_51_51 bitb_51_51 word51_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_51 q_52_51 qb_52_51 bit_52_51 bitb_52_51 word52_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_51 q_53_51 qb_53_51 bit_53_51 bitb_53_51 word53_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_51 q_54_51 qb_54_51 bit_54_51 bitb_54_51 word54_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_51 q_55_51 qb_55_51 bit_55_51 bitb_55_51 word55_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_51 q_56_51 qb_56_51 bit_56_51 bitb_56_51 word56_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_51 q_57_51 qb_57_51 bit_57_51 bitb_57_51 word57_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_51 q_58_51 qb_58_51 bit_58_51 bitb_58_51 word58_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_51 q_59_51 qb_59_51 bit_59_51 bitb_59_51 word59_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_51 q_60_51 qb_60_51 bit_60_51 bitb_60_51 word60_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_51 q_61_51 qb_61_51 bit_61_51 bitb_61_51 word61_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_51 q_62_51 qb_62_51 bit_62_51 bitb_62_51 word62_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_51 q_63_51 qb_63_51 bit_63_51 bitb_63_51 word63_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_51 q_64_51 qb_64_51 bit_64_51 bitb_64_51 word64_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_51 q_65_51 qb_65_51 bit_65_51 bitb_65_51 word65_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_51 q_66_51 qb_66_51 bit_66_51 bitb_66_51 word66_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_51 q_67_51 qb_67_51 bit_67_51 bitb_67_51 word67_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_51 q_68_51 qb_68_51 bit_68_51 bitb_68_51 word68_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_51 q_69_51 qb_69_51 bit_69_51 bitb_69_51 word69_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_51 q_70_51 qb_70_51 bit_70_51 bitb_70_51 word70_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_51 q_71_51 qb_71_51 bit_71_51 bitb_71_51 word71_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_51 q_72_51 qb_72_51 bit_72_51 bitb_72_51 word72_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_51 q_73_51 qb_73_51 bit_73_51 bitb_73_51 word73_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_51 q_74_51 qb_74_51 bit_74_51 bitb_74_51 word74_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_51 q_75_51 qb_75_51 bit_75_51 bitb_75_51 word75_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_51 q_76_51 qb_76_51 bit_76_51 bitb_76_51 word76_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_51 q_77_51 qb_77_51 bit_77_51 bitb_77_51 word77_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_51 q_78_51 qb_78_51 bit_78_51 bitb_78_51 word78_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_51 q_79_51 qb_79_51 bit_79_51 bitb_79_51 word79_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_51 q_80_51 qb_80_51 bit_80_51 bitb_80_51 word80_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_51 q_81_51 qb_81_51 bit_81_51 bitb_81_51 word81_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_51 q_82_51 qb_82_51 bit_82_51 bitb_82_51 word82_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_51 q_83_51 qb_83_51 bit_83_51 bitb_83_51 word83_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_51 q_84_51 qb_84_51 bit_84_51 bitb_84_51 word84_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_51 q_85_51 qb_85_51 bit_85_51 bitb_85_51 word85_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_51 q_86_51 qb_86_51 bit_86_51 bitb_86_51 word86_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_51 q_87_51 qb_87_51 bit_87_51 bitb_87_51 word87_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_51 q_88_51 qb_88_51 bit_88_51 bitb_88_51 word88_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_51 q_89_51 qb_89_51 bit_89_51 bitb_89_51 word89_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_51 q_90_51 qb_90_51 bit_90_51 bitb_90_51 word90_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_51 q_91_51 qb_91_51 bit_91_51 bitb_91_51 word91_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_51 q_92_51 qb_92_51 bit_92_51 bitb_92_51 word92_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_51 q_93_51 qb_93_51 bit_93_51 bitb_93_51 word93_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_51 q_94_51 qb_94_51 bit_94_51 bitb_94_51 word94_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_51 q_95_51 qb_95_51 bit_95_51 bitb_95_51 word95_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_51 q_96_51 qb_96_51 bit_96_51 bitb_96_51 word96_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_51 q_97_51 qb_97_51 bit_97_51 bitb_97_51 word97_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_51 q_98_51 qb_98_51 bit_98_51 bitb_98_51 word98_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_51 q_99_51 qb_99_51 bit_99_51 bitb_99_51 word99_51 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_52 q_0_52 qb_0_52 bit_0_52 bitb_0_52 word0_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_52 q_1_52 qb_1_52 bit_1_52 bitb_1_52 word1_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_52 q_2_52 qb_2_52 bit_2_52 bitb_2_52 word2_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_52 q_3_52 qb_3_52 bit_3_52 bitb_3_52 word3_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_52 q_4_52 qb_4_52 bit_4_52 bitb_4_52 word4_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_52 q_5_52 qb_5_52 bit_5_52 bitb_5_52 word5_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_52 q_6_52 qb_6_52 bit_6_52 bitb_6_52 word6_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_52 q_7_52 qb_7_52 bit_7_52 bitb_7_52 word7_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_52 q_8_52 qb_8_52 bit_8_52 bitb_8_52 word8_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_52 q_9_52 qb_9_52 bit_9_52 bitb_9_52 word9_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_52 q_10_52 qb_10_52 bit_10_52 bitb_10_52 word10_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_52 q_11_52 qb_11_52 bit_11_52 bitb_11_52 word11_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_52 q_12_52 qb_12_52 bit_12_52 bitb_12_52 word12_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_52 q_13_52 qb_13_52 bit_13_52 bitb_13_52 word13_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_52 q_14_52 qb_14_52 bit_14_52 bitb_14_52 word14_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_52 q_15_52 qb_15_52 bit_15_52 bitb_15_52 word15_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_52 q_16_52 qb_16_52 bit_16_52 bitb_16_52 word16_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_52 q_17_52 qb_17_52 bit_17_52 bitb_17_52 word17_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_52 q_18_52 qb_18_52 bit_18_52 bitb_18_52 word18_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_52 q_19_52 qb_19_52 bit_19_52 bitb_19_52 word19_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_52 q_20_52 qb_20_52 bit_20_52 bitb_20_52 word20_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_52 q_21_52 qb_21_52 bit_21_52 bitb_21_52 word21_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_52 q_22_52 qb_22_52 bit_22_52 bitb_22_52 word22_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_52 q_23_52 qb_23_52 bit_23_52 bitb_23_52 word23_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_52 q_24_52 qb_24_52 bit_24_52 bitb_24_52 word24_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_52 q_25_52 qb_25_52 bit_25_52 bitb_25_52 word25_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_52 q_26_52 qb_26_52 bit_26_52 bitb_26_52 word26_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_52 q_27_52 qb_27_52 bit_27_52 bitb_27_52 word27_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_52 q_28_52 qb_28_52 bit_28_52 bitb_28_52 word28_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_52 q_29_52 qb_29_52 bit_29_52 bitb_29_52 word29_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_52 q_30_52 qb_30_52 bit_30_52 bitb_30_52 word30_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_52 q_31_52 qb_31_52 bit_31_52 bitb_31_52 word31_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_52 q_32_52 qb_32_52 bit_32_52 bitb_32_52 word32_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_52 q_33_52 qb_33_52 bit_33_52 bitb_33_52 word33_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_52 q_34_52 qb_34_52 bit_34_52 bitb_34_52 word34_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_52 q_35_52 qb_35_52 bit_35_52 bitb_35_52 word35_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_52 q_36_52 qb_36_52 bit_36_52 bitb_36_52 word36_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_52 q_37_52 qb_37_52 bit_37_52 bitb_37_52 word37_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_52 q_38_52 qb_38_52 bit_38_52 bitb_38_52 word38_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_52 q_39_52 qb_39_52 bit_39_52 bitb_39_52 word39_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_52 q_40_52 qb_40_52 bit_40_52 bitb_40_52 word40_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_52 q_41_52 qb_41_52 bit_41_52 bitb_41_52 word41_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_52 q_42_52 qb_42_52 bit_42_52 bitb_42_52 word42_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_52 q_43_52 qb_43_52 bit_43_52 bitb_43_52 word43_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_52 q_44_52 qb_44_52 bit_44_52 bitb_44_52 word44_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_52 q_45_52 qb_45_52 bit_45_52 bitb_45_52 word45_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_52 q_46_52 qb_46_52 bit_46_52 bitb_46_52 word46_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_52 q_47_52 qb_47_52 bit_47_52 bitb_47_52 word47_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_52 q_48_52 qb_48_52 bit_48_52 bitb_48_52 word48_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_52 q_49_52 qb_49_52 bit_49_52 bitb_49_52 word49_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_52 q_50_52 qb_50_52 bit_50_52 bitb_50_52 word50_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_52 q_51_52 qb_51_52 bit_51_52 bitb_51_52 word51_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_52 q_52_52 qb_52_52 bit_52_52 bitb_52_52 word52_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_52 q_53_52 qb_53_52 bit_53_52 bitb_53_52 word53_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_52 q_54_52 qb_54_52 bit_54_52 bitb_54_52 word54_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_52 q_55_52 qb_55_52 bit_55_52 bitb_55_52 word55_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_52 q_56_52 qb_56_52 bit_56_52 bitb_56_52 word56_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_52 q_57_52 qb_57_52 bit_57_52 bitb_57_52 word57_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_52 q_58_52 qb_58_52 bit_58_52 bitb_58_52 word58_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_52 q_59_52 qb_59_52 bit_59_52 bitb_59_52 word59_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_52 q_60_52 qb_60_52 bit_60_52 bitb_60_52 word60_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_52 q_61_52 qb_61_52 bit_61_52 bitb_61_52 word61_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_52 q_62_52 qb_62_52 bit_62_52 bitb_62_52 word62_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_52 q_63_52 qb_63_52 bit_63_52 bitb_63_52 word63_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_52 q_64_52 qb_64_52 bit_64_52 bitb_64_52 word64_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_52 q_65_52 qb_65_52 bit_65_52 bitb_65_52 word65_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_52 q_66_52 qb_66_52 bit_66_52 bitb_66_52 word66_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_52 q_67_52 qb_67_52 bit_67_52 bitb_67_52 word67_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_52 q_68_52 qb_68_52 bit_68_52 bitb_68_52 word68_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_52 q_69_52 qb_69_52 bit_69_52 bitb_69_52 word69_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_52 q_70_52 qb_70_52 bit_70_52 bitb_70_52 word70_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_52 q_71_52 qb_71_52 bit_71_52 bitb_71_52 word71_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_52 q_72_52 qb_72_52 bit_72_52 bitb_72_52 word72_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_52 q_73_52 qb_73_52 bit_73_52 bitb_73_52 word73_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_52 q_74_52 qb_74_52 bit_74_52 bitb_74_52 word74_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_52 q_75_52 qb_75_52 bit_75_52 bitb_75_52 word75_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_52 q_76_52 qb_76_52 bit_76_52 bitb_76_52 word76_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_52 q_77_52 qb_77_52 bit_77_52 bitb_77_52 word77_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_52 q_78_52 qb_78_52 bit_78_52 bitb_78_52 word78_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_52 q_79_52 qb_79_52 bit_79_52 bitb_79_52 word79_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_52 q_80_52 qb_80_52 bit_80_52 bitb_80_52 word80_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_52 q_81_52 qb_81_52 bit_81_52 bitb_81_52 word81_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_52 q_82_52 qb_82_52 bit_82_52 bitb_82_52 word82_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_52 q_83_52 qb_83_52 bit_83_52 bitb_83_52 word83_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_52 q_84_52 qb_84_52 bit_84_52 bitb_84_52 word84_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_52 q_85_52 qb_85_52 bit_85_52 bitb_85_52 word85_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_52 q_86_52 qb_86_52 bit_86_52 bitb_86_52 word86_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_52 q_87_52 qb_87_52 bit_87_52 bitb_87_52 word87_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_52 q_88_52 qb_88_52 bit_88_52 bitb_88_52 word88_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_52 q_89_52 qb_89_52 bit_89_52 bitb_89_52 word89_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_52 q_90_52 qb_90_52 bit_90_52 bitb_90_52 word90_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_52 q_91_52 qb_91_52 bit_91_52 bitb_91_52 word91_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_52 q_92_52 qb_92_52 bit_92_52 bitb_92_52 word92_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_52 q_93_52 qb_93_52 bit_93_52 bitb_93_52 word93_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_52 q_94_52 qb_94_52 bit_94_52 bitb_94_52 word94_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_52 q_95_52 qb_95_52 bit_95_52 bitb_95_52 word95_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_52 q_96_52 qb_96_52 bit_96_52 bitb_96_52 word96_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_52 q_97_52 qb_97_52 bit_97_52 bitb_97_52 word97_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_52 q_98_52 qb_98_52 bit_98_52 bitb_98_52 word98_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_52 q_99_52 qb_99_52 bit_99_52 bitb_99_52 word99_52 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_53 q_0_53 qb_0_53 bit_0_53 bitb_0_53 word0_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_53 q_1_53 qb_1_53 bit_1_53 bitb_1_53 word1_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_53 q_2_53 qb_2_53 bit_2_53 bitb_2_53 word2_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_53 q_3_53 qb_3_53 bit_3_53 bitb_3_53 word3_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_53 q_4_53 qb_4_53 bit_4_53 bitb_4_53 word4_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_53 q_5_53 qb_5_53 bit_5_53 bitb_5_53 word5_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_53 q_6_53 qb_6_53 bit_6_53 bitb_6_53 word6_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_53 q_7_53 qb_7_53 bit_7_53 bitb_7_53 word7_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_53 q_8_53 qb_8_53 bit_8_53 bitb_8_53 word8_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_53 q_9_53 qb_9_53 bit_9_53 bitb_9_53 word9_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_53 q_10_53 qb_10_53 bit_10_53 bitb_10_53 word10_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_53 q_11_53 qb_11_53 bit_11_53 bitb_11_53 word11_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_53 q_12_53 qb_12_53 bit_12_53 bitb_12_53 word12_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_53 q_13_53 qb_13_53 bit_13_53 bitb_13_53 word13_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_53 q_14_53 qb_14_53 bit_14_53 bitb_14_53 word14_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_53 q_15_53 qb_15_53 bit_15_53 bitb_15_53 word15_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_53 q_16_53 qb_16_53 bit_16_53 bitb_16_53 word16_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_53 q_17_53 qb_17_53 bit_17_53 bitb_17_53 word17_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_53 q_18_53 qb_18_53 bit_18_53 bitb_18_53 word18_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_53 q_19_53 qb_19_53 bit_19_53 bitb_19_53 word19_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_53 q_20_53 qb_20_53 bit_20_53 bitb_20_53 word20_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_53 q_21_53 qb_21_53 bit_21_53 bitb_21_53 word21_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_53 q_22_53 qb_22_53 bit_22_53 bitb_22_53 word22_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_53 q_23_53 qb_23_53 bit_23_53 bitb_23_53 word23_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_53 q_24_53 qb_24_53 bit_24_53 bitb_24_53 word24_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_53 q_25_53 qb_25_53 bit_25_53 bitb_25_53 word25_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_53 q_26_53 qb_26_53 bit_26_53 bitb_26_53 word26_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_53 q_27_53 qb_27_53 bit_27_53 bitb_27_53 word27_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_53 q_28_53 qb_28_53 bit_28_53 bitb_28_53 word28_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_53 q_29_53 qb_29_53 bit_29_53 bitb_29_53 word29_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_53 q_30_53 qb_30_53 bit_30_53 bitb_30_53 word30_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_53 q_31_53 qb_31_53 bit_31_53 bitb_31_53 word31_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_53 q_32_53 qb_32_53 bit_32_53 bitb_32_53 word32_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_53 q_33_53 qb_33_53 bit_33_53 bitb_33_53 word33_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_53 q_34_53 qb_34_53 bit_34_53 bitb_34_53 word34_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_53 q_35_53 qb_35_53 bit_35_53 bitb_35_53 word35_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_53 q_36_53 qb_36_53 bit_36_53 bitb_36_53 word36_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_53 q_37_53 qb_37_53 bit_37_53 bitb_37_53 word37_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_53 q_38_53 qb_38_53 bit_38_53 bitb_38_53 word38_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_53 q_39_53 qb_39_53 bit_39_53 bitb_39_53 word39_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_53 q_40_53 qb_40_53 bit_40_53 bitb_40_53 word40_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_53 q_41_53 qb_41_53 bit_41_53 bitb_41_53 word41_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_53 q_42_53 qb_42_53 bit_42_53 bitb_42_53 word42_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_53 q_43_53 qb_43_53 bit_43_53 bitb_43_53 word43_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_53 q_44_53 qb_44_53 bit_44_53 bitb_44_53 word44_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_53 q_45_53 qb_45_53 bit_45_53 bitb_45_53 word45_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_53 q_46_53 qb_46_53 bit_46_53 bitb_46_53 word46_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_53 q_47_53 qb_47_53 bit_47_53 bitb_47_53 word47_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_53 q_48_53 qb_48_53 bit_48_53 bitb_48_53 word48_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_53 q_49_53 qb_49_53 bit_49_53 bitb_49_53 word49_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_53 q_50_53 qb_50_53 bit_50_53 bitb_50_53 word50_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_53 q_51_53 qb_51_53 bit_51_53 bitb_51_53 word51_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_53 q_52_53 qb_52_53 bit_52_53 bitb_52_53 word52_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_53 q_53_53 qb_53_53 bit_53_53 bitb_53_53 word53_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_53 q_54_53 qb_54_53 bit_54_53 bitb_54_53 word54_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_53 q_55_53 qb_55_53 bit_55_53 bitb_55_53 word55_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_53 q_56_53 qb_56_53 bit_56_53 bitb_56_53 word56_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_53 q_57_53 qb_57_53 bit_57_53 bitb_57_53 word57_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_53 q_58_53 qb_58_53 bit_58_53 bitb_58_53 word58_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_53 q_59_53 qb_59_53 bit_59_53 bitb_59_53 word59_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_53 q_60_53 qb_60_53 bit_60_53 bitb_60_53 word60_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_53 q_61_53 qb_61_53 bit_61_53 bitb_61_53 word61_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_53 q_62_53 qb_62_53 bit_62_53 bitb_62_53 word62_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_53 q_63_53 qb_63_53 bit_63_53 bitb_63_53 word63_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_53 q_64_53 qb_64_53 bit_64_53 bitb_64_53 word64_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_53 q_65_53 qb_65_53 bit_65_53 bitb_65_53 word65_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_53 q_66_53 qb_66_53 bit_66_53 bitb_66_53 word66_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_53 q_67_53 qb_67_53 bit_67_53 bitb_67_53 word67_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_53 q_68_53 qb_68_53 bit_68_53 bitb_68_53 word68_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_53 q_69_53 qb_69_53 bit_69_53 bitb_69_53 word69_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_53 q_70_53 qb_70_53 bit_70_53 bitb_70_53 word70_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_53 q_71_53 qb_71_53 bit_71_53 bitb_71_53 word71_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_53 q_72_53 qb_72_53 bit_72_53 bitb_72_53 word72_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_53 q_73_53 qb_73_53 bit_73_53 bitb_73_53 word73_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_53 q_74_53 qb_74_53 bit_74_53 bitb_74_53 word74_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_53 q_75_53 qb_75_53 bit_75_53 bitb_75_53 word75_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_53 q_76_53 qb_76_53 bit_76_53 bitb_76_53 word76_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_53 q_77_53 qb_77_53 bit_77_53 bitb_77_53 word77_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_53 q_78_53 qb_78_53 bit_78_53 bitb_78_53 word78_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_53 q_79_53 qb_79_53 bit_79_53 bitb_79_53 word79_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_53 q_80_53 qb_80_53 bit_80_53 bitb_80_53 word80_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_53 q_81_53 qb_81_53 bit_81_53 bitb_81_53 word81_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_53 q_82_53 qb_82_53 bit_82_53 bitb_82_53 word82_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_53 q_83_53 qb_83_53 bit_83_53 bitb_83_53 word83_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_53 q_84_53 qb_84_53 bit_84_53 bitb_84_53 word84_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_53 q_85_53 qb_85_53 bit_85_53 bitb_85_53 word85_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_53 q_86_53 qb_86_53 bit_86_53 bitb_86_53 word86_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_53 q_87_53 qb_87_53 bit_87_53 bitb_87_53 word87_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_53 q_88_53 qb_88_53 bit_88_53 bitb_88_53 word88_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_53 q_89_53 qb_89_53 bit_89_53 bitb_89_53 word89_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_53 q_90_53 qb_90_53 bit_90_53 bitb_90_53 word90_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_53 q_91_53 qb_91_53 bit_91_53 bitb_91_53 word91_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_53 q_92_53 qb_92_53 bit_92_53 bitb_92_53 word92_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_53 q_93_53 qb_93_53 bit_93_53 bitb_93_53 word93_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_53 q_94_53 qb_94_53 bit_94_53 bitb_94_53 word94_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_53 q_95_53 qb_95_53 bit_95_53 bitb_95_53 word95_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_53 q_96_53 qb_96_53 bit_96_53 bitb_96_53 word96_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_53 q_97_53 qb_97_53 bit_97_53 bitb_97_53 word97_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_53 q_98_53 qb_98_53 bit_98_53 bitb_98_53 word98_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_53 q_99_53 qb_99_53 bit_99_53 bitb_99_53 word99_53 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_54 q_0_54 qb_0_54 bit_0_54 bitb_0_54 word0_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_54 q_1_54 qb_1_54 bit_1_54 bitb_1_54 word1_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_54 q_2_54 qb_2_54 bit_2_54 bitb_2_54 word2_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_54 q_3_54 qb_3_54 bit_3_54 bitb_3_54 word3_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_54 q_4_54 qb_4_54 bit_4_54 bitb_4_54 word4_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_54 q_5_54 qb_5_54 bit_5_54 bitb_5_54 word5_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_54 q_6_54 qb_6_54 bit_6_54 bitb_6_54 word6_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_54 q_7_54 qb_7_54 bit_7_54 bitb_7_54 word7_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_54 q_8_54 qb_8_54 bit_8_54 bitb_8_54 word8_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_54 q_9_54 qb_9_54 bit_9_54 bitb_9_54 word9_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_54 q_10_54 qb_10_54 bit_10_54 bitb_10_54 word10_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_54 q_11_54 qb_11_54 bit_11_54 bitb_11_54 word11_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_54 q_12_54 qb_12_54 bit_12_54 bitb_12_54 word12_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_54 q_13_54 qb_13_54 bit_13_54 bitb_13_54 word13_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_54 q_14_54 qb_14_54 bit_14_54 bitb_14_54 word14_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_54 q_15_54 qb_15_54 bit_15_54 bitb_15_54 word15_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_54 q_16_54 qb_16_54 bit_16_54 bitb_16_54 word16_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_54 q_17_54 qb_17_54 bit_17_54 bitb_17_54 word17_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_54 q_18_54 qb_18_54 bit_18_54 bitb_18_54 word18_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_54 q_19_54 qb_19_54 bit_19_54 bitb_19_54 word19_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_54 q_20_54 qb_20_54 bit_20_54 bitb_20_54 word20_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_54 q_21_54 qb_21_54 bit_21_54 bitb_21_54 word21_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_54 q_22_54 qb_22_54 bit_22_54 bitb_22_54 word22_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_54 q_23_54 qb_23_54 bit_23_54 bitb_23_54 word23_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_54 q_24_54 qb_24_54 bit_24_54 bitb_24_54 word24_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_54 q_25_54 qb_25_54 bit_25_54 bitb_25_54 word25_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_54 q_26_54 qb_26_54 bit_26_54 bitb_26_54 word26_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_54 q_27_54 qb_27_54 bit_27_54 bitb_27_54 word27_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_54 q_28_54 qb_28_54 bit_28_54 bitb_28_54 word28_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_54 q_29_54 qb_29_54 bit_29_54 bitb_29_54 word29_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_54 q_30_54 qb_30_54 bit_30_54 bitb_30_54 word30_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_54 q_31_54 qb_31_54 bit_31_54 bitb_31_54 word31_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_54 q_32_54 qb_32_54 bit_32_54 bitb_32_54 word32_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_54 q_33_54 qb_33_54 bit_33_54 bitb_33_54 word33_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_54 q_34_54 qb_34_54 bit_34_54 bitb_34_54 word34_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_54 q_35_54 qb_35_54 bit_35_54 bitb_35_54 word35_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_54 q_36_54 qb_36_54 bit_36_54 bitb_36_54 word36_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_54 q_37_54 qb_37_54 bit_37_54 bitb_37_54 word37_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_54 q_38_54 qb_38_54 bit_38_54 bitb_38_54 word38_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_54 q_39_54 qb_39_54 bit_39_54 bitb_39_54 word39_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_54 q_40_54 qb_40_54 bit_40_54 bitb_40_54 word40_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_54 q_41_54 qb_41_54 bit_41_54 bitb_41_54 word41_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_54 q_42_54 qb_42_54 bit_42_54 bitb_42_54 word42_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_54 q_43_54 qb_43_54 bit_43_54 bitb_43_54 word43_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_54 q_44_54 qb_44_54 bit_44_54 bitb_44_54 word44_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_54 q_45_54 qb_45_54 bit_45_54 bitb_45_54 word45_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_54 q_46_54 qb_46_54 bit_46_54 bitb_46_54 word46_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_54 q_47_54 qb_47_54 bit_47_54 bitb_47_54 word47_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_54 q_48_54 qb_48_54 bit_48_54 bitb_48_54 word48_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_54 q_49_54 qb_49_54 bit_49_54 bitb_49_54 word49_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_54 q_50_54 qb_50_54 bit_50_54 bitb_50_54 word50_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_54 q_51_54 qb_51_54 bit_51_54 bitb_51_54 word51_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_54 q_52_54 qb_52_54 bit_52_54 bitb_52_54 word52_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_54 q_53_54 qb_53_54 bit_53_54 bitb_53_54 word53_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_54 q_54_54 qb_54_54 bit_54_54 bitb_54_54 word54_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_54 q_55_54 qb_55_54 bit_55_54 bitb_55_54 word55_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_54 q_56_54 qb_56_54 bit_56_54 bitb_56_54 word56_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_54 q_57_54 qb_57_54 bit_57_54 bitb_57_54 word57_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_54 q_58_54 qb_58_54 bit_58_54 bitb_58_54 word58_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_54 q_59_54 qb_59_54 bit_59_54 bitb_59_54 word59_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_54 q_60_54 qb_60_54 bit_60_54 bitb_60_54 word60_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_54 q_61_54 qb_61_54 bit_61_54 bitb_61_54 word61_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_54 q_62_54 qb_62_54 bit_62_54 bitb_62_54 word62_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_54 q_63_54 qb_63_54 bit_63_54 bitb_63_54 word63_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_54 q_64_54 qb_64_54 bit_64_54 bitb_64_54 word64_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_54 q_65_54 qb_65_54 bit_65_54 bitb_65_54 word65_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_54 q_66_54 qb_66_54 bit_66_54 bitb_66_54 word66_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_54 q_67_54 qb_67_54 bit_67_54 bitb_67_54 word67_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_54 q_68_54 qb_68_54 bit_68_54 bitb_68_54 word68_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_54 q_69_54 qb_69_54 bit_69_54 bitb_69_54 word69_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_54 q_70_54 qb_70_54 bit_70_54 bitb_70_54 word70_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_54 q_71_54 qb_71_54 bit_71_54 bitb_71_54 word71_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_54 q_72_54 qb_72_54 bit_72_54 bitb_72_54 word72_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_54 q_73_54 qb_73_54 bit_73_54 bitb_73_54 word73_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_54 q_74_54 qb_74_54 bit_74_54 bitb_74_54 word74_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_54 q_75_54 qb_75_54 bit_75_54 bitb_75_54 word75_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_54 q_76_54 qb_76_54 bit_76_54 bitb_76_54 word76_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_54 q_77_54 qb_77_54 bit_77_54 bitb_77_54 word77_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_54 q_78_54 qb_78_54 bit_78_54 bitb_78_54 word78_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_54 q_79_54 qb_79_54 bit_79_54 bitb_79_54 word79_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_54 q_80_54 qb_80_54 bit_80_54 bitb_80_54 word80_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_54 q_81_54 qb_81_54 bit_81_54 bitb_81_54 word81_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_54 q_82_54 qb_82_54 bit_82_54 bitb_82_54 word82_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_54 q_83_54 qb_83_54 bit_83_54 bitb_83_54 word83_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_54 q_84_54 qb_84_54 bit_84_54 bitb_84_54 word84_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_54 q_85_54 qb_85_54 bit_85_54 bitb_85_54 word85_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_54 q_86_54 qb_86_54 bit_86_54 bitb_86_54 word86_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_54 q_87_54 qb_87_54 bit_87_54 bitb_87_54 word87_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_54 q_88_54 qb_88_54 bit_88_54 bitb_88_54 word88_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_54 q_89_54 qb_89_54 bit_89_54 bitb_89_54 word89_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_54 q_90_54 qb_90_54 bit_90_54 bitb_90_54 word90_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_54 q_91_54 qb_91_54 bit_91_54 bitb_91_54 word91_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_54 q_92_54 qb_92_54 bit_92_54 bitb_92_54 word92_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_54 q_93_54 qb_93_54 bit_93_54 bitb_93_54 word93_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_54 q_94_54 qb_94_54 bit_94_54 bitb_94_54 word94_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_54 q_95_54 qb_95_54 bit_95_54 bitb_95_54 word95_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_54 q_96_54 qb_96_54 bit_96_54 bitb_96_54 word96_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_54 q_97_54 qb_97_54 bit_97_54 bitb_97_54 word97_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_54 q_98_54 qb_98_54 bit_98_54 bitb_98_54 word98_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_54 q_99_54 qb_99_54 bit_99_54 bitb_99_54 word99_54 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_55 q_0_55 qb_0_55 bit_0_55 bitb_0_55 word0_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_55 q_1_55 qb_1_55 bit_1_55 bitb_1_55 word1_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_55 q_2_55 qb_2_55 bit_2_55 bitb_2_55 word2_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_55 q_3_55 qb_3_55 bit_3_55 bitb_3_55 word3_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_55 q_4_55 qb_4_55 bit_4_55 bitb_4_55 word4_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_55 q_5_55 qb_5_55 bit_5_55 bitb_5_55 word5_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_55 q_6_55 qb_6_55 bit_6_55 bitb_6_55 word6_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_55 q_7_55 qb_7_55 bit_7_55 bitb_7_55 word7_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_55 q_8_55 qb_8_55 bit_8_55 bitb_8_55 word8_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_55 q_9_55 qb_9_55 bit_9_55 bitb_9_55 word9_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_55 q_10_55 qb_10_55 bit_10_55 bitb_10_55 word10_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_55 q_11_55 qb_11_55 bit_11_55 bitb_11_55 word11_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_55 q_12_55 qb_12_55 bit_12_55 bitb_12_55 word12_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_55 q_13_55 qb_13_55 bit_13_55 bitb_13_55 word13_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_55 q_14_55 qb_14_55 bit_14_55 bitb_14_55 word14_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_55 q_15_55 qb_15_55 bit_15_55 bitb_15_55 word15_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_55 q_16_55 qb_16_55 bit_16_55 bitb_16_55 word16_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_55 q_17_55 qb_17_55 bit_17_55 bitb_17_55 word17_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_55 q_18_55 qb_18_55 bit_18_55 bitb_18_55 word18_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_55 q_19_55 qb_19_55 bit_19_55 bitb_19_55 word19_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_55 q_20_55 qb_20_55 bit_20_55 bitb_20_55 word20_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_55 q_21_55 qb_21_55 bit_21_55 bitb_21_55 word21_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_55 q_22_55 qb_22_55 bit_22_55 bitb_22_55 word22_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_55 q_23_55 qb_23_55 bit_23_55 bitb_23_55 word23_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_55 q_24_55 qb_24_55 bit_24_55 bitb_24_55 word24_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_55 q_25_55 qb_25_55 bit_25_55 bitb_25_55 word25_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_55 q_26_55 qb_26_55 bit_26_55 bitb_26_55 word26_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_55 q_27_55 qb_27_55 bit_27_55 bitb_27_55 word27_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_55 q_28_55 qb_28_55 bit_28_55 bitb_28_55 word28_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_55 q_29_55 qb_29_55 bit_29_55 bitb_29_55 word29_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_55 q_30_55 qb_30_55 bit_30_55 bitb_30_55 word30_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_55 q_31_55 qb_31_55 bit_31_55 bitb_31_55 word31_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_55 q_32_55 qb_32_55 bit_32_55 bitb_32_55 word32_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_55 q_33_55 qb_33_55 bit_33_55 bitb_33_55 word33_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_55 q_34_55 qb_34_55 bit_34_55 bitb_34_55 word34_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_55 q_35_55 qb_35_55 bit_35_55 bitb_35_55 word35_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_55 q_36_55 qb_36_55 bit_36_55 bitb_36_55 word36_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_55 q_37_55 qb_37_55 bit_37_55 bitb_37_55 word37_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_55 q_38_55 qb_38_55 bit_38_55 bitb_38_55 word38_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_55 q_39_55 qb_39_55 bit_39_55 bitb_39_55 word39_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_55 q_40_55 qb_40_55 bit_40_55 bitb_40_55 word40_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_55 q_41_55 qb_41_55 bit_41_55 bitb_41_55 word41_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_55 q_42_55 qb_42_55 bit_42_55 bitb_42_55 word42_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_55 q_43_55 qb_43_55 bit_43_55 bitb_43_55 word43_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_55 q_44_55 qb_44_55 bit_44_55 bitb_44_55 word44_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_55 q_45_55 qb_45_55 bit_45_55 bitb_45_55 word45_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_55 q_46_55 qb_46_55 bit_46_55 bitb_46_55 word46_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_55 q_47_55 qb_47_55 bit_47_55 bitb_47_55 word47_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_55 q_48_55 qb_48_55 bit_48_55 bitb_48_55 word48_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_55 q_49_55 qb_49_55 bit_49_55 bitb_49_55 word49_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_55 q_50_55 qb_50_55 bit_50_55 bitb_50_55 word50_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_55 q_51_55 qb_51_55 bit_51_55 bitb_51_55 word51_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_55 q_52_55 qb_52_55 bit_52_55 bitb_52_55 word52_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_55 q_53_55 qb_53_55 bit_53_55 bitb_53_55 word53_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_55 q_54_55 qb_54_55 bit_54_55 bitb_54_55 word54_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_55 q_55_55 qb_55_55 bit_55_55 bitb_55_55 word55_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_55 q_56_55 qb_56_55 bit_56_55 bitb_56_55 word56_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_55 q_57_55 qb_57_55 bit_57_55 bitb_57_55 word57_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_55 q_58_55 qb_58_55 bit_58_55 bitb_58_55 word58_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_55 q_59_55 qb_59_55 bit_59_55 bitb_59_55 word59_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_55 q_60_55 qb_60_55 bit_60_55 bitb_60_55 word60_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_55 q_61_55 qb_61_55 bit_61_55 bitb_61_55 word61_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_55 q_62_55 qb_62_55 bit_62_55 bitb_62_55 word62_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_55 q_63_55 qb_63_55 bit_63_55 bitb_63_55 word63_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_55 q_64_55 qb_64_55 bit_64_55 bitb_64_55 word64_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_55 q_65_55 qb_65_55 bit_65_55 bitb_65_55 word65_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_55 q_66_55 qb_66_55 bit_66_55 bitb_66_55 word66_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_55 q_67_55 qb_67_55 bit_67_55 bitb_67_55 word67_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_55 q_68_55 qb_68_55 bit_68_55 bitb_68_55 word68_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_55 q_69_55 qb_69_55 bit_69_55 bitb_69_55 word69_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_55 q_70_55 qb_70_55 bit_70_55 bitb_70_55 word70_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_55 q_71_55 qb_71_55 bit_71_55 bitb_71_55 word71_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_55 q_72_55 qb_72_55 bit_72_55 bitb_72_55 word72_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_55 q_73_55 qb_73_55 bit_73_55 bitb_73_55 word73_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_55 q_74_55 qb_74_55 bit_74_55 bitb_74_55 word74_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_55 q_75_55 qb_75_55 bit_75_55 bitb_75_55 word75_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_55 q_76_55 qb_76_55 bit_76_55 bitb_76_55 word76_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_55 q_77_55 qb_77_55 bit_77_55 bitb_77_55 word77_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_55 q_78_55 qb_78_55 bit_78_55 bitb_78_55 word78_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_55 q_79_55 qb_79_55 bit_79_55 bitb_79_55 word79_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_55 q_80_55 qb_80_55 bit_80_55 bitb_80_55 word80_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_55 q_81_55 qb_81_55 bit_81_55 bitb_81_55 word81_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_55 q_82_55 qb_82_55 bit_82_55 bitb_82_55 word82_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_55 q_83_55 qb_83_55 bit_83_55 bitb_83_55 word83_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_55 q_84_55 qb_84_55 bit_84_55 bitb_84_55 word84_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_55 q_85_55 qb_85_55 bit_85_55 bitb_85_55 word85_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_55 q_86_55 qb_86_55 bit_86_55 bitb_86_55 word86_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_55 q_87_55 qb_87_55 bit_87_55 bitb_87_55 word87_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_55 q_88_55 qb_88_55 bit_88_55 bitb_88_55 word88_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_55 q_89_55 qb_89_55 bit_89_55 bitb_89_55 word89_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_55 q_90_55 qb_90_55 bit_90_55 bitb_90_55 word90_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_55 q_91_55 qb_91_55 bit_91_55 bitb_91_55 word91_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_55 q_92_55 qb_92_55 bit_92_55 bitb_92_55 word92_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_55 q_93_55 qb_93_55 bit_93_55 bitb_93_55 word93_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_55 q_94_55 qb_94_55 bit_94_55 bitb_94_55 word94_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_55 q_95_55 qb_95_55 bit_95_55 bitb_95_55 word95_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_55 q_96_55 qb_96_55 bit_96_55 bitb_96_55 word96_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_55 q_97_55 qb_97_55 bit_97_55 bitb_97_55 word97_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_55 q_98_55 qb_98_55 bit_98_55 bitb_98_55 word98_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_55 q_99_55 qb_99_55 bit_99_55 bitb_99_55 word99_55 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_56 q_0_56 qb_0_56 bit_0_56 bitb_0_56 word0_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_56 q_1_56 qb_1_56 bit_1_56 bitb_1_56 word1_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_56 q_2_56 qb_2_56 bit_2_56 bitb_2_56 word2_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_56 q_3_56 qb_3_56 bit_3_56 bitb_3_56 word3_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_56 q_4_56 qb_4_56 bit_4_56 bitb_4_56 word4_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_56 q_5_56 qb_5_56 bit_5_56 bitb_5_56 word5_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_56 q_6_56 qb_6_56 bit_6_56 bitb_6_56 word6_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_56 q_7_56 qb_7_56 bit_7_56 bitb_7_56 word7_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_56 q_8_56 qb_8_56 bit_8_56 bitb_8_56 word8_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_56 q_9_56 qb_9_56 bit_9_56 bitb_9_56 word9_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_56 q_10_56 qb_10_56 bit_10_56 bitb_10_56 word10_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_56 q_11_56 qb_11_56 bit_11_56 bitb_11_56 word11_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_56 q_12_56 qb_12_56 bit_12_56 bitb_12_56 word12_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_56 q_13_56 qb_13_56 bit_13_56 bitb_13_56 word13_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_56 q_14_56 qb_14_56 bit_14_56 bitb_14_56 word14_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_56 q_15_56 qb_15_56 bit_15_56 bitb_15_56 word15_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_56 q_16_56 qb_16_56 bit_16_56 bitb_16_56 word16_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_56 q_17_56 qb_17_56 bit_17_56 bitb_17_56 word17_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_56 q_18_56 qb_18_56 bit_18_56 bitb_18_56 word18_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_56 q_19_56 qb_19_56 bit_19_56 bitb_19_56 word19_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_56 q_20_56 qb_20_56 bit_20_56 bitb_20_56 word20_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_56 q_21_56 qb_21_56 bit_21_56 bitb_21_56 word21_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_56 q_22_56 qb_22_56 bit_22_56 bitb_22_56 word22_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_56 q_23_56 qb_23_56 bit_23_56 bitb_23_56 word23_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_56 q_24_56 qb_24_56 bit_24_56 bitb_24_56 word24_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_56 q_25_56 qb_25_56 bit_25_56 bitb_25_56 word25_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_56 q_26_56 qb_26_56 bit_26_56 bitb_26_56 word26_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_56 q_27_56 qb_27_56 bit_27_56 bitb_27_56 word27_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_56 q_28_56 qb_28_56 bit_28_56 bitb_28_56 word28_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_56 q_29_56 qb_29_56 bit_29_56 bitb_29_56 word29_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_56 q_30_56 qb_30_56 bit_30_56 bitb_30_56 word30_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_56 q_31_56 qb_31_56 bit_31_56 bitb_31_56 word31_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_56 q_32_56 qb_32_56 bit_32_56 bitb_32_56 word32_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_56 q_33_56 qb_33_56 bit_33_56 bitb_33_56 word33_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_56 q_34_56 qb_34_56 bit_34_56 bitb_34_56 word34_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_56 q_35_56 qb_35_56 bit_35_56 bitb_35_56 word35_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_56 q_36_56 qb_36_56 bit_36_56 bitb_36_56 word36_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_56 q_37_56 qb_37_56 bit_37_56 bitb_37_56 word37_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_56 q_38_56 qb_38_56 bit_38_56 bitb_38_56 word38_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_56 q_39_56 qb_39_56 bit_39_56 bitb_39_56 word39_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_56 q_40_56 qb_40_56 bit_40_56 bitb_40_56 word40_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_56 q_41_56 qb_41_56 bit_41_56 bitb_41_56 word41_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_56 q_42_56 qb_42_56 bit_42_56 bitb_42_56 word42_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_56 q_43_56 qb_43_56 bit_43_56 bitb_43_56 word43_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_56 q_44_56 qb_44_56 bit_44_56 bitb_44_56 word44_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_56 q_45_56 qb_45_56 bit_45_56 bitb_45_56 word45_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_56 q_46_56 qb_46_56 bit_46_56 bitb_46_56 word46_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_56 q_47_56 qb_47_56 bit_47_56 bitb_47_56 word47_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_56 q_48_56 qb_48_56 bit_48_56 bitb_48_56 word48_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_56 q_49_56 qb_49_56 bit_49_56 bitb_49_56 word49_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_56 q_50_56 qb_50_56 bit_50_56 bitb_50_56 word50_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_56 q_51_56 qb_51_56 bit_51_56 bitb_51_56 word51_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_56 q_52_56 qb_52_56 bit_52_56 bitb_52_56 word52_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_56 q_53_56 qb_53_56 bit_53_56 bitb_53_56 word53_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_56 q_54_56 qb_54_56 bit_54_56 bitb_54_56 word54_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_56 q_55_56 qb_55_56 bit_55_56 bitb_55_56 word55_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_56 q_56_56 qb_56_56 bit_56_56 bitb_56_56 word56_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_56 q_57_56 qb_57_56 bit_57_56 bitb_57_56 word57_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_56 q_58_56 qb_58_56 bit_58_56 bitb_58_56 word58_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_56 q_59_56 qb_59_56 bit_59_56 bitb_59_56 word59_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_56 q_60_56 qb_60_56 bit_60_56 bitb_60_56 word60_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_56 q_61_56 qb_61_56 bit_61_56 bitb_61_56 word61_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_56 q_62_56 qb_62_56 bit_62_56 bitb_62_56 word62_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_56 q_63_56 qb_63_56 bit_63_56 bitb_63_56 word63_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_56 q_64_56 qb_64_56 bit_64_56 bitb_64_56 word64_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_56 q_65_56 qb_65_56 bit_65_56 bitb_65_56 word65_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_56 q_66_56 qb_66_56 bit_66_56 bitb_66_56 word66_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_56 q_67_56 qb_67_56 bit_67_56 bitb_67_56 word67_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_56 q_68_56 qb_68_56 bit_68_56 bitb_68_56 word68_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_56 q_69_56 qb_69_56 bit_69_56 bitb_69_56 word69_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_56 q_70_56 qb_70_56 bit_70_56 bitb_70_56 word70_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_56 q_71_56 qb_71_56 bit_71_56 bitb_71_56 word71_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_56 q_72_56 qb_72_56 bit_72_56 bitb_72_56 word72_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_56 q_73_56 qb_73_56 bit_73_56 bitb_73_56 word73_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_56 q_74_56 qb_74_56 bit_74_56 bitb_74_56 word74_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_56 q_75_56 qb_75_56 bit_75_56 bitb_75_56 word75_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_56 q_76_56 qb_76_56 bit_76_56 bitb_76_56 word76_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_56 q_77_56 qb_77_56 bit_77_56 bitb_77_56 word77_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_56 q_78_56 qb_78_56 bit_78_56 bitb_78_56 word78_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_56 q_79_56 qb_79_56 bit_79_56 bitb_79_56 word79_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_56 q_80_56 qb_80_56 bit_80_56 bitb_80_56 word80_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_56 q_81_56 qb_81_56 bit_81_56 bitb_81_56 word81_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_56 q_82_56 qb_82_56 bit_82_56 bitb_82_56 word82_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_56 q_83_56 qb_83_56 bit_83_56 bitb_83_56 word83_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_56 q_84_56 qb_84_56 bit_84_56 bitb_84_56 word84_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_56 q_85_56 qb_85_56 bit_85_56 bitb_85_56 word85_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_56 q_86_56 qb_86_56 bit_86_56 bitb_86_56 word86_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_56 q_87_56 qb_87_56 bit_87_56 bitb_87_56 word87_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_56 q_88_56 qb_88_56 bit_88_56 bitb_88_56 word88_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_56 q_89_56 qb_89_56 bit_89_56 bitb_89_56 word89_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_56 q_90_56 qb_90_56 bit_90_56 bitb_90_56 word90_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_56 q_91_56 qb_91_56 bit_91_56 bitb_91_56 word91_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_56 q_92_56 qb_92_56 bit_92_56 bitb_92_56 word92_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_56 q_93_56 qb_93_56 bit_93_56 bitb_93_56 word93_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_56 q_94_56 qb_94_56 bit_94_56 bitb_94_56 word94_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_56 q_95_56 qb_95_56 bit_95_56 bitb_95_56 word95_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_56 q_96_56 qb_96_56 bit_96_56 bitb_96_56 word96_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_56 q_97_56 qb_97_56 bit_97_56 bitb_97_56 word97_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_56 q_98_56 qb_98_56 bit_98_56 bitb_98_56 word98_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_56 q_99_56 qb_99_56 bit_99_56 bitb_99_56 word99_56 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_57 q_0_57 qb_0_57 bit_0_57 bitb_0_57 word0_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_57 q_1_57 qb_1_57 bit_1_57 bitb_1_57 word1_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_57 q_2_57 qb_2_57 bit_2_57 bitb_2_57 word2_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_57 q_3_57 qb_3_57 bit_3_57 bitb_3_57 word3_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_57 q_4_57 qb_4_57 bit_4_57 bitb_4_57 word4_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_57 q_5_57 qb_5_57 bit_5_57 bitb_5_57 word5_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_57 q_6_57 qb_6_57 bit_6_57 bitb_6_57 word6_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_57 q_7_57 qb_7_57 bit_7_57 bitb_7_57 word7_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_57 q_8_57 qb_8_57 bit_8_57 bitb_8_57 word8_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_57 q_9_57 qb_9_57 bit_9_57 bitb_9_57 word9_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_57 q_10_57 qb_10_57 bit_10_57 bitb_10_57 word10_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_57 q_11_57 qb_11_57 bit_11_57 bitb_11_57 word11_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_57 q_12_57 qb_12_57 bit_12_57 bitb_12_57 word12_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_57 q_13_57 qb_13_57 bit_13_57 bitb_13_57 word13_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_57 q_14_57 qb_14_57 bit_14_57 bitb_14_57 word14_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_57 q_15_57 qb_15_57 bit_15_57 bitb_15_57 word15_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_57 q_16_57 qb_16_57 bit_16_57 bitb_16_57 word16_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_57 q_17_57 qb_17_57 bit_17_57 bitb_17_57 word17_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_57 q_18_57 qb_18_57 bit_18_57 bitb_18_57 word18_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_57 q_19_57 qb_19_57 bit_19_57 bitb_19_57 word19_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_57 q_20_57 qb_20_57 bit_20_57 bitb_20_57 word20_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_57 q_21_57 qb_21_57 bit_21_57 bitb_21_57 word21_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_57 q_22_57 qb_22_57 bit_22_57 bitb_22_57 word22_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_57 q_23_57 qb_23_57 bit_23_57 bitb_23_57 word23_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_57 q_24_57 qb_24_57 bit_24_57 bitb_24_57 word24_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_57 q_25_57 qb_25_57 bit_25_57 bitb_25_57 word25_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_57 q_26_57 qb_26_57 bit_26_57 bitb_26_57 word26_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_57 q_27_57 qb_27_57 bit_27_57 bitb_27_57 word27_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_57 q_28_57 qb_28_57 bit_28_57 bitb_28_57 word28_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_57 q_29_57 qb_29_57 bit_29_57 bitb_29_57 word29_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_57 q_30_57 qb_30_57 bit_30_57 bitb_30_57 word30_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_57 q_31_57 qb_31_57 bit_31_57 bitb_31_57 word31_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_57 q_32_57 qb_32_57 bit_32_57 bitb_32_57 word32_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_57 q_33_57 qb_33_57 bit_33_57 bitb_33_57 word33_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_57 q_34_57 qb_34_57 bit_34_57 bitb_34_57 word34_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_57 q_35_57 qb_35_57 bit_35_57 bitb_35_57 word35_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_57 q_36_57 qb_36_57 bit_36_57 bitb_36_57 word36_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_57 q_37_57 qb_37_57 bit_37_57 bitb_37_57 word37_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_57 q_38_57 qb_38_57 bit_38_57 bitb_38_57 word38_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_57 q_39_57 qb_39_57 bit_39_57 bitb_39_57 word39_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_57 q_40_57 qb_40_57 bit_40_57 bitb_40_57 word40_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_57 q_41_57 qb_41_57 bit_41_57 bitb_41_57 word41_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_57 q_42_57 qb_42_57 bit_42_57 bitb_42_57 word42_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_57 q_43_57 qb_43_57 bit_43_57 bitb_43_57 word43_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_57 q_44_57 qb_44_57 bit_44_57 bitb_44_57 word44_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_57 q_45_57 qb_45_57 bit_45_57 bitb_45_57 word45_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_57 q_46_57 qb_46_57 bit_46_57 bitb_46_57 word46_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_57 q_47_57 qb_47_57 bit_47_57 bitb_47_57 word47_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_57 q_48_57 qb_48_57 bit_48_57 bitb_48_57 word48_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_57 q_49_57 qb_49_57 bit_49_57 bitb_49_57 word49_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_57 q_50_57 qb_50_57 bit_50_57 bitb_50_57 word50_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_57 q_51_57 qb_51_57 bit_51_57 bitb_51_57 word51_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_57 q_52_57 qb_52_57 bit_52_57 bitb_52_57 word52_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_57 q_53_57 qb_53_57 bit_53_57 bitb_53_57 word53_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_57 q_54_57 qb_54_57 bit_54_57 bitb_54_57 word54_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_57 q_55_57 qb_55_57 bit_55_57 bitb_55_57 word55_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_57 q_56_57 qb_56_57 bit_56_57 bitb_56_57 word56_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_57 q_57_57 qb_57_57 bit_57_57 bitb_57_57 word57_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_57 q_58_57 qb_58_57 bit_58_57 bitb_58_57 word58_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_57 q_59_57 qb_59_57 bit_59_57 bitb_59_57 word59_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_57 q_60_57 qb_60_57 bit_60_57 bitb_60_57 word60_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_57 q_61_57 qb_61_57 bit_61_57 bitb_61_57 word61_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_57 q_62_57 qb_62_57 bit_62_57 bitb_62_57 word62_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_57 q_63_57 qb_63_57 bit_63_57 bitb_63_57 word63_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_57 q_64_57 qb_64_57 bit_64_57 bitb_64_57 word64_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_57 q_65_57 qb_65_57 bit_65_57 bitb_65_57 word65_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_57 q_66_57 qb_66_57 bit_66_57 bitb_66_57 word66_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_57 q_67_57 qb_67_57 bit_67_57 bitb_67_57 word67_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_57 q_68_57 qb_68_57 bit_68_57 bitb_68_57 word68_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_57 q_69_57 qb_69_57 bit_69_57 bitb_69_57 word69_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_57 q_70_57 qb_70_57 bit_70_57 bitb_70_57 word70_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_57 q_71_57 qb_71_57 bit_71_57 bitb_71_57 word71_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_57 q_72_57 qb_72_57 bit_72_57 bitb_72_57 word72_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_57 q_73_57 qb_73_57 bit_73_57 bitb_73_57 word73_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_57 q_74_57 qb_74_57 bit_74_57 bitb_74_57 word74_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_57 q_75_57 qb_75_57 bit_75_57 bitb_75_57 word75_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_57 q_76_57 qb_76_57 bit_76_57 bitb_76_57 word76_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_57 q_77_57 qb_77_57 bit_77_57 bitb_77_57 word77_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_57 q_78_57 qb_78_57 bit_78_57 bitb_78_57 word78_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_57 q_79_57 qb_79_57 bit_79_57 bitb_79_57 word79_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_57 q_80_57 qb_80_57 bit_80_57 bitb_80_57 word80_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_57 q_81_57 qb_81_57 bit_81_57 bitb_81_57 word81_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_57 q_82_57 qb_82_57 bit_82_57 bitb_82_57 word82_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_57 q_83_57 qb_83_57 bit_83_57 bitb_83_57 word83_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_57 q_84_57 qb_84_57 bit_84_57 bitb_84_57 word84_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_57 q_85_57 qb_85_57 bit_85_57 bitb_85_57 word85_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_57 q_86_57 qb_86_57 bit_86_57 bitb_86_57 word86_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_57 q_87_57 qb_87_57 bit_87_57 bitb_87_57 word87_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_57 q_88_57 qb_88_57 bit_88_57 bitb_88_57 word88_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_57 q_89_57 qb_89_57 bit_89_57 bitb_89_57 word89_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_57 q_90_57 qb_90_57 bit_90_57 bitb_90_57 word90_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_57 q_91_57 qb_91_57 bit_91_57 bitb_91_57 word91_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_57 q_92_57 qb_92_57 bit_92_57 bitb_92_57 word92_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_57 q_93_57 qb_93_57 bit_93_57 bitb_93_57 word93_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_57 q_94_57 qb_94_57 bit_94_57 bitb_94_57 word94_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_57 q_95_57 qb_95_57 bit_95_57 bitb_95_57 word95_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_57 q_96_57 qb_96_57 bit_96_57 bitb_96_57 word96_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_57 q_97_57 qb_97_57 bit_97_57 bitb_97_57 word97_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_57 q_98_57 qb_98_57 bit_98_57 bitb_98_57 word98_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_57 q_99_57 qb_99_57 bit_99_57 bitb_99_57 word99_57 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_58 q_0_58 qb_0_58 bit_0_58 bitb_0_58 word0_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_58 q_1_58 qb_1_58 bit_1_58 bitb_1_58 word1_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_58 q_2_58 qb_2_58 bit_2_58 bitb_2_58 word2_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_58 q_3_58 qb_3_58 bit_3_58 bitb_3_58 word3_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_58 q_4_58 qb_4_58 bit_4_58 bitb_4_58 word4_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_58 q_5_58 qb_5_58 bit_5_58 bitb_5_58 word5_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_58 q_6_58 qb_6_58 bit_6_58 bitb_6_58 word6_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_58 q_7_58 qb_7_58 bit_7_58 bitb_7_58 word7_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_58 q_8_58 qb_8_58 bit_8_58 bitb_8_58 word8_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_58 q_9_58 qb_9_58 bit_9_58 bitb_9_58 word9_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_58 q_10_58 qb_10_58 bit_10_58 bitb_10_58 word10_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_58 q_11_58 qb_11_58 bit_11_58 bitb_11_58 word11_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_58 q_12_58 qb_12_58 bit_12_58 bitb_12_58 word12_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_58 q_13_58 qb_13_58 bit_13_58 bitb_13_58 word13_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_58 q_14_58 qb_14_58 bit_14_58 bitb_14_58 word14_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_58 q_15_58 qb_15_58 bit_15_58 bitb_15_58 word15_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_58 q_16_58 qb_16_58 bit_16_58 bitb_16_58 word16_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_58 q_17_58 qb_17_58 bit_17_58 bitb_17_58 word17_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_58 q_18_58 qb_18_58 bit_18_58 bitb_18_58 word18_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_58 q_19_58 qb_19_58 bit_19_58 bitb_19_58 word19_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_58 q_20_58 qb_20_58 bit_20_58 bitb_20_58 word20_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_58 q_21_58 qb_21_58 bit_21_58 bitb_21_58 word21_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_58 q_22_58 qb_22_58 bit_22_58 bitb_22_58 word22_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_58 q_23_58 qb_23_58 bit_23_58 bitb_23_58 word23_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_58 q_24_58 qb_24_58 bit_24_58 bitb_24_58 word24_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_58 q_25_58 qb_25_58 bit_25_58 bitb_25_58 word25_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_58 q_26_58 qb_26_58 bit_26_58 bitb_26_58 word26_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_58 q_27_58 qb_27_58 bit_27_58 bitb_27_58 word27_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_58 q_28_58 qb_28_58 bit_28_58 bitb_28_58 word28_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_58 q_29_58 qb_29_58 bit_29_58 bitb_29_58 word29_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_58 q_30_58 qb_30_58 bit_30_58 bitb_30_58 word30_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_58 q_31_58 qb_31_58 bit_31_58 bitb_31_58 word31_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_58 q_32_58 qb_32_58 bit_32_58 bitb_32_58 word32_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_58 q_33_58 qb_33_58 bit_33_58 bitb_33_58 word33_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_58 q_34_58 qb_34_58 bit_34_58 bitb_34_58 word34_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_58 q_35_58 qb_35_58 bit_35_58 bitb_35_58 word35_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_58 q_36_58 qb_36_58 bit_36_58 bitb_36_58 word36_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_58 q_37_58 qb_37_58 bit_37_58 bitb_37_58 word37_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_58 q_38_58 qb_38_58 bit_38_58 bitb_38_58 word38_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_58 q_39_58 qb_39_58 bit_39_58 bitb_39_58 word39_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_58 q_40_58 qb_40_58 bit_40_58 bitb_40_58 word40_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_58 q_41_58 qb_41_58 bit_41_58 bitb_41_58 word41_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_58 q_42_58 qb_42_58 bit_42_58 bitb_42_58 word42_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_58 q_43_58 qb_43_58 bit_43_58 bitb_43_58 word43_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_58 q_44_58 qb_44_58 bit_44_58 bitb_44_58 word44_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_58 q_45_58 qb_45_58 bit_45_58 bitb_45_58 word45_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_58 q_46_58 qb_46_58 bit_46_58 bitb_46_58 word46_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_58 q_47_58 qb_47_58 bit_47_58 bitb_47_58 word47_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_58 q_48_58 qb_48_58 bit_48_58 bitb_48_58 word48_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_58 q_49_58 qb_49_58 bit_49_58 bitb_49_58 word49_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_58 q_50_58 qb_50_58 bit_50_58 bitb_50_58 word50_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_58 q_51_58 qb_51_58 bit_51_58 bitb_51_58 word51_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_58 q_52_58 qb_52_58 bit_52_58 bitb_52_58 word52_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_58 q_53_58 qb_53_58 bit_53_58 bitb_53_58 word53_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_58 q_54_58 qb_54_58 bit_54_58 bitb_54_58 word54_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_58 q_55_58 qb_55_58 bit_55_58 bitb_55_58 word55_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_58 q_56_58 qb_56_58 bit_56_58 bitb_56_58 word56_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_58 q_57_58 qb_57_58 bit_57_58 bitb_57_58 word57_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_58 q_58_58 qb_58_58 bit_58_58 bitb_58_58 word58_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_58 q_59_58 qb_59_58 bit_59_58 bitb_59_58 word59_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_58 q_60_58 qb_60_58 bit_60_58 bitb_60_58 word60_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_58 q_61_58 qb_61_58 bit_61_58 bitb_61_58 word61_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_58 q_62_58 qb_62_58 bit_62_58 bitb_62_58 word62_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_58 q_63_58 qb_63_58 bit_63_58 bitb_63_58 word63_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_58 q_64_58 qb_64_58 bit_64_58 bitb_64_58 word64_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_58 q_65_58 qb_65_58 bit_65_58 bitb_65_58 word65_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_58 q_66_58 qb_66_58 bit_66_58 bitb_66_58 word66_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_58 q_67_58 qb_67_58 bit_67_58 bitb_67_58 word67_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_58 q_68_58 qb_68_58 bit_68_58 bitb_68_58 word68_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_58 q_69_58 qb_69_58 bit_69_58 bitb_69_58 word69_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_58 q_70_58 qb_70_58 bit_70_58 bitb_70_58 word70_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_58 q_71_58 qb_71_58 bit_71_58 bitb_71_58 word71_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_58 q_72_58 qb_72_58 bit_72_58 bitb_72_58 word72_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_58 q_73_58 qb_73_58 bit_73_58 bitb_73_58 word73_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_58 q_74_58 qb_74_58 bit_74_58 bitb_74_58 word74_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_58 q_75_58 qb_75_58 bit_75_58 bitb_75_58 word75_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_58 q_76_58 qb_76_58 bit_76_58 bitb_76_58 word76_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_58 q_77_58 qb_77_58 bit_77_58 bitb_77_58 word77_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_58 q_78_58 qb_78_58 bit_78_58 bitb_78_58 word78_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_58 q_79_58 qb_79_58 bit_79_58 bitb_79_58 word79_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_58 q_80_58 qb_80_58 bit_80_58 bitb_80_58 word80_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_58 q_81_58 qb_81_58 bit_81_58 bitb_81_58 word81_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_58 q_82_58 qb_82_58 bit_82_58 bitb_82_58 word82_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_58 q_83_58 qb_83_58 bit_83_58 bitb_83_58 word83_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_58 q_84_58 qb_84_58 bit_84_58 bitb_84_58 word84_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_58 q_85_58 qb_85_58 bit_85_58 bitb_85_58 word85_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_58 q_86_58 qb_86_58 bit_86_58 bitb_86_58 word86_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_58 q_87_58 qb_87_58 bit_87_58 bitb_87_58 word87_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_58 q_88_58 qb_88_58 bit_88_58 bitb_88_58 word88_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_58 q_89_58 qb_89_58 bit_89_58 bitb_89_58 word89_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_58 q_90_58 qb_90_58 bit_90_58 bitb_90_58 word90_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_58 q_91_58 qb_91_58 bit_91_58 bitb_91_58 word91_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_58 q_92_58 qb_92_58 bit_92_58 bitb_92_58 word92_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_58 q_93_58 qb_93_58 bit_93_58 bitb_93_58 word93_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_58 q_94_58 qb_94_58 bit_94_58 bitb_94_58 word94_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_58 q_95_58 qb_95_58 bit_95_58 bitb_95_58 word95_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_58 q_96_58 qb_96_58 bit_96_58 bitb_96_58 word96_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_58 q_97_58 qb_97_58 bit_97_58 bitb_97_58 word97_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_58 q_98_58 qb_98_58 bit_98_58 bitb_98_58 word98_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_58 q_99_58 qb_99_58 bit_99_58 bitb_99_58 word99_58 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_59 q_0_59 qb_0_59 bit_0_59 bitb_0_59 word0_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_59 q_1_59 qb_1_59 bit_1_59 bitb_1_59 word1_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_59 q_2_59 qb_2_59 bit_2_59 bitb_2_59 word2_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_59 q_3_59 qb_3_59 bit_3_59 bitb_3_59 word3_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_59 q_4_59 qb_4_59 bit_4_59 bitb_4_59 word4_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_59 q_5_59 qb_5_59 bit_5_59 bitb_5_59 word5_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_59 q_6_59 qb_6_59 bit_6_59 bitb_6_59 word6_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_59 q_7_59 qb_7_59 bit_7_59 bitb_7_59 word7_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_59 q_8_59 qb_8_59 bit_8_59 bitb_8_59 word8_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_59 q_9_59 qb_9_59 bit_9_59 bitb_9_59 word9_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_59 q_10_59 qb_10_59 bit_10_59 bitb_10_59 word10_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_59 q_11_59 qb_11_59 bit_11_59 bitb_11_59 word11_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_59 q_12_59 qb_12_59 bit_12_59 bitb_12_59 word12_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_59 q_13_59 qb_13_59 bit_13_59 bitb_13_59 word13_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_59 q_14_59 qb_14_59 bit_14_59 bitb_14_59 word14_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_59 q_15_59 qb_15_59 bit_15_59 bitb_15_59 word15_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_59 q_16_59 qb_16_59 bit_16_59 bitb_16_59 word16_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_59 q_17_59 qb_17_59 bit_17_59 bitb_17_59 word17_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_59 q_18_59 qb_18_59 bit_18_59 bitb_18_59 word18_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_59 q_19_59 qb_19_59 bit_19_59 bitb_19_59 word19_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_59 q_20_59 qb_20_59 bit_20_59 bitb_20_59 word20_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_59 q_21_59 qb_21_59 bit_21_59 bitb_21_59 word21_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_59 q_22_59 qb_22_59 bit_22_59 bitb_22_59 word22_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_59 q_23_59 qb_23_59 bit_23_59 bitb_23_59 word23_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_59 q_24_59 qb_24_59 bit_24_59 bitb_24_59 word24_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_59 q_25_59 qb_25_59 bit_25_59 bitb_25_59 word25_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_59 q_26_59 qb_26_59 bit_26_59 bitb_26_59 word26_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_59 q_27_59 qb_27_59 bit_27_59 bitb_27_59 word27_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_59 q_28_59 qb_28_59 bit_28_59 bitb_28_59 word28_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_59 q_29_59 qb_29_59 bit_29_59 bitb_29_59 word29_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_59 q_30_59 qb_30_59 bit_30_59 bitb_30_59 word30_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_59 q_31_59 qb_31_59 bit_31_59 bitb_31_59 word31_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_59 q_32_59 qb_32_59 bit_32_59 bitb_32_59 word32_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_59 q_33_59 qb_33_59 bit_33_59 bitb_33_59 word33_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_59 q_34_59 qb_34_59 bit_34_59 bitb_34_59 word34_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_59 q_35_59 qb_35_59 bit_35_59 bitb_35_59 word35_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_59 q_36_59 qb_36_59 bit_36_59 bitb_36_59 word36_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_59 q_37_59 qb_37_59 bit_37_59 bitb_37_59 word37_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_59 q_38_59 qb_38_59 bit_38_59 bitb_38_59 word38_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_59 q_39_59 qb_39_59 bit_39_59 bitb_39_59 word39_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_59 q_40_59 qb_40_59 bit_40_59 bitb_40_59 word40_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_59 q_41_59 qb_41_59 bit_41_59 bitb_41_59 word41_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_59 q_42_59 qb_42_59 bit_42_59 bitb_42_59 word42_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_59 q_43_59 qb_43_59 bit_43_59 bitb_43_59 word43_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_59 q_44_59 qb_44_59 bit_44_59 bitb_44_59 word44_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_59 q_45_59 qb_45_59 bit_45_59 bitb_45_59 word45_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_59 q_46_59 qb_46_59 bit_46_59 bitb_46_59 word46_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_59 q_47_59 qb_47_59 bit_47_59 bitb_47_59 word47_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_59 q_48_59 qb_48_59 bit_48_59 bitb_48_59 word48_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_59 q_49_59 qb_49_59 bit_49_59 bitb_49_59 word49_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_59 q_50_59 qb_50_59 bit_50_59 bitb_50_59 word50_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_59 q_51_59 qb_51_59 bit_51_59 bitb_51_59 word51_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_59 q_52_59 qb_52_59 bit_52_59 bitb_52_59 word52_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_59 q_53_59 qb_53_59 bit_53_59 bitb_53_59 word53_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_59 q_54_59 qb_54_59 bit_54_59 bitb_54_59 word54_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_59 q_55_59 qb_55_59 bit_55_59 bitb_55_59 word55_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_59 q_56_59 qb_56_59 bit_56_59 bitb_56_59 word56_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_59 q_57_59 qb_57_59 bit_57_59 bitb_57_59 word57_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_59 q_58_59 qb_58_59 bit_58_59 bitb_58_59 word58_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_59 q_59_59 qb_59_59 bit_59_59 bitb_59_59 word59_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_59 q_60_59 qb_60_59 bit_60_59 bitb_60_59 word60_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_59 q_61_59 qb_61_59 bit_61_59 bitb_61_59 word61_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_59 q_62_59 qb_62_59 bit_62_59 bitb_62_59 word62_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_59 q_63_59 qb_63_59 bit_63_59 bitb_63_59 word63_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_59 q_64_59 qb_64_59 bit_64_59 bitb_64_59 word64_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_59 q_65_59 qb_65_59 bit_65_59 bitb_65_59 word65_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_59 q_66_59 qb_66_59 bit_66_59 bitb_66_59 word66_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_59 q_67_59 qb_67_59 bit_67_59 bitb_67_59 word67_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_59 q_68_59 qb_68_59 bit_68_59 bitb_68_59 word68_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_59 q_69_59 qb_69_59 bit_69_59 bitb_69_59 word69_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_59 q_70_59 qb_70_59 bit_70_59 bitb_70_59 word70_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_59 q_71_59 qb_71_59 bit_71_59 bitb_71_59 word71_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_59 q_72_59 qb_72_59 bit_72_59 bitb_72_59 word72_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_59 q_73_59 qb_73_59 bit_73_59 bitb_73_59 word73_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_59 q_74_59 qb_74_59 bit_74_59 bitb_74_59 word74_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_59 q_75_59 qb_75_59 bit_75_59 bitb_75_59 word75_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_59 q_76_59 qb_76_59 bit_76_59 bitb_76_59 word76_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_59 q_77_59 qb_77_59 bit_77_59 bitb_77_59 word77_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_59 q_78_59 qb_78_59 bit_78_59 bitb_78_59 word78_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_59 q_79_59 qb_79_59 bit_79_59 bitb_79_59 word79_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_59 q_80_59 qb_80_59 bit_80_59 bitb_80_59 word80_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_59 q_81_59 qb_81_59 bit_81_59 bitb_81_59 word81_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_59 q_82_59 qb_82_59 bit_82_59 bitb_82_59 word82_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_59 q_83_59 qb_83_59 bit_83_59 bitb_83_59 word83_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_59 q_84_59 qb_84_59 bit_84_59 bitb_84_59 word84_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_59 q_85_59 qb_85_59 bit_85_59 bitb_85_59 word85_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_59 q_86_59 qb_86_59 bit_86_59 bitb_86_59 word86_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_59 q_87_59 qb_87_59 bit_87_59 bitb_87_59 word87_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_59 q_88_59 qb_88_59 bit_88_59 bitb_88_59 word88_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_59 q_89_59 qb_89_59 bit_89_59 bitb_89_59 word89_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_59 q_90_59 qb_90_59 bit_90_59 bitb_90_59 word90_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_59 q_91_59 qb_91_59 bit_91_59 bitb_91_59 word91_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_59 q_92_59 qb_92_59 bit_92_59 bitb_92_59 word92_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_59 q_93_59 qb_93_59 bit_93_59 bitb_93_59 word93_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_59 q_94_59 qb_94_59 bit_94_59 bitb_94_59 word94_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_59 q_95_59 qb_95_59 bit_95_59 bitb_95_59 word95_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_59 q_96_59 qb_96_59 bit_96_59 bitb_96_59 word96_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_59 q_97_59 qb_97_59 bit_97_59 bitb_97_59 word97_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_59 q_98_59 qb_98_59 bit_98_59 bitb_98_59 word98_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_59 q_99_59 qb_99_59 bit_99_59 bitb_99_59 word99_59 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_60 q_0_60 qb_0_60 bit_0_60 bitb_0_60 word0_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_60 q_1_60 qb_1_60 bit_1_60 bitb_1_60 word1_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_60 q_2_60 qb_2_60 bit_2_60 bitb_2_60 word2_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_60 q_3_60 qb_3_60 bit_3_60 bitb_3_60 word3_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_60 q_4_60 qb_4_60 bit_4_60 bitb_4_60 word4_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_60 q_5_60 qb_5_60 bit_5_60 bitb_5_60 word5_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_60 q_6_60 qb_6_60 bit_6_60 bitb_6_60 word6_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_60 q_7_60 qb_7_60 bit_7_60 bitb_7_60 word7_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_60 q_8_60 qb_8_60 bit_8_60 bitb_8_60 word8_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_60 q_9_60 qb_9_60 bit_9_60 bitb_9_60 word9_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_60 q_10_60 qb_10_60 bit_10_60 bitb_10_60 word10_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_60 q_11_60 qb_11_60 bit_11_60 bitb_11_60 word11_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_60 q_12_60 qb_12_60 bit_12_60 bitb_12_60 word12_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_60 q_13_60 qb_13_60 bit_13_60 bitb_13_60 word13_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_60 q_14_60 qb_14_60 bit_14_60 bitb_14_60 word14_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_60 q_15_60 qb_15_60 bit_15_60 bitb_15_60 word15_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_60 q_16_60 qb_16_60 bit_16_60 bitb_16_60 word16_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_60 q_17_60 qb_17_60 bit_17_60 bitb_17_60 word17_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_60 q_18_60 qb_18_60 bit_18_60 bitb_18_60 word18_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_60 q_19_60 qb_19_60 bit_19_60 bitb_19_60 word19_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_60 q_20_60 qb_20_60 bit_20_60 bitb_20_60 word20_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_60 q_21_60 qb_21_60 bit_21_60 bitb_21_60 word21_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_60 q_22_60 qb_22_60 bit_22_60 bitb_22_60 word22_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_60 q_23_60 qb_23_60 bit_23_60 bitb_23_60 word23_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_60 q_24_60 qb_24_60 bit_24_60 bitb_24_60 word24_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_60 q_25_60 qb_25_60 bit_25_60 bitb_25_60 word25_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_60 q_26_60 qb_26_60 bit_26_60 bitb_26_60 word26_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_60 q_27_60 qb_27_60 bit_27_60 bitb_27_60 word27_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_60 q_28_60 qb_28_60 bit_28_60 bitb_28_60 word28_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_60 q_29_60 qb_29_60 bit_29_60 bitb_29_60 word29_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_60 q_30_60 qb_30_60 bit_30_60 bitb_30_60 word30_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_60 q_31_60 qb_31_60 bit_31_60 bitb_31_60 word31_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_60 q_32_60 qb_32_60 bit_32_60 bitb_32_60 word32_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_60 q_33_60 qb_33_60 bit_33_60 bitb_33_60 word33_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_60 q_34_60 qb_34_60 bit_34_60 bitb_34_60 word34_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_60 q_35_60 qb_35_60 bit_35_60 bitb_35_60 word35_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_60 q_36_60 qb_36_60 bit_36_60 bitb_36_60 word36_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_60 q_37_60 qb_37_60 bit_37_60 bitb_37_60 word37_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_60 q_38_60 qb_38_60 bit_38_60 bitb_38_60 word38_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_60 q_39_60 qb_39_60 bit_39_60 bitb_39_60 word39_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_60 q_40_60 qb_40_60 bit_40_60 bitb_40_60 word40_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_60 q_41_60 qb_41_60 bit_41_60 bitb_41_60 word41_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_60 q_42_60 qb_42_60 bit_42_60 bitb_42_60 word42_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_60 q_43_60 qb_43_60 bit_43_60 bitb_43_60 word43_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_60 q_44_60 qb_44_60 bit_44_60 bitb_44_60 word44_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_60 q_45_60 qb_45_60 bit_45_60 bitb_45_60 word45_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_60 q_46_60 qb_46_60 bit_46_60 bitb_46_60 word46_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_60 q_47_60 qb_47_60 bit_47_60 bitb_47_60 word47_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_60 q_48_60 qb_48_60 bit_48_60 bitb_48_60 word48_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_60 q_49_60 qb_49_60 bit_49_60 bitb_49_60 word49_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_60 q_50_60 qb_50_60 bit_50_60 bitb_50_60 word50_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_60 q_51_60 qb_51_60 bit_51_60 bitb_51_60 word51_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_60 q_52_60 qb_52_60 bit_52_60 bitb_52_60 word52_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_60 q_53_60 qb_53_60 bit_53_60 bitb_53_60 word53_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_60 q_54_60 qb_54_60 bit_54_60 bitb_54_60 word54_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_60 q_55_60 qb_55_60 bit_55_60 bitb_55_60 word55_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_60 q_56_60 qb_56_60 bit_56_60 bitb_56_60 word56_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_60 q_57_60 qb_57_60 bit_57_60 bitb_57_60 word57_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_60 q_58_60 qb_58_60 bit_58_60 bitb_58_60 word58_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_60 q_59_60 qb_59_60 bit_59_60 bitb_59_60 word59_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_60 q_60_60 qb_60_60 bit_60_60 bitb_60_60 word60_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_60 q_61_60 qb_61_60 bit_61_60 bitb_61_60 word61_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_60 q_62_60 qb_62_60 bit_62_60 bitb_62_60 word62_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_60 q_63_60 qb_63_60 bit_63_60 bitb_63_60 word63_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_60 q_64_60 qb_64_60 bit_64_60 bitb_64_60 word64_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_60 q_65_60 qb_65_60 bit_65_60 bitb_65_60 word65_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_60 q_66_60 qb_66_60 bit_66_60 bitb_66_60 word66_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_60 q_67_60 qb_67_60 bit_67_60 bitb_67_60 word67_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_60 q_68_60 qb_68_60 bit_68_60 bitb_68_60 word68_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_60 q_69_60 qb_69_60 bit_69_60 bitb_69_60 word69_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_60 q_70_60 qb_70_60 bit_70_60 bitb_70_60 word70_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_60 q_71_60 qb_71_60 bit_71_60 bitb_71_60 word71_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_60 q_72_60 qb_72_60 bit_72_60 bitb_72_60 word72_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_60 q_73_60 qb_73_60 bit_73_60 bitb_73_60 word73_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_60 q_74_60 qb_74_60 bit_74_60 bitb_74_60 word74_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_60 q_75_60 qb_75_60 bit_75_60 bitb_75_60 word75_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_60 q_76_60 qb_76_60 bit_76_60 bitb_76_60 word76_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_60 q_77_60 qb_77_60 bit_77_60 bitb_77_60 word77_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_60 q_78_60 qb_78_60 bit_78_60 bitb_78_60 word78_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_60 q_79_60 qb_79_60 bit_79_60 bitb_79_60 word79_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_60 q_80_60 qb_80_60 bit_80_60 bitb_80_60 word80_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_60 q_81_60 qb_81_60 bit_81_60 bitb_81_60 word81_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_60 q_82_60 qb_82_60 bit_82_60 bitb_82_60 word82_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_60 q_83_60 qb_83_60 bit_83_60 bitb_83_60 word83_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_60 q_84_60 qb_84_60 bit_84_60 bitb_84_60 word84_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_60 q_85_60 qb_85_60 bit_85_60 bitb_85_60 word85_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_60 q_86_60 qb_86_60 bit_86_60 bitb_86_60 word86_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_60 q_87_60 qb_87_60 bit_87_60 bitb_87_60 word87_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_60 q_88_60 qb_88_60 bit_88_60 bitb_88_60 word88_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_60 q_89_60 qb_89_60 bit_89_60 bitb_89_60 word89_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_60 q_90_60 qb_90_60 bit_90_60 bitb_90_60 word90_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_60 q_91_60 qb_91_60 bit_91_60 bitb_91_60 word91_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_60 q_92_60 qb_92_60 bit_92_60 bitb_92_60 word92_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_60 q_93_60 qb_93_60 bit_93_60 bitb_93_60 word93_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_60 q_94_60 qb_94_60 bit_94_60 bitb_94_60 word94_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_60 q_95_60 qb_95_60 bit_95_60 bitb_95_60 word95_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_60 q_96_60 qb_96_60 bit_96_60 bitb_96_60 word96_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_60 q_97_60 qb_97_60 bit_97_60 bitb_97_60 word97_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_60 q_98_60 qb_98_60 bit_98_60 bitb_98_60 word98_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_60 q_99_60 qb_99_60 bit_99_60 bitb_99_60 word99_60 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_61 q_0_61 qb_0_61 bit_0_61 bitb_0_61 word0_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_61 q_1_61 qb_1_61 bit_1_61 bitb_1_61 word1_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_61 q_2_61 qb_2_61 bit_2_61 bitb_2_61 word2_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_61 q_3_61 qb_3_61 bit_3_61 bitb_3_61 word3_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_61 q_4_61 qb_4_61 bit_4_61 bitb_4_61 word4_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_61 q_5_61 qb_5_61 bit_5_61 bitb_5_61 word5_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_61 q_6_61 qb_6_61 bit_6_61 bitb_6_61 word6_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_61 q_7_61 qb_7_61 bit_7_61 bitb_7_61 word7_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_61 q_8_61 qb_8_61 bit_8_61 bitb_8_61 word8_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_61 q_9_61 qb_9_61 bit_9_61 bitb_9_61 word9_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_61 q_10_61 qb_10_61 bit_10_61 bitb_10_61 word10_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_61 q_11_61 qb_11_61 bit_11_61 bitb_11_61 word11_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_61 q_12_61 qb_12_61 bit_12_61 bitb_12_61 word12_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_61 q_13_61 qb_13_61 bit_13_61 bitb_13_61 word13_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_61 q_14_61 qb_14_61 bit_14_61 bitb_14_61 word14_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_61 q_15_61 qb_15_61 bit_15_61 bitb_15_61 word15_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_61 q_16_61 qb_16_61 bit_16_61 bitb_16_61 word16_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_61 q_17_61 qb_17_61 bit_17_61 bitb_17_61 word17_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_61 q_18_61 qb_18_61 bit_18_61 bitb_18_61 word18_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_61 q_19_61 qb_19_61 bit_19_61 bitb_19_61 word19_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_61 q_20_61 qb_20_61 bit_20_61 bitb_20_61 word20_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_61 q_21_61 qb_21_61 bit_21_61 bitb_21_61 word21_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_61 q_22_61 qb_22_61 bit_22_61 bitb_22_61 word22_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_61 q_23_61 qb_23_61 bit_23_61 bitb_23_61 word23_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_61 q_24_61 qb_24_61 bit_24_61 bitb_24_61 word24_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_61 q_25_61 qb_25_61 bit_25_61 bitb_25_61 word25_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_61 q_26_61 qb_26_61 bit_26_61 bitb_26_61 word26_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_61 q_27_61 qb_27_61 bit_27_61 bitb_27_61 word27_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_61 q_28_61 qb_28_61 bit_28_61 bitb_28_61 word28_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_61 q_29_61 qb_29_61 bit_29_61 bitb_29_61 word29_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_61 q_30_61 qb_30_61 bit_30_61 bitb_30_61 word30_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_61 q_31_61 qb_31_61 bit_31_61 bitb_31_61 word31_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_61 q_32_61 qb_32_61 bit_32_61 bitb_32_61 word32_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_61 q_33_61 qb_33_61 bit_33_61 bitb_33_61 word33_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_61 q_34_61 qb_34_61 bit_34_61 bitb_34_61 word34_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_61 q_35_61 qb_35_61 bit_35_61 bitb_35_61 word35_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_61 q_36_61 qb_36_61 bit_36_61 bitb_36_61 word36_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_61 q_37_61 qb_37_61 bit_37_61 bitb_37_61 word37_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_61 q_38_61 qb_38_61 bit_38_61 bitb_38_61 word38_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_61 q_39_61 qb_39_61 bit_39_61 bitb_39_61 word39_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_61 q_40_61 qb_40_61 bit_40_61 bitb_40_61 word40_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_61 q_41_61 qb_41_61 bit_41_61 bitb_41_61 word41_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_61 q_42_61 qb_42_61 bit_42_61 bitb_42_61 word42_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_61 q_43_61 qb_43_61 bit_43_61 bitb_43_61 word43_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_61 q_44_61 qb_44_61 bit_44_61 bitb_44_61 word44_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_61 q_45_61 qb_45_61 bit_45_61 bitb_45_61 word45_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_61 q_46_61 qb_46_61 bit_46_61 bitb_46_61 word46_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_61 q_47_61 qb_47_61 bit_47_61 bitb_47_61 word47_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_61 q_48_61 qb_48_61 bit_48_61 bitb_48_61 word48_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_61 q_49_61 qb_49_61 bit_49_61 bitb_49_61 word49_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_61 q_50_61 qb_50_61 bit_50_61 bitb_50_61 word50_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_61 q_51_61 qb_51_61 bit_51_61 bitb_51_61 word51_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_61 q_52_61 qb_52_61 bit_52_61 bitb_52_61 word52_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_61 q_53_61 qb_53_61 bit_53_61 bitb_53_61 word53_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_61 q_54_61 qb_54_61 bit_54_61 bitb_54_61 word54_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_61 q_55_61 qb_55_61 bit_55_61 bitb_55_61 word55_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_61 q_56_61 qb_56_61 bit_56_61 bitb_56_61 word56_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_61 q_57_61 qb_57_61 bit_57_61 bitb_57_61 word57_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_61 q_58_61 qb_58_61 bit_58_61 bitb_58_61 word58_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_61 q_59_61 qb_59_61 bit_59_61 bitb_59_61 word59_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_61 q_60_61 qb_60_61 bit_60_61 bitb_60_61 word60_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_61 q_61_61 qb_61_61 bit_61_61 bitb_61_61 word61_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_61 q_62_61 qb_62_61 bit_62_61 bitb_62_61 word62_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_61 q_63_61 qb_63_61 bit_63_61 bitb_63_61 word63_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_61 q_64_61 qb_64_61 bit_64_61 bitb_64_61 word64_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_61 q_65_61 qb_65_61 bit_65_61 bitb_65_61 word65_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_61 q_66_61 qb_66_61 bit_66_61 bitb_66_61 word66_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_61 q_67_61 qb_67_61 bit_67_61 bitb_67_61 word67_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_61 q_68_61 qb_68_61 bit_68_61 bitb_68_61 word68_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_61 q_69_61 qb_69_61 bit_69_61 bitb_69_61 word69_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_61 q_70_61 qb_70_61 bit_70_61 bitb_70_61 word70_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_61 q_71_61 qb_71_61 bit_71_61 bitb_71_61 word71_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_61 q_72_61 qb_72_61 bit_72_61 bitb_72_61 word72_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_61 q_73_61 qb_73_61 bit_73_61 bitb_73_61 word73_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_61 q_74_61 qb_74_61 bit_74_61 bitb_74_61 word74_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_61 q_75_61 qb_75_61 bit_75_61 bitb_75_61 word75_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_61 q_76_61 qb_76_61 bit_76_61 bitb_76_61 word76_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_61 q_77_61 qb_77_61 bit_77_61 bitb_77_61 word77_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_61 q_78_61 qb_78_61 bit_78_61 bitb_78_61 word78_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_61 q_79_61 qb_79_61 bit_79_61 bitb_79_61 word79_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_61 q_80_61 qb_80_61 bit_80_61 bitb_80_61 word80_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_61 q_81_61 qb_81_61 bit_81_61 bitb_81_61 word81_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_61 q_82_61 qb_82_61 bit_82_61 bitb_82_61 word82_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_61 q_83_61 qb_83_61 bit_83_61 bitb_83_61 word83_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_61 q_84_61 qb_84_61 bit_84_61 bitb_84_61 word84_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_61 q_85_61 qb_85_61 bit_85_61 bitb_85_61 word85_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_61 q_86_61 qb_86_61 bit_86_61 bitb_86_61 word86_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_61 q_87_61 qb_87_61 bit_87_61 bitb_87_61 word87_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_61 q_88_61 qb_88_61 bit_88_61 bitb_88_61 word88_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_61 q_89_61 qb_89_61 bit_89_61 bitb_89_61 word89_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_61 q_90_61 qb_90_61 bit_90_61 bitb_90_61 word90_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_61 q_91_61 qb_91_61 bit_91_61 bitb_91_61 word91_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_61 q_92_61 qb_92_61 bit_92_61 bitb_92_61 word92_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_61 q_93_61 qb_93_61 bit_93_61 bitb_93_61 word93_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_61 q_94_61 qb_94_61 bit_94_61 bitb_94_61 word94_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_61 q_95_61 qb_95_61 bit_95_61 bitb_95_61 word95_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_61 q_96_61 qb_96_61 bit_96_61 bitb_96_61 word96_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_61 q_97_61 qb_97_61 bit_97_61 bitb_97_61 word97_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_61 q_98_61 qb_98_61 bit_98_61 bitb_98_61 word98_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_61 q_99_61 qb_99_61 bit_99_61 bitb_99_61 word99_61 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_62 q_0_62 qb_0_62 bit_0_62 bitb_0_62 word0_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_62 q_1_62 qb_1_62 bit_1_62 bitb_1_62 word1_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_62 q_2_62 qb_2_62 bit_2_62 bitb_2_62 word2_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_62 q_3_62 qb_3_62 bit_3_62 bitb_3_62 word3_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_62 q_4_62 qb_4_62 bit_4_62 bitb_4_62 word4_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_62 q_5_62 qb_5_62 bit_5_62 bitb_5_62 word5_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_62 q_6_62 qb_6_62 bit_6_62 bitb_6_62 word6_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_62 q_7_62 qb_7_62 bit_7_62 bitb_7_62 word7_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_62 q_8_62 qb_8_62 bit_8_62 bitb_8_62 word8_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_62 q_9_62 qb_9_62 bit_9_62 bitb_9_62 word9_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_62 q_10_62 qb_10_62 bit_10_62 bitb_10_62 word10_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_62 q_11_62 qb_11_62 bit_11_62 bitb_11_62 word11_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_62 q_12_62 qb_12_62 bit_12_62 bitb_12_62 word12_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_62 q_13_62 qb_13_62 bit_13_62 bitb_13_62 word13_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_62 q_14_62 qb_14_62 bit_14_62 bitb_14_62 word14_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_62 q_15_62 qb_15_62 bit_15_62 bitb_15_62 word15_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_62 q_16_62 qb_16_62 bit_16_62 bitb_16_62 word16_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_62 q_17_62 qb_17_62 bit_17_62 bitb_17_62 word17_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_62 q_18_62 qb_18_62 bit_18_62 bitb_18_62 word18_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_62 q_19_62 qb_19_62 bit_19_62 bitb_19_62 word19_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_62 q_20_62 qb_20_62 bit_20_62 bitb_20_62 word20_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_62 q_21_62 qb_21_62 bit_21_62 bitb_21_62 word21_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_62 q_22_62 qb_22_62 bit_22_62 bitb_22_62 word22_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_62 q_23_62 qb_23_62 bit_23_62 bitb_23_62 word23_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_62 q_24_62 qb_24_62 bit_24_62 bitb_24_62 word24_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_62 q_25_62 qb_25_62 bit_25_62 bitb_25_62 word25_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_62 q_26_62 qb_26_62 bit_26_62 bitb_26_62 word26_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_62 q_27_62 qb_27_62 bit_27_62 bitb_27_62 word27_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_62 q_28_62 qb_28_62 bit_28_62 bitb_28_62 word28_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_62 q_29_62 qb_29_62 bit_29_62 bitb_29_62 word29_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_62 q_30_62 qb_30_62 bit_30_62 bitb_30_62 word30_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_62 q_31_62 qb_31_62 bit_31_62 bitb_31_62 word31_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_62 q_32_62 qb_32_62 bit_32_62 bitb_32_62 word32_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_62 q_33_62 qb_33_62 bit_33_62 bitb_33_62 word33_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_62 q_34_62 qb_34_62 bit_34_62 bitb_34_62 word34_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_62 q_35_62 qb_35_62 bit_35_62 bitb_35_62 word35_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_62 q_36_62 qb_36_62 bit_36_62 bitb_36_62 word36_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_62 q_37_62 qb_37_62 bit_37_62 bitb_37_62 word37_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_62 q_38_62 qb_38_62 bit_38_62 bitb_38_62 word38_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_62 q_39_62 qb_39_62 bit_39_62 bitb_39_62 word39_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_62 q_40_62 qb_40_62 bit_40_62 bitb_40_62 word40_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_62 q_41_62 qb_41_62 bit_41_62 bitb_41_62 word41_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_62 q_42_62 qb_42_62 bit_42_62 bitb_42_62 word42_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_62 q_43_62 qb_43_62 bit_43_62 bitb_43_62 word43_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_62 q_44_62 qb_44_62 bit_44_62 bitb_44_62 word44_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_62 q_45_62 qb_45_62 bit_45_62 bitb_45_62 word45_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_62 q_46_62 qb_46_62 bit_46_62 bitb_46_62 word46_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_62 q_47_62 qb_47_62 bit_47_62 bitb_47_62 word47_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_62 q_48_62 qb_48_62 bit_48_62 bitb_48_62 word48_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_62 q_49_62 qb_49_62 bit_49_62 bitb_49_62 word49_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_62 q_50_62 qb_50_62 bit_50_62 bitb_50_62 word50_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_62 q_51_62 qb_51_62 bit_51_62 bitb_51_62 word51_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_62 q_52_62 qb_52_62 bit_52_62 bitb_52_62 word52_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_62 q_53_62 qb_53_62 bit_53_62 bitb_53_62 word53_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_62 q_54_62 qb_54_62 bit_54_62 bitb_54_62 word54_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_62 q_55_62 qb_55_62 bit_55_62 bitb_55_62 word55_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_62 q_56_62 qb_56_62 bit_56_62 bitb_56_62 word56_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_62 q_57_62 qb_57_62 bit_57_62 bitb_57_62 word57_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_62 q_58_62 qb_58_62 bit_58_62 bitb_58_62 word58_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_62 q_59_62 qb_59_62 bit_59_62 bitb_59_62 word59_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_62 q_60_62 qb_60_62 bit_60_62 bitb_60_62 word60_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_62 q_61_62 qb_61_62 bit_61_62 bitb_61_62 word61_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_62 q_62_62 qb_62_62 bit_62_62 bitb_62_62 word62_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_62 q_63_62 qb_63_62 bit_63_62 bitb_63_62 word63_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_62 q_64_62 qb_64_62 bit_64_62 bitb_64_62 word64_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_62 q_65_62 qb_65_62 bit_65_62 bitb_65_62 word65_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_62 q_66_62 qb_66_62 bit_66_62 bitb_66_62 word66_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_62 q_67_62 qb_67_62 bit_67_62 bitb_67_62 word67_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_62 q_68_62 qb_68_62 bit_68_62 bitb_68_62 word68_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_62 q_69_62 qb_69_62 bit_69_62 bitb_69_62 word69_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_62 q_70_62 qb_70_62 bit_70_62 bitb_70_62 word70_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_62 q_71_62 qb_71_62 bit_71_62 bitb_71_62 word71_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_62 q_72_62 qb_72_62 bit_72_62 bitb_72_62 word72_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_62 q_73_62 qb_73_62 bit_73_62 bitb_73_62 word73_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_62 q_74_62 qb_74_62 bit_74_62 bitb_74_62 word74_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_62 q_75_62 qb_75_62 bit_75_62 bitb_75_62 word75_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_62 q_76_62 qb_76_62 bit_76_62 bitb_76_62 word76_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_62 q_77_62 qb_77_62 bit_77_62 bitb_77_62 word77_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_62 q_78_62 qb_78_62 bit_78_62 bitb_78_62 word78_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_62 q_79_62 qb_79_62 bit_79_62 bitb_79_62 word79_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_62 q_80_62 qb_80_62 bit_80_62 bitb_80_62 word80_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_62 q_81_62 qb_81_62 bit_81_62 bitb_81_62 word81_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_62 q_82_62 qb_82_62 bit_82_62 bitb_82_62 word82_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_62 q_83_62 qb_83_62 bit_83_62 bitb_83_62 word83_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_62 q_84_62 qb_84_62 bit_84_62 bitb_84_62 word84_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_62 q_85_62 qb_85_62 bit_85_62 bitb_85_62 word85_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_62 q_86_62 qb_86_62 bit_86_62 bitb_86_62 word86_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_62 q_87_62 qb_87_62 bit_87_62 bitb_87_62 word87_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_62 q_88_62 qb_88_62 bit_88_62 bitb_88_62 word88_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_62 q_89_62 qb_89_62 bit_89_62 bitb_89_62 word89_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_62 q_90_62 qb_90_62 bit_90_62 bitb_90_62 word90_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_62 q_91_62 qb_91_62 bit_91_62 bitb_91_62 word91_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_62 q_92_62 qb_92_62 bit_92_62 bitb_92_62 word92_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_62 q_93_62 qb_93_62 bit_93_62 bitb_93_62 word93_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_62 q_94_62 qb_94_62 bit_94_62 bitb_94_62 word94_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_62 q_95_62 qb_95_62 bit_95_62 bitb_95_62 word95_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_62 q_96_62 qb_96_62 bit_96_62 bitb_96_62 word96_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_62 q_97_62 qb_97_62 bit_97_62 bitb_97_62 word97_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_62 q_98_62 qb_98_62 bit_98_62 bitb_98_62 word98_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_62 q_99_62 qb_99_62 bit_99_62 bitb_99_62 word99_62 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_63 q_0_63 qb_0_63 bit_0_63 bitb_0_63 word0_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_63 q_1_63 qb_1_63 bit_1_63 bitb_1_63 word1_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_63 q_2_63 qb_2_63 bit_2_63 bitb_2_63 word2_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_63 q_3_63 qb_3_63 bit_3_63 bitb_3_63 word3_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_63 q_4_63 qb_4_63 bit_4_63 bitb_4_63 word4_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_63 q_5_63 qb_5_63 bit_5_63 bitb_5_63 word5_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_63 q_6_63 qb_6_63 bit_6_63 bitb_6_63 word6_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_63 q_7_63 qb_7_63 bit_7_63 bitb_7_63 word7_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_63 q_8_63 qb_8_63 bit_8_63 bitb_8_63 word8_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_63 q_9_63 qb_9_63 bit_9_63 bitb_9_63 word9_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_63 q_10_63 qb_10_63 bit_10_63 bitb_10_63 word10_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_63 q_11_63 qb_11_63 bit_11_63 bitb_11_63 word11_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_63 q_12_63 qb_12_63 bit_12_63 bitb_12_63 word12_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_63 q_13_63 qb_13_63 bit_13_63 bitb_13_63 word13_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_63 q_14_63 qb_14_63 bit_14_63 bitb_14_63 word14_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_63 q_15_63 qb_15_63 bit_15_63 bitb_15_63 word15_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_63 q_16_63 qb_16_63 bit_16_63 bitb_16_63 word16_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_63 q_17_63 qb_17_63 bit_17_63 bitb_17_63 word17_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_63 q_18_63 qb_18_63 bit_18_63 bitb_18_63 word18_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_63 q_19_63 qb_19_63 bit_19_63 bitb_19_63 word19_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_63 q_20_63 qb_20_63 bit_20_63 bitb_20_63 word20_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_63 q_21_63 qb_21_63 bit_21_63 bitb_21_63 word21_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_63 q_22_63 qb_22_63 bit_22_63 bitb_22_63 word22_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_63 q_23_63 qb_23_63 bit_23_63 bitb_23_63 word23_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_63 q_24_63 qb_24_63 bit_24_63 bitb_24_63 word24_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_63 q_25_63 qb_25_63 bit_25_63 bitb_25_63 word25_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_63 q_26_63 qb_26_63 bit_26_63 bitb_26_63 word26_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_63 q_27_63 qb_27_63 bit_27_63 bitb_27_63 word27_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_63 q_28_63 qb_28_63 bit_28_63 bitb_28_63 word28_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_63 q_29_63 qb_29_63 bit_29_63 bitb_29_63 word29_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_63 q_30_63 qb_30_63 bit_30_63 bitb_30_63 word30_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_63 q_31_63 qb_31_63 bit_31_63 bitb_31_63 word31_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_63 q_32_63 qb_32_63 bit_32_63 bitb_32_63 word32_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_63 q_33_63 qb_33_63 bit_33_63 bitb_33_63 word33_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_63 q_34_63 qb_34_63 bit_34_63 bitb_34_63 word34_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_63 q_35_63 qb_35_63 bit_35_63 bitb_35_63 word35_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_63 q_36_63 qb_36_63 bit_36_63 bitb_36_63 word36_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_63 q_37_63 qb_37_63 bit_37_63 bitb_37_63 word37_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_63 q_38_63 qb_38_63 bit_38_63 bitb_38_63 word38_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_63 q_39_63 qb_39_63 bit_39_63 bitb_39_63 word39_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_63 q_40_63 qb_40_63 bit_40_63 bitb_40_63 word40_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_63 q_41_63 qb_41_63 bit_41_63 bitb_41_63 word41_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_63 q_42_63 qb_42_63 bit_42_63 bitb_42_63 word42_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_63 q_43_63 qb_43_63 bit_43_63 bitb_43_63 word43_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_63 q_44_63 qb_44_63 bit_44_63 bitb_44_63 word44_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_63 q_45_63 qb_45_63 bit_45_63 bitb_45_63 word45_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_63 q_46_63 qb_46_63 bit_46_63 bitb_46_63 word46_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_63 q_47_63 qb_47_63 bit_47_63 bitb_47_63 word47_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_63 q_48_63 qb_48_63 bit_48_63 bitb_48_63 word48_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_63 q_49_63 qb_49_63 bit_49_63 bitb_49_63 word49_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_63 q_50_63 qb_50_63 bit_50_63 bitb_50_63 word50_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_63 q_51_63 qb_51_63 bit_51_63 bitb_51_63 word51_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_63 q_52_63 qb_52_63 bit_52_63 bitb_52_63 word52_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_63 q_53_63 qb_53_63 bit_53_63 bitb_53_63 word53_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_63 q_54_63 qb_54_63 bit_54_63 bitb_54_63 word54_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_63 q_55_63 qb_55_63 bit_55_63 bitb_55_63 word55_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_63 q_56_63 qb_56_63 bit_56_63 bitb_56_63 word56_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_63 q_57_63 qb_57_63 bit_57_63 bitb_57_63 word57_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_63 q_58_63 qb_58_63 bit_58_63 bitb_58_63 word58_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_63 q_59_63 qb_59_63 bit_59_63 bitb_59_63 word59_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_63 q_60_63 qb_60_63 bit_60_63 bitb_60_63 word60_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_63 q_61_63 qb_61_63 bit_61_63 bitb_61_63 word61_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_63 q_62_63 qb_62_63 bit_62_63 bitb_62_63 word62_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_63 q_63_63 qb_63_63 bit_63_63 bitb_63_63 word63_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_63 q_64_63 qb_64_63 bit_64_63 bitb_64_63 word64_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_63 q_65_63 qb_65_63 bit_65_63 bitb_65_63 word65_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_63 q_66_63 qb_66_63 bit_66_63 bitb_66_63 word66_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_63 q_67_63 qb_67_63 bit_67_63 bitb_67_63 word67_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_63 q_68_63 qb_68_63 bit_68_63 bitb_68_63 word68_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_63 q_69_63 qb_69_63 bit_69_63 bitb_69_63 word69_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_63 q_70_63 qb_70_63 bit_70_63 bitb_70_63 word70_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_63 q_71_63 qb_71_63 bit_71_63 bitb_71_63 word71_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_63 q_72_63 qb_72_63 bit_72_63 bitb_72_63 word72_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_63 q_73_63 qb_73_63 bit_73_63 bitb_73_63 word73_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_63 q_74_63 qb_74_63 bit_74_63 bitb_74_63 word74_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_63 q_75_63 qb_75_63 bit_75_63 bitb_75_63 word75_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_63 q_76_63 qb_76_63 bit_76_63 bitb_76_63 word76_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_63 q_77_63 qb_77_63 bit_77_63 bitb_77_63 word77_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_63 q_78_63 qb_78_63 bit_78_63 bitb_78_63 word78_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_63 q_79_63 qb_79_63 bit_79_63 bitb_79_63 word79_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_63 q_80_63 qb_80_63 bit_80_63 bitb_80_63 word80_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_63 q_81_63 qb_81_63 bit_81_63 bitb_81_63 word81_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_63 q_82_63 qb_82_63 bit_82_63 bitb_82_63 word82_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_63 q_83_63 qb_83_63 bit_83_63 bitb_83_63 word83_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_63 q_84_63 qb_84_63 bit_84_63 bitb_84_63 word84_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_63 q_85_63 qb_85_63 bit_85_63 bitb_85_63 word85_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_63 q_86_63 qb_86_63 bit_86_63 bitb_86_63 word86_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_63 q_87_63 qb_87_63 bit_87_63 bitb_87_63 word87_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_63 q_88_63 qb_88_63 bit_88_63 bitb_88_63 word88_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_63 q_89_63 qb_89_63 bit_89_63 bitb_89_63 word89_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_63 q_90_63 qb_90_63 bit_90_63 bitb_90_63 word90_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_63 q_91_63 qb_91_63 bit_91_63 bitb_91_63 word91_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_63 q_92_63 qb_92_63 bit_92_63 bitb_92_63 word92_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_63 q_93_63 qb_93_63 bit_93_63 bitb_93_63 word93_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_63 q_94_63 qb_94_63 bit_94_63 bitb_94_63 word94_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_63 q_95_63 qb_95_63 bit_95_63 bitb_95_63 word95_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_63 q_96_63 qb_96_63 bit_96_63 bitb_96_63 word96_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_63 q_97_63 qb_97_63 bit_97_63 bitb_97_63 word97_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_63 q_98_63 qb_98_63 bit_98_63 bitb_98_63 word98_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_63 q_99_63 qb_99_63 bit_99_63 bitb_99_63 word99_63 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_64 q_0_64 qb_0_64 bit_0_64 bitb_0_64 word0_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_64 q_1_64 qb_1_64 bit_1_64 bitb_1_64 word1_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_64 q_2_64 qb_2_64 bit_2_64 bitb_2_64 word2_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_64 q_3_64 qb_3_64 bit_3_64 bitb_3_64 word3_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_64 q_4_64 qb_4_64 bit_4_64 bitb_4_64 word4_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_64 q_5_64 qb_5_64 bit_5_64 bitb_5_64 word5_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_64 q_6_64 qb_6_64 bit_6_64 bitb_6_64 word6_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_64 q_7_64 qb_7_64 bit_7_64 bitb_7_64 word7_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_64 q_8_64 qb_8_64 bit_8_64 bitb_8_64 word8_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_64 q_9_64 qb_9_64 bit_9_64 bitb_9_64 word9_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_64 q_10_64 qb_10_64 bit_10_64 bitb_10_64 word10_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_64 q_11_64 qb_11_64 bit_11_64 bitb_11_64 word11_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_64 q_12_64 qb_12_64 bit_12_64 bitb_12_64 word12_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_64 q_13_64 qb_13_64 bit_13_64 bitb_13_64 word13_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_64 q_14_64 qb_14_64 bit_14_64 bitb_14_64 word14_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_64 q_15_64 qb_15_64 bit_15_64 bitb_15_64 word15_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_64 q_16_64 qb_16_64 bit_16_64 bitb_16_64 word16_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_64 q_17_64 qb_17_64 bit_17_64 bitb_17_64 word17_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_64 q_18_64 qb_18_64 bit_18_64 bitb_18_64 word18_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_64 q_19_64 qb_19_64 bit_19_64 bitb_19_64 word19_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_64 q_20_64 qb_20_64 bit_20_64 bitb_20_64 word20_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_64 q_21_64 qb_21_64 bit_21_64 bitb_21_64 word21_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_64 q_22_64 qb_22_64 bit_22_64 bitb_22_64 word22_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_64 q_23_64 qb_23_64 bit_23_64 bitb_23_64 word23_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_64 q_24_64 qb_24_64 bit_24_64 bitb_24_64 word24_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_64 q_25_64 qb_25_64 bit_25_64 bitb_25_64 word25_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_64 q_26_64 qb_26_64 bit_26_64 bitb_26_64 word26_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_64 q_27_64 qb_27_64 bit_27_64 bitb_27_64 word27_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_64 q_28_64 qb_28_64 bit_28_64 bitb_28_64 word28_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_64 q_29_64 qb_29_64 bit_29_64 bitb_29_64 word29_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_64 q_30_64 qb_30_64 bit_30_64 bitb_30_64 word30_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_64 q_31_64 qb_31_64 bit_31_64 bitb_31_64 word31_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_64 q_32_64 qb_32_64 bit_32_64 bitb_32_64 word32_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_64 q_33_64 qb_33_64 bit_33_64 bitb_33_64 word33_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_64 q_34_64 qb_34_64 bit_34_64 bitb_34_64 word34_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_64 q_35_64 qb_35_64 bit_35_64 bitb_35_64 word35_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_64 q_36_64 qb_36_64 bit_36_64 bitb_36_64 word36_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_64 q_37_64 qb_37_64 bit_37_64 bitb_37_64 word37_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_64 q_38_64 qb_38_64 bit_38_64 bitb_38_64 word38_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_64 q_39_64 qb_39_64 bit_39_64 bitb_39_64 word39_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_64 q_40_64 qb_40_64 bit_40_64 bitb_40_64 word40_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_64 q_41_64 qb_41_64 bit_41_64 bitb_41_64 word41_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_64 q_42_64 qb_42_64 bit_42_64 bitb_42_64 word42_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_64 q_43_64 qb_43_64 bit_43_64 bitb_43_64 word43_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_64 q_44_64 qb_44_64 bit_44_64 bitb_44_64 word44_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_64 q_45_64 qb_45_64 bit_45_64 bitb_45_64 word45_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_64 q_46_64 qb_46_64 bit_46_64 bitb_46_64 word46_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_64 q_47_64 qb_47_64 bit_47_64 bitb_47_64 word47_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_64 q_48_64 qb_48_64 bit_48_64 bitb_48_64 word48_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_64 q_49_64 qb_49_64 bit_49_64 bitb_49_64 word49_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_64 q_50_64 qb_50_64 bit_50_64 bitb_50_64 word50_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_64 q_51_64 qb_51_64 bit_51_64 bitb_51_64 word51_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_64 q_52_64 qb_52_64 bit_52_64 bitb_52_64 word52_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_64 q_53_64 qb_53_64 bit_53_64 bitb_53_64 word53_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_64 q_54_64 qb_54_64 bit_54_64 bitb_54_64 word54_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_64 q_55_64 qb_55_64 bit_55_64 bitb_55_64 word55_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_64 q_56_64 qb_56_64 bit_56_64 bitb_56_64 word56_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_64 q_57_64 qb_57_64 bit_57_64 bitb_57_64 word57_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_64 q_58_64 qb_58_64 bit_58_64 bitb_58_64 word58_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_64 q_59_64 qb_59_64 bit_59_64 bitb_59_64 word59_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_64 q_60_64 qb_60_64 bit_60_64 bitb_60_64 word60_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_64 q_61_64 qb_61_64 bit_61_64 bitb_61_64 word61_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_64 q_62_64 qb_62_64 bit_62_64 bitb_62_64 word62_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_64 q_63_64 qb_63_64 bit_63_64 bitb_63_64 word63_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_64 q_64_64 qb_64_64 bit_64_64 bitb_64_64 word64_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_64 q_65_64 qb_65_64 bit_65_64 bitb_65_64 word65_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_64 q_66_64 qb_66_64 bit_66_64 bitb_66_64 word66_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_64 q_67_64 qb_67_64 bit_67_64 bitb_67_64 word67_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_64 q_68_64 qb_68_64 bit_68_64 bitb_68_64 word68_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_64 q_69_64 qb_69_64 bit_69_64 bitb_69_64 word69_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_64 q_70_64 qb_70_64 bit_70_64 bitb_70_64 word70_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_64 q_71_64 qb_71_64 bit_71_64 bitb_71_64 word71_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_64 q_72_64 qb_72_64 bit_72_64 bitb_72_64 word72_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_64 q_73_64 qb_73_64 bit_73_64 bitb_73_64 word73_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_64 q_74_64 qb_74_64 bit_74_64 bitb_74_64 word74_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_64 q_75_64 qb_75_64 bit_75_64 bitb_75_64 word75_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_64 q_76_64 qb_76_64 bit_76_64 bitb_76_64 word76_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_64 q_77_64 qb_77_64 bit_77_64 bitb_77_64 word77_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_64 q_78_64 qb_78_64 bit_78_64 bitb_78_64 word78_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_64 q_79_64 qb_79_64 bit_79_64 bitb_79_64 word79_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_64 q_80_64 qb_80_64 bit_80_64 bitb_80_64 word80_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_64 q_81_64 qb_81_64 bit_81_64 bitb_81_64 word81_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_64 q_82_64 qb_82_64 bit_82_64 bitb_82_64 word82_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_64 q_83_64 qb_83_64 bit_83_64 bitb_83_64 word83_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_64 q_84_64 qb_84_64 bit_84_64 bitb_84_64 word84_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_64 q_85_64 qb_85_64 bit_85_64 bitb_85_64 word85_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_64 q_86_64 qb_86_64 bit_86_64 bitb_86_64 word86_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_64 q_87_64 qb_87_64 bit_87_64 bitb_87_64 word87_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_64 q_88_64 qb_88_64 bit_88_64 bitb_88_64 word88_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_64 q_89_64 qb_89_64 bit_89_64 bitb_89_64 word89_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_64 q_90_64 qb_90_64 bit_90_64 bitb_90_64 word90_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_64 q_91_64 qb_91_64 bit_91_64 bitb_91_64 word91_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_64 q_92_64 qb_92_64 bit_92_64 bitb_92_64 word92_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_64 q_93_64 qb_93_64 bit_93_64 bitb_93_64 word93_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_64 q_94_64 qb_94_64 bit_94_64 bitb_94_64 word94_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_64 q_95_64 qb_95_64 bit_95_64 bitb_95_64 word95_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_64 q_96_64 qb_96_64 bit_96_64 bitb_96_64 word96_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_64 q_97_64 qb_97_64 bit_97_64 bitb_97_64 word97_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_64 q_98_64 qb_98_64 bit_98_64 bitb_98_64 word98_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_64 q_99_64 qb_99_64 bit_99_64 bitb_99_64 word99_64 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_65 q_0_65 qb_0_65 bit_0_65 bitb_0_65 word0_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_65 q_1_65 qb_1_65 bit_1_65 bitb_1_65 word1_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_65 q_2_65 qb_2_65 bit_2_65 bitb_2_65 word2_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_65 q_3_65 qb_3_65 bit_3_65 bitb_3_65 word3_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_65 q_4_65 qb_4_65 bit_4_65 bitb_4_65 word4_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_65 q_5_65 qb_5_65 bit_5_65 bitb_5_65 word5_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_65 q_6_65 qb_6_65 bit_6_65 bitb_6_65 word6_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_65 q_7_65 qb_7_65 bit_7_65 bitb_7_65 word7_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_65 q_8_65 qb_8_65 bit_8_65 bitb_8_65 word8_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_65 q_9_65 qb_9_65 bit_9_65 bitb_9_65 word9_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_65 q_10_65 qb_10_65 bit_10_65 bitb_10_65 word10_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_65 q_11_65 qb_11_65 bit_11_65 bitb_11_65 word11_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_65 q_12_65 qb_12_65 bit_12_65 bitb_12_65 word12_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_65 q_13_65 qb_13_65 bit_13_65 bitb_13_65 word13_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_65 q_14_65 qb_14_65 bit_14_65 bitb_14_65 word14_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_65 q_15_65 qb_15_65 bit_15_65 bitb_15_65 word15_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_65 q_16_65 qb_16_65 bit_16_65 bitb_16_65 word16_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_65 q_17_65 qb_17_65 bit_17_65 bitb_17_65 word17_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_65 q_18_65 qb_18_65 bit_18_65 bitb_18_65 word18_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_65 q_19_65 qb_19_65 bit_19_65 bitb_19_65 word19_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_65 q_20_65 qb_20_65 bit_20_65 bitb_20_65 word20_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_65 q_21_65 qb_21_65 bit_21_65 bitb_21_65 word21_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_65 q_22_65 qb_22_65 bit_22_65 bitb_22_65 word22_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_65 q_23_65 qb_23_65 bit_23_65 bitb_23_65 word23_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_65 q_24_65 qb_24_65 bit_24_65 bitb_24_65 word24_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_65 q_25_65 qb_25_65 bit_25_65 bitb_25_65 word25_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_65 q_26_65 qb_26_65 bit_26_65 bitb_26_65 word26_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_65 q_27_65 qb_27_65 bit_27_65 bitb_27_65 word27_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_65 q_28_65 qb_28_65 bit_28_65 bitb_28_65 word28_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_65 q_29_65 qb_29_65 bit_29_65 bitb_29_65 word29_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_65 q_30_65 qb_30_65 bit_30_65 bitb_30_65 word30_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_65 q_31_65 qb_31_65 bit_31_65 bitb_31_65 word31_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_65 q_32_65 qb_32_65 bit_32_65 bitb_32_65 word32_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_65 q_33_65 qb_33_65 bit_33_65 bitb_33_65 word33_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_65 q_34_65 qb_34_65 bit_34_65 bitb_34_65 word34_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_65 q_35_65 qb_35_65 bit_35_65 bitb_35_65 word35_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_65 q_36_65 qb_36_65 bit_36_65 bitb_36_65 word36_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_65 q_37_65 qb_37_65 bit_37_65 bitb_37_65 word37_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_65 q_38_65 qb_38_65 bit_38_65 bitb_38_65 word38_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_65 q_39_65 qb_39_65 bit_39_65 bitb_39_65 word39_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_65 q_40_65 qb_40_65 bit_40_65 bitb_40_65 word40_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_65 q_41_65 qb_41_65 bit_41_65 bitb_41_65 word41_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_65 q_42_65 qb_42_65 bit_42_65 bitb_42_65 word42_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_65 q_43_65 qb_43_65 bit_43_65 bitb_43_65 word43_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_65 q_44_65 qb_44_65 bit_44_65 bitb_44_65 word44_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_65 q_45_65 qb_45_65 bit_45_65 bitb_45_65 word45_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_65 q_46_65 qb_46_65 bit_46_65 bitb_46_65 word46_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_65 q_47_65 qb_47_65 bit_47_65 bitb_47_65 word47_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_65 q_48_65 qb_48_65 bit_48_65 bitb_48_65 word48_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_65 q_49_65 qb_49_65 bit_49_65 bitb_49_65 word49_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_65 q_50_65 qb_50_65 bit_50_65 bitb_50_65 word50_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_65 q_51_65 qb_51_65 bit_51_65 bitb_51_65 word51_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_65 q_52_65 qb_52_65 bit_52_65 bitb_52_65 word52_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_65 q_53_65 qb_53_65 bit_53_65 bitb_53_65 word53_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_65 q_54_65 qb_54_65 bit_54_65 bitb_54_65 word54_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_65 q_55_65 qb_55_65 bit_55_65 bitb_55_65 word55_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_65 q_56_65 qb_56_65 bit_56_65 bitb_56_65 word56_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_65 q_57_65 qb_57_65 bit_57_65 bitb_57_65 word57_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_65 q_58_65 qb_58_65 bit_58_65 bitb_58_65 word58_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_65 q_59_65 qb_59_65 bit_59_65 bitb_59_65 word59_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_65 q_60_65 qb_60_65 bit_60_65 bitb_60_65 word60_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_65 q_61_65 qb_61_65 bit_61_65 bitb_61_65 word61_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_65 q_62_65 qb_62_65 bit_62_65 bitb_62_65 word62_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_65 q_63_65 qb_63_65 bit_63_65 bitb_63_65 word63_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_65 q_64_65 qb_64_65 bit_64_65 bitb_64_65 word64_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_65 q_65_65 qb_65_65 bit_65_65 bitb_65_65 word65_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_65 q_66_65 qb_66_65 bit_66_65 bitb_66_65 word66_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_65 q_67_65 qb_67_65 bit_67_65 bitb_67_65 word67_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_65 q_68_65 qb_68_65 bit_68_65 bitb_68_65 word68_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_65 q_69_65 qb_69_65 bit_69_65 bitb_69_65 word69_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_65 q_70_65 qb_70_65 bit_70_65 bitb_70_65 word70_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_65 q_71_65 qb_71_65 bit_71_65 bitb_71_65 word71_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_65 q_72_65 qb_72_65 bit_72_65 bitb_72_65 word72_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_65 q_73_65 qb_73_65 bit_73_65 bitb_73_65 word73_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_65 q_74_65 qb_74_65 bit_74_65 bitb_74_65 word74_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_65 q_75_65 qb_75_65 bit_75_65 bitb_75_65 word75_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_65 q_76_65 qb_76_65 bit_76_65 bitb_76_65 word76_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_65 q_77_65 qb_77_65 bit_77_65 bitb_77_65 word77_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_65 q_78_65 qb_78_65 bit_78_65 bitb_78_65 word78_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_65 q_79_65 qb_79_65 bit_79_65 bitb_79_65 word79_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_65 q_80_65 qb_80_65 bit_80_65 bitb_80_65 word80_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_65 q_81_65 qb_81_65 bit_81_65 bitb_81_65 word81_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_65 q_82_65 qb_82_65 bit_82_65 bitb_82_65 word82_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_65 q_83_65 qb_83_65 bit_83_65 bitb_83_65 word83_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_65 q_84_65 qb_84_65 bit_84_65 bitb_84_65 word84_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_65 q_85_65 qb_85_65 bit_85_65 bitb_85_65 word85_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_65 q_86_65 qb_86_65 bit_86_65 bitb_86_65 word86_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_65 q_87_65 qb_87_65 bit_87_65 bitb_87_65 word87_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_65 q_88_65 qb_88_65 bit_88_65 bitb_88_65 word88_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_65 q_89_65 qb_89_65 bit_89_65 bitb_89_65 word89_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_65 q_90_65 qb_90_65 bit_90_65 bitb_90_65 word90_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_65 q_91_65 qb_91_65 bit_91_65 bitb_91_65 word91_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_65 q_92_65 qb_92_65 bit_92_65 bitb_92_65 word92_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_65 q_93_65 qb_93_65 bit_93_65 bitb_93_65 word93_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_65 q_94_65 qb_94_65 bit_94_65 bitb_94_65 word94_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_65 q_95_65 qb_95_65 bit_95_65 bitb_95_65 word95_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_65 q_96_65 qb_96_65 bit_96_65 bitb_96_65 word96_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_65 q_97_65 qb_97_65 bit_97_65 bitb_97_65 word97_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_65 q_98_65 qb_98_65 bit_98_65 bitb_98_65 word98_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_65 q_99_65 qb_99_65 bit_99_65 bitb_99_65 word99_65 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_66 q_0_66 qb_0_66 bit_0_66 bitb_0_66 word0_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_66 q_1_66 qb_1_66 bit_1_66 bitb_1_66 word1_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_66 q_2_66 qb_2_66 bit_2_66 bitb_2_66 word2_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_66 q_3_66 qb_3_66 bit_3_66 bitb_3_66 word3_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_66 q_4_66 qb_4_66 bit_4_66 bitb_4_66 word4_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_66 q_5_66 qb_5_66 bit_5_66 bitb_5_66 word5_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_66 q_6_66 qb_6_66 bit_6_66 bitb_6_66 word6_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_66 q_7_66 qb_7_66 bit_7_66 bitb_7_66 word7_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_66 q_8_66 qb_8_66 bit_8_66 bitb_8_66 word8_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_66 q_9_66 qb_9_66 bit_9_66 bitb_9_66 word9_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_66 q_10_66 qb_10_66 bit_10_66 bitb_10_66 word10_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_66 q_11_66 qb_11_66 bit_11_66 bitb_11_66 word11_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_66 q_12_66 qb_12_66 bit_12_66 bitb_12_66 word12_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_66 q_13_66 qb_13_66 bit_13_66 bitb_13_66 word13_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_66 q_14_66 qb_14_66 bit_14_66 bitb_14_66 word14_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_66 q_15_66 qb_15_66 bit_15_66 bitb_15_66 word15_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_66 q_16_66 qb_16_66 bit_16_66 bitb_16_66 word16_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_66 q_17_66 qb_17_66 bit_17_66 bitb_17_66 word17_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_66 q_18_66 qb_18_66 bit_18_66 bitb_18_66 word18_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_66 q_19_66 qb_19_66 bit_19_66 bitb_19_66 word19_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_66 q_20_66 qb_20_66 bit_20_66 bitb_20_66 word20_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_66 q_21_66 qb_21_66 bit_21_66 bitb_21_66 word21_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_66 q_22_66 qb_22_66 bit_22_66 bitb_22_66 word22_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_66 q_23_66 qb_23_66 bit_23_66 bitb_23_66 word23_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_66 q_24_66 qb_24_66 bit_24_66 bitb_24_66 word24_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_66 q_25_66 qb_25_66 bit_25_66 bitb_25_66 word25_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_66 q_26_66 qb_26_66 bit_26_66 bitb_26_66 word26_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_66 q_27_66 qb_27_66 bit_27_66 bitb_27_66 word27_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_66 q_28_66 qb_28_66 bit_28_66 bitb_28_66 word28_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_66 q_29_66 qb_29_66 bit_29_66 bitb_29_66 word29_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_66 q_30_66 qb_30_66 bit_30_66 bitb_30_66 word30_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_66 q_31_66 qb_31_66 bit_31_66 bitb_31_66 word31_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_66 q_32_66 qb_32_66 bit_32_66 bitb_32_66 word32_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_66 q_33_66 qb_33_66 bit_33_66 bitb_33_66 word33_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_66 q_34_66 qb_34_66 bit_34_66 bitb_34_66 word34_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_66 q_35_66 qb_35_66 bit_35_66 bitb_35_66 word35_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_66 q_36_66 qb_36_66 bit_36_66 bitb_36_66 word36_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_66 q_37_66 qb_37_66 bit_37_66 bitb_37_66 word37_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_66 q_38_66 qb_38_66 bit_38_66 bitb_38_66 word38_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_66 q_39_66 qb_39_66 bit_39_66 bitb_39_66 word39_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_66 q_40_66 qb_40_66 bit_40_66 bitb_40_66 word40_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_66 q_41_66 qb_41_66 bit_41_66 bitb_41_66 word41_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_66 q_42_66 qb_42_66 bit_42_66 bitb_42_66 word42_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_66 q_43_66 qb_43_66 bit_43_66 bitb_43_66 word43_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_66 q_44_66 qb_44_66 bit_44_66 bitb_44_66 word44_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_66 q_45_66 qb_45_66 bit_45_66 bitb_45_66 word45_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_66 q_46_66 qb_46_66 bit_46_66 bitb_46_66 word46_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_66 q_47_66 qb_47_66 bit_47_66 bitb_47_66 word47_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_66 q_48_66 qb_48_66 bit_48_66 bitb_48_66 word48_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_66 q_49_66 qb_49_66 bit_49_66 bitb_49_66 word49_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_66 q_50_66 qb_50_66 bit_50_66 bitb_50_66 word50_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_66 q_51_66 qb_51_66 bit_51_66 bitb_51_66 word51_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_66 q_52_66 qb_52_66 bit_52_66 bitb_52_66 word52_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_66 q_53_66 qb_53_66 bit_53_66 bitb_53_66 word53_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_66 q_54_66 qb_54_66 bit_54_66 bitb_54_66 word54_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_66 q_55_66 qb_55_66 bit_55_66 bitb_55_66 word55_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_66 q_56_66 qb_56_66 bit_56_66 bitb_56_66 word56_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_66 q_57_66 qb_57_66 bit_57_66 bitb_57_66 word57_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_66 q_58_66 qb_58_66 bit_58_66 bitb_58_66 word58_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_66 q_59_66 qb_59_66 bit_59_66 bitb_59_66 word59_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_66 q_60_66 qb_60_66 bit_60_66 bitb_60_66 word60_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_66 q_61_66 qb_61_66 bit_61_66 bitb_61_66 word61_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_66 q_62_66 qb_62_66 bit_62_66 bitb_62_66 word62_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_66 q_63_66 qb_63_66 bit_63_66 bitb_63_66 word63_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_66 q_64_66 qb_64_66 bit_64_66 bitb_64_66 word64_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_66 q_65_66 qb_65_66 bit_65_66 bitb_65_66 word65_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_66 q_66_66 qb_66_66 bit_66_66 bitb_66_66 word66_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_66 q_67_66 qb_67_66 bit_67_66 bitb_67_66 word67_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_66 q_68_66 qb_68_66 bit_68_66 bitb_68_66 word68_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_66 q_69_66 qb_69_66 bit_69_66 bitb_69_66 word69_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_66 q_70_66 qb_70_66 bit_70_66 bitb_70_66 word70_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_66 q_71_66 qb_71_66 bit_71_66 bitb_71_66 word71_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_66 q_72_66 qb_72_66 bit_72_66 bitb_72_66 word72_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_66 q_73_66 qb_73_66 bit_73_66 bitb_73_66 word73_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_66 q_74_66 qb_74_66 bit_74_66 bitb_74_66 word74_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_66 q_75_66 qb_75_66 bit_75_66 bitb_75_66 word75_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_66 q_76_66 qb_76_66 bit_76_66 bitb_76_66 word76_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_66 q_77_66 qb_77_66 bit_77_66 bitb_77_66 word77_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_66 q_78_66 qb_78_66 bit_78_66 bitb_78_66 word78_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_66 q_79_66 qb_79_66 bit_79_66 bitb_79_66 word79_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_66 q_80_66 qb_80_66 bit_80_66 bitb_80_66 word80_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_66 q_81_66 qb_81_66 bit_81_66 bitb_81_66 word81_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_66 q_82_66 qb_82_66 bit_82_66 bitb_82_66 word82_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_66 q_83_66 qb_83_66 bit_83_66 bitb_83_66 word83_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_66 q_84_66 qb_84_66 bit_84_66 bitb_84_66 word84_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_66 q_85_66 qb_85_66 bit_85_66 bitb_85_66 word85_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_66 q_86_66 qb_86_66 bit_86_66 bitb_86_66 word86_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_66 q_87_66 qb_87_66 bit_87_66 bitb_87_66 word87_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_66 q_88_66 qb_88_66 bit_88_66 bitb_88_66 word88_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_66 q_89_66 qb_89_66 bit_89_66 bitb_89_66 word89_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_66 q_90_66 qb_90_66 bit_90_66 bitb_90_66 word90_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_66 q_91_66 qb_91_66 bit_91_66 bitb_91_66 word91_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_66 q_92_66 qb_92_66 bit_92_66 bitb_92_66 word92_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_66 q_93_66 qb_93_66 bit_93_66 bitb_93_66 word93_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_66 q_94_66 qb_94_66 bit_94_66 bitb_94_66 word94_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_66 q_95_66 qb_95_66 bit_95_66 bitb_95_66 word95_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_66 q_96_66 qb_96_66 bit_96_66 bitb_96_66 word96_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_66 q_97_66 qb_97_66 bit_97_66 bitb_97_66 word97_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_66 q_98_66 qb_98_66 bit_98_66 bitb_98_66 word98_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_66 q_99_66 qb_99_66 bit_99_66 bitb_99_66 word99_66 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_67 q_0_67 qb_0_67 bit_0_67 bitb_0_67 word0_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_67 q_1_67 qb_1_67 bit_1_67 bitb_1_67 word1_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_67 q_2_67 qb_2_67 bit_2_67 bitb_2_67 word2_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_67 q_3_67 qb_3_67 bit_3_67 bitb_3_67 word3_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_67 q_4_67 qb_4_67 bit_4_67 bitb_4_67 word4_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_67 q_5_67 qb_5_67 bit_5_67 bitb_5_67 word5_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_67 q_6_67 qb_6_67 bit_6_67 bitb_6_67 word6_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_67 q_7_67 qb_7_67 bit_7_67 bitb_7_67 word7_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_67 q_8_67 qb_8_67 bit_8_67 bitb_8_67 word8_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_67 q_9_67 qb_9_67 bit_9_67 bitb_9_67 word9_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_67 q_10_67 qb_10_67 bit_10_67 bitb_10_67 word10_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_67 q_11_67 qb_11_67 bit_11_67 bitb_11_67 word11_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_67 q_12_67 qb_12_67 bit_12_67 bitb_12_67 word12_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_67 q_13_67 qb_13_67 bit_13_67 bitb_13_67 word13_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_67 q_14_67 qb_14_67 bit_14_67 bitb_14_67 word14_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_67 q_15_67 qb_15_67 bit_15_67 bitb_15_67 word15_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_67 q_16_67 qb_16_67 bit_16_67 bitb_16_67 word16_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_67 q_17_67 qb_17_67 bit_17_67 bitb_17_67 word17_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_67 q_18_67 qb_18_67 bit_18_67 bitb_18_67 word18_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_67 q_19_67 qb_19_67 bit_19_67 bitb_19_67 word19_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_67 q_20_67 qb_20_67 bit_20_67 bitb_20_67 word20_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_67 q_21_67 qb_21_67 bit_21_67 bitb_21_67 word21_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_67 q_22_67 qb_22_67 bit_22_67 bitb_22_67 word22_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_67 q_23_67 qb_23_67 bit_23_67 bitb_23_67 word23_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_67 q_24_67 qb_24_67 bit_24_67 bitb_24_67 word24_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_67 q_25_67 qb_25_67 bit_25_67 bitb_25_67 word25_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_67 q_26_67 qb_26_67 bit_26_67 bitb_26_67 word26_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_67 q_27_67 qb_27_67 bit_27_67 bitb_27_67 word27_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_67 q_28_67 qb_28_67 bit_28_67 bitb_28_67 word28_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_67 q_29_67 qb_29_67 bit_29_67 bitb_29_67 word29_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_67 q_30_67 qb_30_67 bit_30_67 bitb_30_67 word30_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_67 q_31_67 qb_31_67 bit_31_67 bitb_31_67 word31_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_67 q_32_67 qb_32_67 bit_32_67 bitb_32_67 word32_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_67 q_33_67 qb_33_67 bit_33_67 bitb_33_67 word33_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_67 q_34_67 qb_34_67 bit_34_67 bitb_34_67 word34_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_67 q_35_67 qb_35_67 bit_35_67 bitb_35_67 word35_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_67 q_36_67 qb_36_67 bit_36_67 bitb_36_67 word36_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_67 q_37_67 qb_37_67 bit_37_67 bitb_37_67 word37_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_67 q_38_67 qb_38_67 bit_38_67 bitb_38_67 word38_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_67 q_39_67 qb_39_67 bit_39_67 bitb_39_67 word39_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_67 q_40_67 qb_40_67 bit_40_67 bitb_40_67 word40_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_67 q_41_67 qb_41_67 bit_41_67 bitb_41_67 word41_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_67 q_42_67 qb_42_67 bit_42_67 bitb_42_67 word42_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_67 q_43_67 qb_43_67 bit_43_67 bitb_43_67 word43_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_67 q_44_67 qb_44_67 bit_44_67 bitb_44_67 word44_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_67 q_45_67 qb_45_67 bit_45_67 bitb_45_67 word45_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_67 q_46_67 qb_46_67 bit_46_67 bitb_46_67 word46_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_67 q_47_67 qb_47_67 bit_47_67 bitb_47_67 word47_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_67 q_48_67 qb_48_67 bit_48_67 bitb_48_67 word48_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_67 q_49_67 qb_49_67 bit_49_67 bitb_49_67 word49_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_67 q_50_67 qb_50_67 bit_50_67 bitb_50_67 word50_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_67 q_51_67 qb_51_67 bit_51_67 bitb_51_67 word51_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_67 q_52_67 qb_52_67 bit_52_67 bitb_52_67 word52_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_67 q_53_67 qb_53_67 bit_53_67 bitb_53_67 word53_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_67 q_54_67 qb_54_67 bit_54_67 bitb_54_67 word54_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_67 q_55_67 qb_55_67 bit_55_67 bitb_55_67 word55_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_67 q_56_67 qb_56_67 bit_56_67 bitb_56_67 word56_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_67 q_57_67 qb_57_67 bit_57_67 bitb_57_67 word57_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_67 q_58_67 qb_58_67 bit_58_67 bitb_58_67 word58_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_67 q_59_67 qb_59_67 bit_59_67 bitb_59_67 word59_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_67 q_60_67 qb_60_67 bit_60_67 bitb_60_67 word60_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_67 q_61_67 qb_61_67 bit_61_67 bitb_61_67 word61_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_67 q_62_67 qb_62_67 bit_62_67 bitb_62_67 word62_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_67 q_63_67 qb_63_67 bit_63_67 bitb_63_67 word63_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_67 q_64_67 qb_64_67 bit_64_67 bitb_64_67 word64_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_67 q_65_67 qb_65_67 bit_65_67 bitb_65_67 word65_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_67 q_66_67 qb_66_67 bit_66_67 bitb_66_67 word66_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_67 q_67_67 qb_67_67 bit_67_67 bitb_67_67 word67_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_67 q_68_67 qb_68_67 bit_68_67 bitb_68_67 word68_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_67 q_69_67 qb_69_67 bit_69_67 bitb_69_67 word69_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_67 q_70_67 qb_70_67 bit_70_67 bitb_70_67 word70_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_67 q_71_67 qb_71_67 bit_71_67 bitb_71_67 word71_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_67 q_72_67 qb_72_67 bit_72_67 bitb_72_67 word72_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_67 q_73_67 qb_73_67 bit_73_67 bitb_73_67 word73_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_67 q_74_67 qb_74_67 bit_74_67 bitb_74_67 word74_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_67 q_75_67 qb_75_67 bit_75_67 bitb_75_67 word75_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_67 q_76_67 qb_76_67 bit_76_67 bitb_76_67 word76_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_67 q_77_67 qb_77_67 bit_77_67 bitb_77_67 word77_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_67 q_78_67 qb_78_67 bit_78_67 bitb_78_67 word78_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_67 q_79_67 qb_79_67 bit_79_67 bitb_79_67 word79_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_67 q_80_67 qb_80_67 bit_80_67 bitb_80_67 word80_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_67 q_81_67 qb_81_67 bit_81_67 bitb_81_67 word81_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_67 q_82_67 qb_82_67 bit_82_67 bitb_82_67 word82_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_67 q_83_67 qb_83_67 bit_83_67 bitb_83_67 word83_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_67 q_84_67 qb_84_67 bit_84_67 bitb_84_67 word84_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_67 q_85_67 qb_85_67 bit_85_67 bitb_85_67 word85_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_67 q_86_67 qb_86_67 bit_86_67 bitb_86_67 word86_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_67 q_87_67 qb_87_67 bit_87_67 bitb_87_67 word87_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_67 q_88_67 qb_88_67 bit_88_67 bitb_88_67 word88_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_67 q_89_67 qb_89_67 bit_89_67 bitb_89_67 word89_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_67 q_90_67 qb_90_67 bit_90_67 bitb_90_67 word90_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_67 q_91_67 qb_91_67 bit_91_67 bitb_91_67 word91_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_67 q_92_67 qb_92_67 bit_92_67 bitb_92_67 word92_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_67 q_93_67 qb_93_67 bit_93_67 bitb_93_67 word93_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_67 q_94_67 qb_94_67 bit_94_67 bitb_94_67 word94_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_67 q_95_67 qb_95_67 bit_95_67 bitb_95_67 word95_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_67 q_96_67 qb_96_67 bit_96_67 bitb_96_67 word96_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_67 q_97_67 qb_97_67 bit_97_67 bitb_97_67 word97_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_67 q_98_67 qb_98_67 bit_98_67 bitb_98_67 word98_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_67 q_99_67 qb_99_67 bit_99_67 bitb_99_67 word99_67 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_68 q_0_68 qb_0_68 bit_0_68 bitb_0_68 word0_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_68 q_1_68 qb_1_68 bit_1_68 bitb_1_68 word1_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_68 q_2_68 qb_2_68 bit_2_68 bitb_2_68 word2_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_68 q_3_68 qb_3_68 bit_3_68 bitb_3_68 word3_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_68 q_4_68 qb_4_68 bit_4_68 bitb_4_68 word4_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_68 q_5_68 qb_5_68 bit_5_68 bitb_5_68 word5_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_68 q_6_68 qb_6_68 bit_6_68 bitb_6_68 word6_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_68 q_7_68 qb_7_68 bit_7_68 bitb_7_68 word7_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_68 q_8_68 qb_8_68 bit_8_68 bitb_8_68 word8_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_68 q_9_68 qb_9_68 bit_9_68 bitb_9_68 word9_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_68 q_10_68 qb_10_68 bit_10_68 bitb_10_68 word10_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_68 q_11_68 qb_11_68 bit_11_68 bitb_11_68 word11_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_68 q_12_68 qb_12_68 bit_12_68 bitb_12_68 word12_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_68 q_13_68 qb_13_68 bit_13_68 bitb_13_68 word13_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_68 q_14_68 qb_14_68 bit_14_68 bitb_14_68 word14_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_68 q_15_68 qb_15_68 bit_15_68 bitb_15_68 word15_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_68 q_16_68 qb_16_68 bit_16_68 bitb_16_68 word16_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_68 q_17_68 qb_17_68 bit_17_68 bitb_17_68 word17_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_68 q_18_68 qb_18_68 bit_18_68 bitb_18_68 word18_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_68 q_19_68 qb_19_68 bit_19_68 bitb_19_68 word19_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_68 q_20_68 qb_20_68 bit_20_68 bitb_20_68 word20_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_68 q_21_68 qb_21_68 bit_21_68 bitb_21_68 word21_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_68 q_22_68 qb_22_68 bit_22_68 bitb_22_68 word22_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_68 q_23_68 qb_23_68 bit_23_68 bitb_23_68 word23_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_68 q_24_68 qb_24_68 bit_24_68 bitb_24_68 word24_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_68 q_25_68 qb_25_68 bit_25_68 bitb_25_68 word25_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_68 q_26_68 qb_26_68 bit_26_68 bitb_26_68 word26_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_68 q_27_68 qb_27_68 bit_27_68 bitb_27_68 word27_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_68 q_28_68 qb_28_68 bit_28_68 bitb_28_68 word28_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_68 q_29_68 qb_29_68 bit_29_68 bitb_29_68 word29_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_68 q_30_68 qb_30_68 bit_30_68 bitb_30_68 word30_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_68 q_31_68 qb_31_68 bit_31_68 bitb_31_68 word31_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_68 q_32_68 qb_32_68 bit_32_68 bitb_32_68 word32_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_68 q_33_68 qb_33_68 bit_33_68 bitb_33_68 word33_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_68 q_34_68 qb_34_68 bit_34_68 bitb_34_68 word34_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_68 q_35_68 qb_35_68 bit_35_68 bitb_35_68 word35_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_68 q_36_68 qb_36_68 bit_36_68 bitb_36_68 word36_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_68 q_37_68 qb_37_68 bit_37_68 bitb_37_68 word37_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_68 q_38_68 qb_38_68 bit_38_68 bitb_38_68 word38_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_68 q_39_68 qb_39_68 bit_39_68 bitb_39_68 word39_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_68 q_40_68 qb_40_68 bit_40_68 bitb_40_68 word40_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_68 q_41_68 qb_41_68 bit_41_68 bitb_41_68 word41_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_68 q_42_68 qb_42_68 bit_42_68 bitb_42_68 word42_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_68 q_43_68 qb_43_68 bit_43_68 bitb_43_68 word43_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_68 q_44_68 qb_44_68 bit_44_68 bitb_44_68 word44_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_68 q_45_68 qb_45_68 bit_45_68 bitb_45_68 word45_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_68 q_46_68 qb_46_68 bit_46_68 bitb_46_68 word46_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_68 q_47_68 qb_47_68 bit_47_68 bitb_47_68 word47_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_68 q_48_68 qb_48_68 bit_48_68 bitb_48_68 word48_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_68 q_49_68 qb_49_68 bit_49_68 bitb_49_68 word49_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_68 q_50_68 qb_50_68 bit_50_68 bitb_50_68 word50_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_68 q_51_68 qb_51_68 bit_51_68 bitb_51_68 word51_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_68 q_52_68 qb_52_68 bit_52_68 bitb_52_68 word52_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_68 q_53_68 qb_53_68 bit_53_68 bitb_53_68 word53_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_68 q_54_68 qb_54_68 bit_54_68 bitb_54_68 word54_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_68 q_55_68 qb_55_68 bit_55_68 bitb_55_68 word55_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_68 q_56_68 qb_56_68 bit_56_68 bitb_56_68 word56_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_68 q_57_68 qb_57_68 bit_57_68 bitb_57_68 word57_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_68 q_58_68 qb_58_68 bit_58_68 bitb_58_68 word58_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_68 q_59_68 qb_59_68 bit_59_68 bitb_59_68 word59_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_68 q_60_68 qb_60_68 bit_60_68 bitb_60_68 word60_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_68 q_61_68 qb_61_68 bit_61_68 bitb_61_68 word61_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_68 q_62_68 qb_62_68 bit_62_68 bitb_62_68 word62_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_68 q_63_68 qb_63_68 bit_63_68 bitb_63_68 word63_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_68 q_64_68 qb_64_68 bit_64_68 bitb_64_68 word64_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_68 q_65_68 qb_65_68 bit_65_68 bitb_65_68 word65_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_68 q_66_68 qb_66_68 bit_66_68 bitb_66_68 word66_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_68 q_67_68 qb_67_68 bit_67_68 bitb_67_68 word67_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_68 q_68_68 qb_68_68 bit_68_68 bitb_68_68 word68_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_68 q_69_68 qb_69_68 bit_69_68 bitb_69_68 word69_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_68 q_70_68 qb_70_68 bit_70_68 bitb_70_68 word70_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_68 q_71_68 qb_71_68 bit_71_68 bitb_71_68 word71_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_68 q_72_68 qb_72_68 bit_72_68 bitb_72_68 word72_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_68 q_73_68 qb_73_68 bit_73_68 bitb_73_68 word73_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_68 q_74_68 qb_74_68 bit_74_68 bitb_74_68 word74_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_68 q_75_68 qb_75_68 bit_75_68 bitb_75_68 word75_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_68 q_76_68 qb_76_68 bit_76_68 bitb_76_68 word76_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_68 q_77_68 qb_77_68 bit_77_68 bitb_77_68 word77_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_68 q_78_68 qb_78_68 bit_78_68 bitb_78_68 word78_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_68 q_79_68 qb_79_68 bit_79_68 bitb_79_68 word79_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_68 q_80_68 qb_80_68 bit_80_68 bitb_80_68 word80_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_68 q_81_68 qb_81_68 bit_81_68 bitb_81_68 word81_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_68 q_82_68 qb_82_68 bit_82_68 bitb_82_68 word82_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_68 q_83_68 qb_83_68 bit_83_68 bitb_83_68 word83_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_68 q_84_68 qb_84_68 bit_84_68 bitb_84_68 word84_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_68 q_85_68 qb_85_68 bit_85_68 bitb_85_68 word85_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_68 q_86_68 qb_86_68 bit_86_68 bitb_86_68 word86_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_68 q_87_68 qb_87_68 bit_87_68 bitb_87_68 word87_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_68 q_88_68 qb_88_68 bit_88_68 bitb_88_68 word88_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_68 q_89_68 qb_89_68 bit_89_68 bitb_89_68 word89_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_68 q_90_68 qb_90_68 bit_90_68 bitb_90_68 word90_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_68 q_91_68 qb_91_68 bit_91_68 bitb_91_68 word91_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_68 q_92_68 qb_92_68 bit_92_68 bitb_92_68 word92_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_68 q_93_68 qb_93_68 bit_93_68 bitb_93_68 word93_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_68 q_94_68 qb_94_68 bit_94_68 bitb_94_68 word94_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_68 q_95_68 qb_95_68 bit_95_68 bitb_95_68 word95_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_68 q_96_68 qb_96_68 bit_96_68 bitb_96_68 word96_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_68 q_97_68 qb_97_68 bit_97_68 bitb_97_68 word97_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_68 q_98_68 qb_98_68 bit_98_68 bitb_98_68 word98_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_68 q_99_68 qb_99_68 bit_99_68 bitb_99_68 word99_68 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_69 q_0_69 qb_0_69 bit_0_69 bitb_0_69 word0_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_69 q_1_69 qb_1_69 bit_1_69 bitb_1_69 word1_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_69 q_2_69 qb_2_69 bit_2_69 bitb_2_69 word2_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_69 q_3_69 qb_3_69 bit_3_69 bitb_3_69 word3_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_69 q_4_69 qb_4_69 bit_4_69 bitb_4_69 word4_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_69 q_5_69 qb_5_69 bit_5_69 bitb_5_69 word5_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_69 q_6_69 qb_6_69 bit_6_69 bitb_6_69 word6_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_69 q_7_69 qb_7_69 bit_7_69 bitb_7_69 word7_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_69 q_8_69 qb_8_69 bit_8_69 bitb_8_69 word8_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_69 q_9_69 qb_9_69 bit_9_69 bitb_9_69 word9_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_69 q_10_69 qb_10_69 bit_10_69 bitb_10_69 word10_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_69 q_11_69 qb_11_69 bit_11_69 bitb_11_69 word11_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_69 q_12_69 qb_12_69 bit_12_69 bitb_12_69 word12_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_69 q_13_69 qb_13_69 bit_13_69 bitb_13_69 word13_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_69 q_14_69 qb_14_69 bit_14_69 bitb_14_69 word14_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_69 q_15_69 qb_15_69 bit_15_69 bitb_15_69 word15_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_69 q_16_69 qb_16_69 bit_16_69 bitb_16_69 word16_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_69 q_17_69 qb_17_69 bit_17_69 bitb_17_69 word17_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_69 q_18_69 qb_18_69 bit_18_69 bitb_18_69 word18_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_69 q_19_69 qb_19_69 bit_19_69 bitb_19_69 word19_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_69 q_20_69 qb_20_69 bit_20_69 bitb_20_69 word20_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_69 q_21_69 qb_21_69 bit_21_69 bitb_21_69 word21_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_69 q_22_69 qb_22_69 bit_22_69 bitb_22_69 word22_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_69 q_23_69 qb_23_69 bit_23_69 bitb_23_69 word23_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_69 q_24_69 qb_24_69 bit_24_69 bitb_24_69 word24_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_69 q_25_69 qb_25_69 bit_25_69 bitb_25_69 word25_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_69 q_26_69 qb_26_69 bit_26_69 bitb_26_69 word26_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_69 q_27_69 qb_27_69 bit_27_69 bitb_27_69 word27_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_69 q_28_69 qb_28_69 bit_28_69 bitb_28_69 word28_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_69 q_29_69 qb_29_69 bit_29_69 bitb_29_69 word29_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_69 q_30_69 qb_30_69 bit_30_69 bitb_30_69 word30_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_69 q_31_69 qb_31_69 bit_31_69 bitb_31_69 word31_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_69 q_32_69 qb_32_69 bit_32_69 bitb_32_69 word32_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_69 q_33_69 qb_33_69 bit_33_69 bitb_33_69 word33_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_69 q_34_69 qb_34_69 bit_34_69 bitb_34_69 word34_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_69 q_35_69 qb_35_69 bit_35_69 bitb_35_69 word35_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_69 q_36_69 qb_36_69 bit_36_69 bitb_36_69 word36_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_69 q_37_69 qb_37_69 bit_37_69 bitb_37_69 word37_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_69 q_38_69 qb_38_69 bit_38_69 bitb_38_69 word38_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_69 q_39_69 qb_39_69 bit_39_69 bitb_39_69 word39_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_69 q_40_69 qb_40_69 bit_40_69 bitb_40_69 word40_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_69 q_41_69 qb_41_69 bit_41_69 bitb_41_69 word41_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_69 q_42_69 qb_42_69 bit_42_69 bitb_42_69 word42_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_69 q_43_69 qb_43_69 bit_43_69 bitb_43_69 word43_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_69 q_44_69 qb_44_69 bit_44_69 bitb_44_69 word44_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_69 q_45_69 qb_45_69 bit_45_69 bitb_45_69 word45_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_69 q_46_69 qb_46_69 bit_46_69 bitb_46_69 word46_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_69 q_47_69 qb_47_69 bit_47_69 bitb_47_69 word47_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_69 q_48_69 qb_48_69 bit_48_69 bitb_48_69 word48_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_69 q_49_69 qb_49_69 bit_49_69 bitb_49_69 word49_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_69 q_50_69 qb_50_69 bit_50_69 bitb_50_69 word50_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_69 q_51_69 qb_51_69 bit_51_69 bitb_51_69 word51_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_69 q_52_69 qb_52_69 bit_52_69 bitb_52_69 word52_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_69 q_53_69 qb_53_69 bit_53_69 bitb_53_69 word53_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_69 q_54_69 qb_54_69 bit_54_69 bitb_54_69 word54_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_69 q_55_69 qb_55_69 bit_55_69 bitb_55_69 word55_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_69 q_56_69 qb_56_69 bit_56_69 bitb_56_69 word56_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_69 q_57_69 qb_57_69 bit_57_69 bitb_57_69 word57_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_69 q_58_69 qb_58_69 bit_58_69 bitb_58_69 word58_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_69 q_59_69 qb_59_69 bit_59_69 bitb_59_69 word59_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_69 q_60_69 qb_60_69 bit_60_69 bitb_60_69 word60_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_69 q_61_69 qb_61_69 bit_61_69 bitb_61_69 word61_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_69 q_62_69 qb_62_69 bit_62_69 bitb_62_69 word62_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_69 q_63_69 qb_63_69 bit_63_69 bitb_63_69 word63_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_69 q_64_69 qb_64_69 bit_64_69 bitb_64_69 word64_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_69 q_65_69 qb_65_69 bit_65_69 bitb_65_69 word65_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_69 q_66_69 qb_66_69 bit_66_69 bitb_66_69 word66_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_69 q_67_69 qb_67_69 bit_67_69 bitb_67_69 word67_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_69 q_68_69 qb_68_69 bit_68_69 bitb_68_69 word68_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_69 q_69_69 qb_69_69 bit_69_69 bitb_69_69 word69_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_69 q_70_69 qb_70_69 bit_70_69 bitb_70_69 word70_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_69 q_71_69 qb_71_69 bit_71_69 bitb_71_69 word71_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_69 q_72_69 qb_72_69 bit_72_69 bitb_72_69 word72_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_69 q_73_69 qb_73_69 bit_73_69 bitb_73_69 word73_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_69 q_74_69 qb_74_69 bit_74_69 bitb_74_69 word74_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_69 q_75_69 qb_75_69 bit_75_69 bitb_75_69 word75_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_69 q_76_69 qb_76_69 bit_76_69 bitb_76_69 word76_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_69 q_77_69 qb_77_69 bit_77_69 bitb_77_69 word77_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_69 q_78_69 qb_78_69 bit_78_69 bitb_78_69 word78_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_69 q_79_69 qb_79_69 bit_79_69 bitb_79_69 word79_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_69 q_80_69 qb_80_69 bit_80_69 bitb_80_69 word80_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_69 q_81_69 qb_81_69 bit_81_69 bitb_81_69 word81_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_69 q_82_69 qb_82_69 bit_82_69 bitb_82_69 word82_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_69 q_83_69 qb_83_69 bit_83_69 bitb_83_69 word83_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_69 q_84_69 qb_84_69 bit_84_69 bitb_84_69 word84_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_69 q_85_69 qb_85_69 bit_85_69 bitb_85_69 word85_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_69 q_86_69 qb_86_69 bit_86_69 bitb_86_69 word86_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_69 q_87_69 qb_87_69 bit_87_69 bitb_87_69 word87_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_69 q_88_69 qb_88_69 bit_88_69 bitb_88_69 word88_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_69 q_89_69 qb_89_69 bit_89_69 bitb_89_69 word89_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_69 q_90_69 qb_90_69 bit_90_69 bitb_90_69 word90_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_69 q_91_69 qb_91_69 bit_91_69 bitb_91_69 word91_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_69 q_92_69 qb_92_69 bit_92_69 bitb_92_69 word92_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_69 q_93_69 qb_93_69 bit_93_69 bitb_93_69 word93_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_69 q_94_69 qb_94_69 bit_94_69 bitb_94_69 word94_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_69 q_95_69 qb_95_69 bit_95_69 bitb_95_69 word95_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_69 q_96_69 qb_96_69 bit_96_69 bitb_96_69 word96_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_69 q_97_69 qb_97_69 bit_97_69 bitb_97_69 word97_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_69 q_98_69 qb_98_69 bit_98_69 bitb_98_69 word98_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_69 q_99_69 qb_99_69 bit_99_69 bitb_99_69 word99_69 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_70 q_0_70 qb_0_70 bit_0_70 bitb_0_70 word0_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_70 q_1_70 qb_1_70 bit_1_70 bitb_1_70 word1_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_70 q_2_70 qb_2_70 bit_2_70 bitb_2_70 word2_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_70 q_3_70 qb_3_70 bit_3_70 bitb_3_70 word3_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_70 q_4_70 qb_4_70 bit_4_70 bitb_4_70 word4_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_70 q_5_70 qb_5_70 bit_5_70 bitb_5_70 word5_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_70 q_6_70 qb_6_70 bit_6_70 bitb_6_70 word6_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_70 q_7_70 qb_7_70 bit_7_70 bitb_7_70 word7_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_70 q_8_70 qb_8_70 bit_8_70 bitb_8_70 word8_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_70 q_9_70 qb_9_70 bit_9_70 bitb_9_70 word9_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_70 q_10_70 qb_10_70 bit_10_70 bitb_10_70 word10_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_70 q_11_70 qb_11_70 bit_11_70 bitb_11_70 word11_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_70 q_12_70 qb_12_70 bit_12_70 bitb_12_70 word12_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_70 q_13_70 qb_13_70 bit_13_70 bitb_13_70 word13_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_70 q_14_70 qb_14_70 bit_14_70 bitb_14_70 word14_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_70 q_15_70 qb_15_70 bit_15_70 bitb_15_70 word15_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_70 q_16_70 qb_16_70 bit_16_70 bitb_16_70 word16_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_70 q_17_70 qb_17_70 bit_17_70 bitb_17_70 word17_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_70 q_18_70 qb_18_70 bit_18_70 bitb_18_70 word18_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_70 q_19_70 qb_19_70 bit_19_70 bitb_19_70 word19_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_70 q_20_70 qb_20_70 bit_20_70 bitb_20_70 word20_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_70 q_21_70 qb_21_70 bit_21_70 bitb_21_70 word21_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_70 q_22_70 qb_22_70 bit_22_70 bitb_22_70 word22_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_70 q_23_70 qb_23_70 bit_23_70 bitb_23_70 word23_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_70 q_24_70 qb_24_70 bit_24_70 bitb_24_70 word24_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_70 q_25_70 qb_25_70 bit_25_70 bitb_25_70 word25_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_70 q_26_70 qb_26_70 bit_26_70 bitb_26_70 word26_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_70 q_27_70 qb_27_70 bit_27_70 bitb_27_70 word27_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_70 q_28_70 qb_28_70 bit_28_70 bitb_28_70 word28_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_70 q_29_70 qb_29_70 bit_29_70 bitb_29_70 word29_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_70 q_30_70 qb_30_70 bit_30_70 bitb_30_70 word30_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_70 q_31_70 qb_31_70 bit_31_70 bitb_31_70 word31_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_70 q_32_70 qb_32_70 bit_32_70 bitb_32_70 word32_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_70 q_33_70 qb_33_70 bit_33_70 bitb_33_70 word33_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_70 q_34_70 qb_34_70 bit_34_70 bitb_34_70 word34_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_70 q_35_70 qb_35_70 bit_35_70 bitb_35_70 word35_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_70 q_36_70 qb_36_70 bit_36_70 bitb_36_70 word36_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_70 q_37_70 qb_37_70 bit_37_70 bitb_37_70 word37_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_70 q_38_70 qb_38_70 bit_38_70 bitb_38_70 word38_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_70 q_39_70 qb_39_70 bit_39_70 bitb_39_70 word39_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_70 q_40_70 qb_40_70 bit_40_70 bitb_40_70 word40_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_70 q_41_70 qb_41_70 bit_41_70 bitb_41_70 word41_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_70 q_42_70 qb_42_70 bit_42_70 bitb_42_70 word42_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_70 q_43_70 qb_43_70 bit_43_70 bitb_43_70 word43_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_70 q_44_70 qb_44_70 bit_44_70 bitb_44_70 word44_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_70 q_45_70 qb_45_70 bit_45_70 bitb_45_70 word45_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_70 q_46_70 qb_46_70 bit_46_70 bitb_46_70 word46_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_70 q_47_70 qb_47_70 bit_47_70 bitb_47_70 word47_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_70 q_48_70 qb_48_70 bit_48_70 bitb_48_70 word48_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_70 q_49_70 qb_49_70 bit_49_70 bitb_49_70 word49_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_70 q_50_70 qb_50_70 bit_50_70 bitb_50_70 word50_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_70 q_51_70 qb_51_70 bit_51_70 bitb_51_70 word51_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_70 q_52_70 qb_52_70 bit_52_70 bitb_52_70 word52_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_70 q_53_70 qb_53_70 bit_53_70 bitb_53_70 word53_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_70 q_54_70 qb_54_70 bit_54_70 bitb_54_70 word54_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_70 q_55_70 qb_55_70 bit_55_70 bitb_55_70 word55_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_70 q_56_70 qb_56_70 bit_56_70 bitb_56_70 word56_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_70 q_57_70 qb_57_70 bit_57_70 bitb_57_70 word57_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_70 q_58_70 qb_58_70 bit_58_70 bitb_58_70 word58_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_70 q_59_70 qb_59_70 bit_59_70 bitb_59_70 word59_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_70 q_60_70 qb_60_70 bit_60_70 bitb_60_70 word60_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_70 q_61_70 qb_61_70 bit_61_70 bitb_61_70 word61_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_70 q_62_70 qb_62_70 bit_62_70 bitb_62_70 word62_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_70 q_63_70 qb_63_70 bit_63_70 bitb_63_70 word63_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_70 q_64_70 qb_64_70 bit_64_70 bitb_64_70 word64_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_70 q_65_70 qb_65_70 bit_65_70 bitb_65_70 word65_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_70 q_66_70 qb_66_70 bit_66_70 bitb_66_70 word66_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_70 q_67_70 qb_67_70 bit_67_70 bitb_67_70 word67_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_70 q_68_70 qb_68_70 bit_68_70 bitb_68_70 word68_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_70 q_69_70 qb_69_70 bit_69_70 bitb_69_70 word69_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_70 q_70_70 qb_70_70 bit_70_70 bitb_70_70 word70_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_70 q_71_70 qb_71_70 bit_71_70 bitb_71_70 word71_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_70 q_72_70 qb_72_70 bit_72_70 bitb_72_70 word72_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_70 q_73_70 qb_73_70 bit_73_70 bitb_73_70 word73_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_70 q_74_70 qb_74_70 bit_74_70 bitb_74_70 word74_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_70 q_75_70 qb_75_70 bit_75_70 bitb_75_70 word75_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_70 q_76_70 qb_76_70 bit_76_70 bitb_76_70 word76_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_70 q_77_70 qb_77_70 bit_77_70 bitb_77_70 word77_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_70 q_78_70 qb_78_70 bit_78_70 bitb_78_70 word78_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_70 q_79_70 qb_79_70 bit_79_70 bitb_79_70 word79_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_70 q_80_70 qb_80_70 bit_80_70 bitb_80_70 word80_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_70 q_81_70 qb_81_70 bit_81_70 bitb_81_70 word81_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_70 q_82_70 qb_82_70 bit_82_70 bitb_82_70 word82_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_70 q_83_70 qb_83_70 bit_83_70 bitb_83_70 word83_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_70 q_84_70 qb_84_70 bit_84_70 bitb_84_70 word84_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_70 q_85_70 qb_85_70 bit_85_70 bitb_85_70 word85_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_70 q_86_70 qb_86_70 bit_86_70 bitb_86_70 word86_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_70 q_87_70 qb_87_70 bit_87_70 bitb_87_70 word87_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_70 q_88_70 qb_88_70 bit_88_70 bitb_88_70 word88_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_70 q_89_70 qb_89_70 bit_89_70 bitb_89_70 word89_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_70 q_90_70 qb_90_70 bit_90_70 bitb_90_70 word90_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_70 q_91_70 qb_91_70 bit_91_70 bitb_91_70 word91_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_70 q_92_70 qb_92_70 bit_92_70 bitb_92_70 word92_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_70 q_93_70 qb_93_70 bit_93_70 bitb_93_70 word93_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_70 q_94_70 qb_94_70 bit_94_70 bitb_94_70 word94_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_70 q_95_70 qb_95_70 bit_95_70 bitb_95_70 word95_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_70 q_96_70 qb_96_70 bit_96_70 bitb_96_70 word96_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_70 q_97_70 qb_97_70 bit_97_70 bitb_97_70 word97_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_70 q_98_70 qb_98_70 bit_98_70 bitb_98_70 word98_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_70 q_99_70 qb_99_70 bit_99_70 bitb_99_70 word99_70 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_71 q_0_71 qb_0_71 bit_0_71 bitb_0_71 word0_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_71 q_1_71 qb_1_71 bit_1_71 bitb_1_71 word1_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_71 q_2_71 qb_2_71 bit_2_71 bitb_2_71 word2_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_71 q_3_71 qb_3_71 bit_3_71 bitb_3_71 word3_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_71 q_4_71 qb_4_71 bit_4_71 bitb_4_71 word4_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_71 q_5_71 qb_5_71 bit_5_71 bitb_5_71 word5_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_71 q_6_71 qb_6_71 bit_6_71 bitb_6_71 word6_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_71 q_7_71 qb_7_71 bit_7_71 bitb_7_71 word7_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_71 q_8_71 qb_8_71 bit_8_71 bitb_8_71 word8_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_71 q_9_71 qb_9_71 bit_9_71 bitb_9_71 word9_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_71 q_10_71 qb_10_71 bit_10_71 bitb_10_71 word10_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_71 q_11_71 qb_11_71 bit_11_71 bitb_11_71 word11_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_71 q_12_71 qb_12_71 bit_12_71 bitb_12_71 word12_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_71 q_13_71 qb_13_71 bit_13_71 bitb_13_71 word13_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_71 q_14_71 qb_14_71 bit_14_71 bitb_14_71 word14_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_71 q_15_71 qb_15_71 bit_15_71 bitb_15_71 word15_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_71 q_16_71 qb_16_71 bit_16_71 bitb_16_71 word16_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_71 q_17_71 qb_17_71 bit_17_71 bitb_17_71 word17_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_71 q_18_71 qb_18_71 bit_18_71 bitb_18_71 word18_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_71 q_19_71 qb_19_71 bit_19_71 bitb_19_71 word19_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_71 q_20_71 qb_20_71 bit_20_71 bitb_20_71 word20_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_71 q_21_71 qb_21_71 bit_21_71 bitb_21_71 word21_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_71 q_22_71 qb_22_71 bit_22_71 bitb_22_71 word22_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_71 q_23_71 qb_23_71 bit_23_71 bitb_23_71 word23_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_71 q_24_71 qb_24_71 bit_24_71 bitb_24_71 word24_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_71 q_25_71 qb_25_71 bit_25_71 bitb_25_71 word25_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_71 q_26_71 qb_26_71 bit_26_71 bitb_26_71 word26_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_71 q_27_71 qb_27_71 bit_27_71 bitb_27_71 word27_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_71 q_28_71 qb_28_71 bit_28_71 bitb_28_71 word28_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_71 q_29_71 qb_29_71 bit_29_71 bitb_29_71 word29_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_71 q_30_71 qb_30_71 bit_30_71 bitb_30_71 word30_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_71 q_31_71 qb_31_71 bit_31_71 bitb_31_71 word31_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_71 q_32_71 qb_32_71 bit_32_71 bitb_32_71 word32_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_71 q_33_71 qb_33_71 bit_33_71 bitb_33_71 word33_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_71 q_34_71 qb_34_71 bit_34_71 bitb_34_71 word34_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_71 q_35_71 qb_35_71 bit_35_71 bitb_35_71 word35_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_71 q_36_71 qb_36_71 bit_36_71 bitb_36_71 word36_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_71 q_37_71 qb_37_71 bit_37_71 bitb_37_71 word37_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_71 q_38_71 qb_38_71 bit_38_71 bitb_38_71 word38_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_71 q_39_71 qb_39_71 bit_39_71 bitb_39_71 word39_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_71 q_40_71 qb_40_71 bit_40_71 bitb_40_71 word40_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_71 q_41_71 qb_41_71 bit_41_71 bitb_41_71 word41_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_71 q_42_71 qb_42_71 bit_42_71 bitb_42_71 word42_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_71 q_43_71 qb_43_71 bit_43_71 bitb_43_71 word43_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_71 q_44_71 qb_44_71 bit_44_71 bitb_44_71 word44_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_71 q_45_71 qb_45_71 bit_45_71 bitb_45_71 word45_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_71 q_46_71 qb_46_71 bit_46_71 bitb_46_71 word46_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_71 q_47_71 qb_47_71 bit_47_71 bitb_47_71 word47_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_71 q_48_71 qb_48_71 bit_48_71 bitb_48_71 word48_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_71 q_49_71 qb_49_71 bit_49_71 bitb_49_71 word49_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_71 q_50_71 qb_50_71 bit_50_71 bitb_50_71 word50_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_71 q_51_71 qb_51_71 bit_51_71 bitb_51_71 word51_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_71 q_52_71 qb_52_71 bit_52_71 bitb_52_71 word52_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_71 q_53_71 qb_53_71 bit_53_71 bitb_53_71 word53_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_71 q_54_71 qb_54_71 bit_54_71 bitb_54_71 word54_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_71 q_55_71 qb_55_71 bit_55_71 bitb_55_71 word55_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_71 q_56_71 qb_56_71 bit_56_71 bitb_56_71 word56_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_71 q_57_71 qb_57_71 bit_57_71 bitb_57_71 word57_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_71 q_58_71 qb_58_71 bit_58_71 bitb_58_71 word58_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_71 q_59_71 qb_59_71 bit_59_71 bitb_59_71 word59_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_71 q_60_71 qb_60_71 bit_60_71 bitb_60_71 word60_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_71 q_61_71 qb_61_71 bit_61_71 bitb_61_71 word61_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_71 q_62_71 qb_62_71 bit_62_71 bitb_62_71 word62_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_71 q_63_71 qb_63_71 bit_63_71 bitb_63_71 word63_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_71 q_64_71 qb_64_71 bit_64_71 bitb_64_71 word64_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_71 q_65_71 qb_65_71 bit_65_71 bitb_65_71 word65_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_71 q_66_71 qb_66_71 bit_66_71 bitb_66_71 word66_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_71 q_67_71 qb_67_71 bit_67_71 bitb_67_71 word67_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_71 q_68_71 qb_68_71 bit_68_71 bitb_68_71 word68_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_71 q_69_71 qb_69_71 bit_69_71 bitb_69_71 word69_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_71 q_70_71 qb_70_71 bit_70_71 bitb_70_71 word70_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_71 q_71_71 qb_71_71 bit_71_71 bitb_71_71 word71_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_71 q_72_71 qb_72_71 bit_72_71 bitb_72_71 word72_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_71 q_73_71 qb_73_71 bit_73_71 bitb_73_71 word73_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_71 q_74_71 qb_74_71 bit_74_71 bitb_74_71 word74_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_71 q_75_71 qb_75_71 bit_75_71 bitb_75_71 word75_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_71 q_76_71 qb_76_71 bit_76_71 bitb_76_71 word76_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_71 q_77_71 qb_77_71 bit_77_71 bitb_77_71 word77_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_71 q_78_71 qb_78_71 bit_78_71 bitb_78_71 word78_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_71 q_79_71 qb_79_71 bit_79_71 bitb_79_71 word79_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_71 q_80_71 qb_80_71 bit_80_71 bitb_80_71 word80_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_71 q_81_71 qb_81_71 bit_81_71 bitb_81_71 word81_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_71 q_82_71 qb_82_71 bit_82_71 bitb_82_71 word82_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_71 q_83_71 qb_83_71 bit_83_71 bitb_83_71 word83_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_71 q_84_71 qb_84_71 bit_84_71 bitb_84_71 word84_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_71 q_85_71 qb_85_71 bit_85_71 bitb_85_71 word85_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_71 q_86_71 qb_86_71 bit_86_71 bitb_86_71 word86_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_71 q_87_71 qb_87_71 bit_87_71 bitb_87_71 word87_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_71 q_88_71 qb_88_71 bit_88_71 bitb_88_71 word88_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_71 q_89_71 qb_89_71 bit_89_71 bitb_89_71 word89_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_71 q_90_71 qb_90_71 bit_90_71 bitb_90_71 word90_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_71 q_91_71 qb_91_71 bit_91_71 bitb_91_71 word91_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_71 q_92_71 qb_92_71 bit_92_71 bitb_92_71 word92_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_71 q_93_71 qb_93_71 bit_93_71 bitb_93_71 word93_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_71 q_94_71 qb_94_71 bit_94_71 bitb_94_71 word94_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_71 q_95_71 qb_95_71 bit_95_71 bitb_95_71 word95_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_71 q_96_71 qb_96_71 bit_96_71 bitb_96_71 word96_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_71 q_97_71 qb_97_71 bit_97_71 bitb_97_71 word97_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_71 q_98_71 qb_98_71 bit_98_71 bitb_98_71 word98_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_71 q_99_71 qb_99_71 bit_99_71 bitb_99_71 word99_71 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_72 q_0_72 qb_0_72 bit_0_72 bitb_0_72 word0_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_72 q_1_72 qb_1_72 bit_1_72 bitb_1_72 word1_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_72 q_2_72 qb_2_72 bit_2_72 bitb_2_72 word2_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_72 q_3_72 qb_3_72 bit_3_72 bitb_3_72 word3_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_72 q_4_72 qb_4_72 bit_4_72 bitb_4_72 word4_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_72 q_5_72 qb_5_72 bit_5_72 bitb_5_72 word5_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_72 q_6_72 qb_6_72 bit_6_72 bitb_6_72 word6_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_72 q_7_72 qb_7_72 bit_7_72 bitb_7_72 word7_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_72 q_8_72 qb_8_72 bit_8_72 bitb_8_72 word8_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_72 q_9_72 qb_9_72 bit_9_72 bitb_9_72 word9_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_72 q_10_72 qb_10_72 bit_10_72 bitb_10_72 word10_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_72 q_11_72 qb_11_72 bit_11_72 bitb_11_72 word11_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_72 q_12_72 qb_12_72 bit_12_72 bitb_12_72 word12_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_72 q_13_72 qb_13_72 bit_13_72 bitb_13_72 word13_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_72 q_14_72 qb_14_72 bit_14_72 bitb_14_72 word14_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_72 q_15_72 qb_15_72 bit_15_72 bitb_15_72 word15_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_72 q_16_72 qb_16_72 bit_16_72 bitb_16_72 word16_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_72 q_17_72 qb_17_72 bit_17_72 bitb_17_72 word17_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_72 q_18_72 qb_18_72 bit_18_72 bitb_18_72 word18_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_72 q_19_72 qb_19_72 bit_19_72 bitb_19_72 word19_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_72 q_20_72 qb_20_72 bit_20_72 bitb_20_72 word20_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_72 q_21_72 qb_21_72 bit_21_72 bitb_21_72 word21_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_72 q_22_72 qb_22_72 bit_22_72 bitb_22_72 word22_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_72 q_23_72 qb_23_72 bit_23_72 bitb_23_72 word23_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_72 q_24_72 qb_24_72 bit_24_72 bitb_24_72 word24_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_72 q_25_72 qb_25_72 bit_25_72 bitb_25_72 word25_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_72 q_26_72 qb_26_72 bit_26_72 bitb_26_72 word26_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_72 q_27_72 qb_27_72 bit_27_72 bitb_27_72 word27_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_72 q_28_72 qb_28_72 bit_28_72 bitb_28_72 word28_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_72 q_29_72 qb_29_72 bit_29_72 bitb_29_72 word29_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_72 q_30_72 qb_30_72 bit_30_72 bitb_30_72 word30_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_72 q_31_72 qb_31_72 bit_31_72 bitb_31_72 word31_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_72 q_32_72 qb_32_72 bit_32_72 bitb_32_72 word32_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_72 q_33_72 qb_33_72 bit_33_72 bitb_33_72 word33_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_72 q_34_72 qb_34_72 bit_34_72 bitb_34_72 word34_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_72 q_35_72 qb_35_72 bit_35_72 bitb_35_72 word35_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_72 q_36_72 qb_36_72 bit_36_72 bitb_36_72 word36_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_72 q_37_72 qb_37_72 bit_37_72 bitb_37_72 word37_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_72 q_38_72 qb_38_72 bit_38_72 bitb_38_72 word38_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_72 q_39_72 qb_39_72 bit_39_72 bitb_39_72 word39_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_72 q_40_72 qb_40_72 bit_40_72 bitb_40_72 word40_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_72 q_41_72 qb_41_72 bit_41_72 bitb_41_72 word41_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_72 q_42_72 qb_42_72 bit_42_72 bitb_42_72 word42_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_72 q_43_72 qb_43_72 bit_43_72 bitb_43_72 word43_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_72 q_44_72 qb_44_72 bit_44_72 bitb_44_72 word44_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_72 q_45_72 qb_45_72 bit_45_72 bitb_45_72 word45_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_72 q_46_72 qb_46_72 bit_46_72 bitb_46_72 word46_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_72 q_47_72 qb_47_72 bit_47_72 bitb_47_72 word47_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_72 q_48_72 qb_48_72 bit_48_72 bitb_48_72 word48_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_72 q_49_72 qb_49_72 bit_49_72 bitb_49_72 word49_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_72 q_50_72 qb_50_72 bit_50_72 bitb_50_72 word50_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_72 q_51_72 qb_51_72 bit_51_72 bitb_51_72 word51_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_72 q_52_72 qb_52_72 bit_52_72 bitb_52_72 word52_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_72 q_53_72 qb_53_72 bit_53_72 bitb_53_72 word53_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_72 q_54_72 qb_54_72 bit_54_72 bitb_54_72 word54_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_72 q_55_72 qb_55_72 bit_55_72 bitb_55_72 word55_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_72 q_56_72 qb_56_72 bit_56_72 bitb_56_72 word56_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_72 q_57_72 qb_57_72 bit_57_72 bitb_57_72 word57_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_72 q_58_72 qb_58_72 bit_58_72 bitb_58_72 word58_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_72 q_59_72 qb_59_72 bit_59_72 bitb_59_72 word59_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_72 q_60_72 qb_60_72 bit_60_72 bitb_60_72 word60_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_72 q_61_72 qb_61_72 bit_61_72 bitb_61_72 word61_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_72 q_62_72 qb_62_72 bit_62_72 bitb_62_72 word62_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_72 q_63_72 qb_63_72 bit_63_72 bitb_63_72 word63_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_72 q_64_72 qb_64_72 bit_64_72 bitb_64_72 word64_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_72 q_65_72 qb_65_72 bit_65_72 bitb_65_72 word65_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_72 q_66_72 qb_66_72 bit_66_72 bitb_66_72 word66_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_72 q_67_72 qb_67_72 bit_67_72 bitb_67_72 word67_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_72 q_68_72 qb_68_72 bit_68_72 bitb_68_72 word68_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_72 q_69_72 qb_69_72 bit_69_72 bitb_69_72 word69_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_72 q_70_72 qb_70_72 bit_70_72 bitb_70_72 word70_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_72 q_71_72 qb_71_72 bit_71_72 bitb_71_72 word71_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_72 q_72_72 qb_72_72 bit_72_72 bitb_72_72 word72_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_72 q_73_72 qb_73_72 bit_73_72 bitb_73_72 word73_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_72 q_74_72 qb_74_72 bit_74_72 bitb_74_72 word74_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_72 q_75_72 qb_75_72 bit_75_72 bitb_75_72 word75_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_72 q_76_72 qb_76_72 bit_76_72 bitb_76_72 word76_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_72 q_77_72 qb_77_72 bit_77_72 bitb_77_72 word77_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_72 q_78_72 qb_78_72 bit_78_72 bitb_78_72 word78_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_72 q_79_72 qb_79_72 bit_79_72 bitb_79_72 word79_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_72 q_80_72 qb_80_72 bit_80_72 bitb_80_72 word80_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_72 q_81_72 qb_81_72 bit_81_72 bitb_81_72 word81_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_72 q_82_72 qb_82_72 bit_82_72 bitb_82_72 word82_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_72 q_83_72 qb_83_72 bit_83_72 bitb_83_72 word83_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_72 q_84_72 qb_84_72 bit_84_72 bitb_84_72 word84_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_72 q_85_72 qb_85_72 bit_85_72 bitb_85_72 word85_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_72 q_86_72 qb_86_72 bit_86_72 bitb_86_72 word86_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_72 q_87_72 qb_87_72 bit_87_72 bitb_87_72 word87_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_72 q_88_72 qb_88_72 bit_88_72 bitb_88_72 word88_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_72 q_89_72 qb_89_72 bit_89_72 bitb_89_72 word89_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_72 q_90_72 qb_90_72 bit_90_72 bitb_90_72 word90_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_72 q_91_72 qb_91_72 bit_91_72 bitb_91_72 word91_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_72 q_92_72 qb_92_72 bit_92_72 bitb_92_72 word92_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_72 q_93_72 qb_93_72 bit_93_72 bitb_93_72 word93_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_72 q_94_72 qb_94_72 bit_94_72 bitb_94_72 word94_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_72 q_95_72 qb_95_72 bit_95_72 bitb_95_72 word95_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_72 q_96_72 qb_96_72 bit_96_72 bitb_96_72 word96_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_72 q_97_72 qb_97_72 bit_97_72 bitb_97_72 word97_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_72 q_98_72 qb_98_72 bit_98_72 bitb_98_72 word98_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_72 q_99_72 qb_99_72 bit_99_72 bitb_99_72 word99_72 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_73 q_0_73 qb_0_73 bit_0_73 bitb_0_73 word0_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_73 q_1_73 qb_1_73 bit_1_73 bitb_1_73 word1_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_73 q_2_73 qb_2_73 bit_2_73 bitb_2_73 word2_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_73 q_3_73 qb_3_73 bit_3_73 bitb_3_73 word3_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_73 q_4_73 qb_4_73 bit_4_73 bitb_4_73 word4_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_73 q_5_73 qb_5_73 bit_5_73 bitb_5_73 word5_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_73 q_6_73 qb_6_73 bit_6_73 bitb_6_73 word6_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_73 q_7_73 qb_7_73 bit_7_73 bitb_7_73 word7_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_73 q_8_73 qb_8_73 bit_8_73 bitb_8_73 word8_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_73 q_9_73 qb_9_73 bit_9_73 bitb_9_73 word9_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_73 q_10_73 qb_10_73 bit_10_73 bitb_10_73 word10_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_73 q_11_73 qb_11_73 bit_11_73 bitb_11_73 word11_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_73 q_12_73 qb_12_73 bit_12_73 bitb_12_73 word12_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_73 q_13_73 qb_13_73 bit_13_73 bitb_13_73 word13_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_73 q_14_73 qb_14_73 bit_14_73 bitb_14_73 word14_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_73 q_15_73 qb_15_73 bit_15_73 bitb_15_73 word15_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_73 q_16_73 qb_16_73 bit_16_73 bitb_16_73 word16_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_73 q_17_73 qb_17_73 bit_17_73 bitb_17_73 word17_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_73 q_18_73 qb_18_73 bit_18_73 bitb_18_73 word18_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_73 q_19_73 qb_19_73 bit_19_73 bitb_19_73 word19_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_73 q_20_73 qb_20_73 bit_20_73 bitb_20_73 word20_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_73 q_21_73 qb_21_73 bit_21_73 bitb_21_73 word21_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_73 q_22_73 qb_22_73 bit_22_73 bitb_22_73 word22_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_73 q_23_73 qb_23_73 bit_23_73 bitb_23_73 word23_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_73 q_24_73 qb_24_73 bit_24_73 bitb_24_73 word24_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_73 q_25_73 qb_25_73 bit_25_73 bitb_25_73 word25_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_73 q_26_73 qb_26_73 bit_26_73 bitb_26_73 word26_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_73 q_27_73 qb_27_73 bit_27_73 bitb_27_73 word27_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_73 q_28_73 qb_28_73 bit_28_73 bitb_28_73 word28_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_73 q_29_73 qb_29_73 bit_29_73 bitb_29_73 word29_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_73 q_30_73 qb_30_73 bit_30_73 bitb_30_73 word30_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_73 q_31_73 qb_31_73 bit_31_73 bitb_31_73 word31_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_73 q_32_73 qb_32_73 bit_32_73 bitb_32_73 word32_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_73 q_33_73 qb_33_73 bit_33_73 bitb_33_73 word33_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_73 q_34_73 qb_34_73 bit_34_73 bitb_34_73 word34_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_73 q_35_73 qb_35_73 bit_35_73 bitb_35_73 word35_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_73 q_36_73 qb_36_73 bit_36_73 bitb_36_73 word36_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_73 q_37_73 qb_37_73 bit_37_73 bitb_37_73 word37_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_73 q_38_73 qb_38_73 bit_38_73 bitb_38_73 word38_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_73 q_39_73 qb_39_73 bit_39_73 bitb_39_73 word39_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_73 q_40_73 qb_40_73 bit_40_73 bitb_40_73 word40_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_73 q_41_73 qb_41_73 bit_41_73 bitb_41_73 word41_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_73 q_42_73 qb_42_73 bit_42_73 bitb_42_73 word42_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_73 q_43_73 qb_43_73 bit_43_73 bitb_43_73 word43_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_73 q_44_73 qb_44_73 bit_44_73 bitb_44_73 word44_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_73 q_45_73 qb_45_73 bit_45_73 bitb_45_73 word45_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_73 q_46_73 qb_46_73 bit_46_73 bitb_46_73 word46_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_73 q_47_73 qb_47_73 bit_47_73 bitb_47_73 word47_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_73 q_48_73 qb_48_73 bit_48_73 bitb_48_73 word48_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_73 q_49_73 qb_49_73 bit_49_73 bitb_49_73 word49_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_73 q_50_73 qb_50_73 bit_50_73 bitb_50_73 word50_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_73 q_51_73 qb_51_73 bit_51_73 bitb_51_73 word51_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_73 q_52_73 qb_52_73 bit_52_73 bitb_52_73 word52_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_73 q_53_73 qb_53_73 bit_53_73 bitb_53_73 word53_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_73 q_54_73 qb_54_73 bit_54_73 bitb_54_73 word54_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_73 q_55_73 qb_55_73 bit_55_73 bitb_55_73 word55_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_73 q_56_73 qb_56_73 bit_56_73 bitb_56_73 word56_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_73 q_57_73 qb_57_73 bit_57_73 bitb_57_73 word57_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_73 q_58_73 qb_58_73 bit_58_73 bitb_58_73 word58_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_73 q_59_73 qb_59_73 bit_59_73 bitb_59_73 word59_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_73 q_60_73 qb_60_73 bit_60_73 bitb_60_73 word60_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_73 q_61_73 qb_61_73 bit_61_73 bitb_61_73 word61_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_73 q_62_73 qb_62_73 bit_62_73 bitb_62_73 word62_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_73 q_63_73 qb_63_73 bit_63_73 bitb_63_73 word63_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_73 q_64_73 qb_64_73 bit_64_73 bitb_64_73 word64_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_73 q_65_73 qb_65_73 bit_65_73 bitb_65_73 word65_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_73 q_66_73 qb_66_73 bit_66_73 bitb_66_73 word66_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_73 q_67_73 qb_67_73 bit_67_73 bitb_67_73 word67_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_73 q_68_73 qb_68_73 bit_68_73 bitb_68_73 word68_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_73 q_69_73 qb_69_73 bit_69_73 bitb_69_73 word69_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_73 q_70_73 qb_70_73 bit_70_73 bitb_70_73 word70_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_73 q_71_73 qb_71_73 bit_71_73 bitb_71_73 word71_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_73 q_72_73 qb_72_73 bit_72_73 bitb_72_73 word72_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_73 q_73_73 qb_73_73 bit_73_73 bitb_73_73 word73_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_73 q_74_73 qb_74_73 bit_74_73 bitb_74_73 word74_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_73 q_75_73 qb_75_73 bit_75_73 bitb_75_73 word75_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_73 q_76_73 qb_76_73 bit_76_73 bitb_76_73 word76_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_73 q_77_73 qb_77_73 bit_77_73 bitb_77_73 word77_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_73 q_78_73 qb_78_73 bit_78_73 bitb_78_73 word78_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_73 q_79_73 qb_79_73 bit_79_73 bitb_79_73 word79_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_73 q_80_73 qb_80_73 bit_80_73 bitb_80_73 word80_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_73 q_81_73 qb_81_73 bit_81_73 bitb_81_73 word81_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_73 q_82_73 qb_82_73 bit_82_73 bitb_82_73 word82_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_73 q_83_73 qb_83_73 bit_83_73 bitb_83_73 word83_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_73 q_84_73 qb_84_73 bit_84_73 bitb_84_73 word84_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_73 q_85_73 qb_85_73 bit_85_73 bitb_85_73 word85_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_73 q_86_73 qb_86_73 bit_86_73 bitb_86_73 word86_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_73 q_87_73 qb_87_73 bit_87_73 bitb_87_73 word87_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_73 q_88_73 qb_88_73 bit_88_73 bitb_88_73 word88_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_73 q_89_73 qb_89_73 bit_89_73 bitb_89_73 word89_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_73 q_90_73 qb_90_73 bit_90_73 bitb_90_73 word90_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_73 q_91_73 qb_91_73 bit_91_73 bitb_91_73 word91_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_73 q_92_73 qb_92_73 bit_92_73 bitb_92_73 word92_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_73 q_93_73 qb_93_73 bit_93_73 bitb_93_73 word93_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_73 q_94_73 qb_94_73 bit_94_73 bitb_94_73 word94_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_73 q_95_73 qb_95_73 bit_95_73 bitb_95_73 word95_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_73 q_96_73 qb_96_73 bit_96_73 bitb_96_73 word96_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_73 q_97_73 qb_97_73 bit_97_73 bitb_97_73 word97_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_73 q_98_73 qb_98_73 bit_98_73 bitb_98_73 word98_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_73 q_99_73 qb_99_73 bit_99_73 bitb_99_73 word99_73 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_74 q_0_74 qb_0_74 bit_0_74 bitb_0_74 word0_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_74 q_1_74 qb_1_74 bit_1_74 bitb_1_74 word1_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_74 q_2_74 qb_2_74 bit_2_74 bitb_2_74 word2_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_74 q_3_74 qb_3_74 bit_3_74 bitb_3_74 word3_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_74 q_4_74 qb_4_74 bit_4_74 bitb_4_74 word4_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_74 q_5_74 qb_5_74 bit_5_74 bitb_5_74 word5_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_74 q_6_74 qb_6_74 bit_6_74 bitb_6_74 word6_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_74 q_7_74 qb_7_74 bit_7_74 bitb_7_74 word7_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_74 q_8_74 qb_8_74 bit_8_74 bitb_8_74 word8_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_74 q_9_74 qb_9_74 bit_9_74 bitb_9_74 word9_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_74 q_10_74 qb_10_74 bit_10_74 bitb_10_74 word10_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_74 q_11_74 qb_11_74 bit_11_74 bitb_11_74 word11_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_74 q_12_74 qb_12_74 bit_12_74 bitb_12_74 word12_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_74 q_13_74 qb_13_74 bit_13_74 bitb_13_74 word13_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_74 q_14_74 qb_14_74 bit_14_74 bitb_14_74 word14_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_74 q_15_74 qb_15_74 bit_15_74 bitb_15_74 word15_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_74 q_16_74 qb_16_74 bit_16_74 bitb_16_74 word16_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_74 q_17_74 qb_17_74 bit_17_74 bitb_17_74 word17_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_74 q_18_74 qb_18_74 bit_18_74 bitb_18_74 word18_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_74 q_19_74 qb_19_74 bit_19_74 bitb_19_74 word19_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_74 q_20_74 qb_20_74 bit_20_74 bitb_20_74 word20_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_74 q_21_74 qb_21_74 bit_21_74 bitb_21_74 word21_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_74 q_22_74 qb_22_74 bit_22_74 bitb_22_74 word22_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_74 q_23_74 qb_23_74 bit_23_74 bitb_23_74 word23_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_74 q_24_74 qb_24_74 bit_24_74 bitb_24_74 word24_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_74 q_25_74 qb_25_74 bit_25_74 bitb_25_74 word25_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_74 q_26_74 qb_26_74 bit_26_74 bitb_26_74 word26_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_74 q_27_74 qb_27_74 bit_27_74 bitb_27_74 word27_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_74 q_28_74 qb_28_74 bit_28_74 bitb_28_74 word28_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_74 q_29_74 qb_29_74 bit_29_74 bitb_29_74 word29_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_74 q_30_74 qb_30_74 bit_30_74 bitb_30_74 word30_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_74 q_31_74 qb_31_74 bit_31_74 bitb_31_74 word31_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_74 q_32_74 qb_32_74 bit_32_74 bitb_32_74 word32_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_74 q_33_74 qb_33_74 bit_33_74 bitb_33_74 word33_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_74 q_34_74 qb_34_74 bit_34_74 bitb_34_74 word34_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_74 q_35_74 qb_35_74 bit_35_74 bitb_35_74 word35_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_74 q_36_74 qb_36_74 bit_36_74 bitb_36_74 word36_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_74 q_37_74 qb_37_74 bit_37_74 bitb_37_74 word37_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_74 q_38_74 qb_38_74 bit_38_74 bitb_38_74 word38_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_74 q_39_74 qb_39_74 bit_39_74 bitb_39_74 word39_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_74 q_40_74 qb_40_74 bit_40_74 bitb_40_74 word40_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_74 q_41_74 qb_41_74 bit_41_74 bitb_41_74 word41_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_74 q_42_74 qb_42_74 bit_42_74 bitb_42_74 word42_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_74 q_43_74 qb_43_74 bit_43_74 bitb_43_74 word43_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_74 q_44_74 qb_44_74 bit_44_74 bitb_44_74 word44_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_74 q_45_74 qb_45_74 bit_45_74 bitb_45_74 word45_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_74 q_46_74 qb_46_74 bit_46_74 bitb_46_74 word46_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_74 q_47_74 qb_47_74 bit_47_74 bitb_47_74 word47_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_74 q_48_74 qb_48_74 bit_48_74 bitb_48_74 word48_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_74 q_49_74 qb_49_74 bit_49_74 bitb_49_74 word49_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_74 q_50_74 qb_50_74 bit_50_74 bitb_50_74 word50_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_74 q_51_74 qb_51_74 bit_51_74 bitb_51_74 word51_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_74 q_52_74 qb_52_74 bit_52_74 bitb_52_74 word52_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_74 q_53_74 qb_53_74 bit_53_74 bitb_53_74 word53_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_74 q_54_74 qb_54_74 bit_54_74 bitb_54_74 word54_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_74 q_55_74 qb_55_74 bit_55_74 bitb_55_74 word55_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_74 q_56_74 qb_56_74 bit_56_74 bitb_56_74 word56_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_74 q_57_74 qb_57_74 bit_57_74 bitb_57_74 word57_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_74 q_58_74 qb_58_74 bit_58_74 bitb_58_74 word58_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_74 q_59_74 qb_59_74 bit_59_74 bitb_59_74 word59_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_74 q_60_74 qb_60_74 bit_60_74 bitb_60_74 word60_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_74 q_61_74 qb_61_74 bit_61_74 bitb_61_74 word61_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_74 q_62_74 qb_62_74 bit_62_74 bitb_62_74 word62_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_74 q_63_74 qb_63_74 bit_63_74 bitb_63_74 word63_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_74 q_64_74 qb_64_74 bit_64_74 bitb_64_74 word64_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_74 q_65_74 qb_65_74 bit_65_74 bitb_65_74 word65_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_74 q_66_74 qb_66_74 bit_66_74 bitb_66_74 word66_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_74 q_67_74 qb_67_74 bit_67_74 bitb_67_74 word67_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_74 q_68_74 qb_68_74 bit_68_74 bitb_68_74 word68_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_74 q_69_74 qb_69_74 bit_69_74 bitb_69_74 word69_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_74 q_70_74 qb_70_74 bit_70_74 bitb_70_74 word70_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_74 q_71_74 qb_71_74 bit_71_74 bitb_71_74 word71_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_74 q_72_74 qb_72_74 bit_72_74 bitb_72_74 word72_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_74 q_73_74 qb_73_74 bit_73_74 bitb_73_74 word73_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_74 q_74_74 qb_74_74 bit_74_74 bitb_74_74 word74_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_74 q_75_74 qb_75_74 bit_75_74 bitb_75_74 word75_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_74 q_76_74 qb_76_74 bit_76_74 bitb_76_74 word76_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_74 q_77_74 qb_77_74 bit_77_74 bitb_77_74 word77_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_74 q_78_74 qb_78_74 bit_78_74 bitb_78_74 word78_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_74 q_79_74 qb_79_74 bit_79_74 bitb_79_74 word79_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_74 q_80_74 qb_80_74 bit_80_74 bitb_80_74 word80_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_74 q_81_74 qb_81_74 bit_81_74 bitb_81_74 word81_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_74 q_82_74 qb_82_74 bit_82_74 bitb_82_74 word82_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_74 q_83_74 qb_83_74 bit_83_74 bitb_83_74 word83_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_74 q_84_74 qb_84_74 bit_84_74 bitb_84_74 word84_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_74 q_85_74 qb_85_74 bit_85_74 bitb_85_74 word85_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_74 q_86_74 qb_86_74 bit_86_74 bitb_86_74 word86_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_74 q_87_74 qb_87_74 bit_87_74 bitb_87_74 word87_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_74 q_88_74 qb_88_74 bit_88_74 bitb_88_74 word88_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_74 q_89_74 qb_89_74 bit_89_74 bitb_89_74 word89_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_74 q_90_74 qb_90_74 bit_90_74 bitb_90_74 word90_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_74 q_91_74 qb_91_74 bit_91_74 bitb_91_74 word91_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_74 q_92_74 qb_92_74 bit_92_74 bitb_92_74 word92_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_74 q_93_74 qb_93_74 bit_93_74 bitb_93_74 word93_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_74 q_94_74 qb_94_74 bit_94_74 bitb_94_74 word94_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_74 q_95_74 qb_95_74 bit_95_74 bitb_95_74 word95_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_74 q_96_74 qb_96_74 bit_96_74 bitb_96_74 word96_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_74 q_97_74 qb_97_74 bit_97_74 bitb_97_74 word97_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_74 q_98_74 qb_98_74 bit_98_74 bitb_98_74 word98_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_74 q_99_74 qb_99_74 bit_99_74 bitb_99_74 word99_74 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_75 q_0_75 qb_0_75 bit_0_75 bitb_0_75 word0_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_75 q_1_75 qb_1_75 bit_1_75 bitb_1_75 word1_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_75 q_2_75 qb_2_75 bit_2_75 bitb_2_75 word2_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_75 q_3_75 qb_3_75 bit_3_75 bitb_3_75 word3_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_75 q_4_75 qb_4_75 bit_4_75 bitb_4_75 word4_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_75 q_5_75 qb_5_75 bit_5_75 bitb_5_75 word5_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_75 q_6_75 qb_6_75 bit_6_75 bitb_6_75 word6_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_75 q_7_75 qb_7_75 bit_7_75 bitb_7_75 word7_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_75 q_8_75 qb_8_75 bit_8_75 bitb_8_75 word8_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_75 q_9_75 qb_9_75 bit_9_75 bitb_9_75 word9_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_75 q_10_75 qb_10_75 bit_10_75 bitb_10_75 word10_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_75 q_11_75 qb_11_75 bit_11_75 bitb_11_75 word11_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_75 q_12_75 qb_12_75 bit_12_75 bitb_12_75 word12_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_75 q_13_75 qb_13_75 bit_13_75 bitb_13_75 word13_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_75 q_14_75 qb_14_75 bit_14_75 bitb_14_75 word14_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_75 q_15_75 qb_15_75 bit_15_75 bitb_15_75 word15_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_75 q_16_75 qb_16_75 bit_16_75 bitb_16_75 word16_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_75 q_17_75 qb_17_75 bit_17_75 bitb_17_75 word17_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_75 q_18_75 qb_18_75 bit_18_75 bitb_18_75 word18_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_75 q_19_75 qb_19_75 bit_19_75 bitb_19_75 word19_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_75 q_20_75 qb_20_75 bit_20_75 bitb_20_75 word20_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_75 q_21_75 qb_21_75 bit_21_75 bitb_21_75 word21_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_75 q_22_75 qb_22_75 bit_22_75 bitb_22_75 word22_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_75 q_23_75 qb_23_75 bit_23_75 bitb_23_75 word23_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_75 q_24_75 qb_24_75 bit_24_75 bitb_24_75 word24_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_75 q_25_75 qb_25_75 bit_25_75 bitb_25_75 word25_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_75 q_26_75 qb_26_75 bit_26_75 bitb_26_75 word26_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_75 q_27_75 qb_27_75 bit_27_75 bitb_27_75 word27_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_75 q_28_75 qb_28_75 bit_28_75 bitb_28_75 word28_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_75 q_29_75 qb_29_75 bit_29_75 bitb_29_75 word29_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_75 q_30_75 qb_30_75 bit_30_75 bitb_30_75 word30_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_75 q_31_75 qb_31_75 bit_31_75 bitb_31_75 word31_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_75 q_32_75 qb_32_75 bit_32_75 bitb_32_75 word32_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_75 q_33_75 qb_33_75 bit_33_75 bitb_33_75 word33_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_75 q_34_75 qb_34_75 bit_34_75 bitb_34_75 word34_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_75 q_35_75 qb_35_75 bit_35_75 bitb_35_75 word35_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_75 q_36_75 qb_36_75 bit_36_75 bitb_36_75 word36_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_75 q_37_75 qb_37_75 bit_37_75 bitb_37_75 word37_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_75 q_38_75 qb_38_75 bit_38_75 bitb_38_75 word38_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_75 q_39_75 qb_39_75 bit_39_75 bitb_39_75 word39_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_75 q_40_75 qb_40_75 bit_40_75 bitb_40_75 word40_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_75 q_41_75 qb_41_75 bit_41_75 bitb_41_75 word41_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_75 q_42_75 qb_42_75 bit_42_75 bitb_42_75 word42_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_75 q_43_75 qb_43_75 bit_43_75 bitb_43_75 word43_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_75 q_44_75 qb_44_75 bit_44_75 bitb_44_75 word44_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_75 q_45_75 qb_45_75 bit_45_75 bitb_45_75 word45_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_75 q_46_75 qb_46_75 bit_46_75 bitb_46_75 word46_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_75 q_47_75 qb_47_75 bit_47_75 bitb_47_75 word47_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_75 q_48_75 qb_48_75 bit_48_75 bitb_48_75 word48_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_75 q_49_75 qb_49_75 bit_49_75 bitb_49_75 word49_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_75 q_50_75 qb_50_75 bit_50_75 bitb_50_75 word50_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_75 q_51_75 qb_51_75 bit_51_75 bitb_51_75 word51_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_75 q_52_75 qb_52_75 bit_52_75 bitb_52_75 word52_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_75 q_53_75 qb_53_75 bit_53_75 bitb_53_75 word53_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_75 q_54_75 qb_54_75 bit_54_75 bitb_54_75 word54_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_75 q_55_75 qb_55_75 bit_55_75 bitb_55_75 word55_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_75 q_56_75 qb_56_75 bit_56_75 bitb_56_75 word56_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_75 q_57_75 qb_57_75 bit_57_75 bitb_57_75 word57_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_75 q_58_75 qb_58_75 bit_58_75 bitb_58_75 word58_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_75 q_59_75 qb_59_75 bit_59_75 bitb_59_75 word59_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_75 q_60_75 qb_60_75 bit_60_75 bitb_60_75 word60_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_75 q_61_75 qb_61_75 bit_61_75 bitb_61_75 word61_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_75 q_62_75 qb_62_75 bit_62_75 bitb_62_75 word62_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_75 q_63_75 qb_63_75 bit_63_75 bitb_63_75 word63_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_75 q_64_75 qb_64_75 bit_64_75 bitb_64_75 word64_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_75 q_65_75 qb_65_75 bit_65_75 bitb_65_75 word65_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_75 q_66_75 qb_66_75 bit_66_75 bitb_66_75 word66_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_75 q_67_75 qb_67_75 bit_67_75 bitb_67_75 word67_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_75 q_68_75 qb_68_75 bit_68_75 bitb_68_75 word68_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_75 q_69_75 qb_69_75 bit_69_75 bitb_69_75 word69_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_75 q_70_75 qb_70_75 bit_70_75 bitb_70_75 word70_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_75 q_71_75 qb_71_75 bit_71_75 bitb_71_75 word71_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_75 q_72_75 qb_72_75 bit_72_75 bitb_72_75 word72_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_75 q_73_75 qb_73_75 bit_73_75 bitb_73_75 word73_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_75 q_74_75 qb_74_75 bit_74_75 bitb_74_75 word74_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_75 q_75_75 qb_75_75 bit_75_75 bitb_75_75 word75_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_75 q_76_75 qb_76_75 bit_76_75 bitb_76_75 word76_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_75 q_77_75 qb_77_75 bit_77_75 bitb_77_75 word77_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_75 q_78_75 qb_78_75 bit_78_75 bitb_78_75 word78_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_75 q_79_75 qb_79_75 bit_79_75 bitb_79_75 word79_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_75 q_80_75 qb_80_75 bit_80_75 bitb_80_75 word80_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_75 q_81_75 qb_81_75 bit_81_75 bitb_81_75 word81_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_75 q_82_75 qb_82_75 bit_82_75 bitb_82_75 word82_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_75 q_83_75 qb_83_75 bit_83_75 bitb_83_75 word83_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_75 q_84_75 qb_84_75 bit_84_75 bitb_84_75 word84_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_75 q_85_75 qb_85_75 bit_85_75 bitb_85_75 word85_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_75 q_86_75 qb_86_75 bit_86_75 bitb_86_75 word86_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_75 q_87_75 qb_87_75 bit_87_75 bitb_87_75 word87_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_75 q_88_75 qb_88_75 bit_88_75 bitb_88_75 word88_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_75 q_89_75 qb_89_75 bit_89_75 bitb_89_75 word89_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_75 q_90_75 qb_90_75 bit_90_75 bitb_90_75 word90_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_75 q_91_75 qb_91_75 bit_91_75 bitb_91_75 word91_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_75 q_92_75 qb_92_75 bit_92_75 bitb_92_75 word92_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_75 q_93_75 qb_93_75 bit_93_75 bitb_93_75 word93_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_75 q_94_75 qb_94_75 bit_94_75 bitb_94_75 word94_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_75 q_95_75 qb_95_75 bit_95_75 bitb_95_75 word95_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_75 q_96_75 qb_96_75 bit_96_75 bitb_96_75 word96_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_75 q_97_75 qb_97_75 bit_97_75 bitb_97_75 word97_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_75 q_98_75 qb_98_75 bit_98_75 bitb_98_75 word98_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_75 q_99_75 qb_99_75 bit_99_75 bitb_99_75 word99_75 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_76 q_0_76 qb_0_76 bit_0_76 bitb_0_76 word0_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_76 q_1_76 qb_1_76 bit_1_76 bitb_1_76 word1_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_76 q_2_76 qb_2_76 bit_2_76 bitb_2_76 word2_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_76 q_3_76 qb_3_76 bit_3_76 bitb_3_76 word3_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_76 q_4_76 qb_4_76 bit_4_76 bitb_4_76 word4_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_76 q_5_76 qb_5_76 bit_5_76 bitb_5_76 word5_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_76 q_6_76 qb_6_76 bit_6_76 bitb_6_76 word6_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_76 q_7_76 qb_7_76 bit_7_76 bitb_7_76 word7_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_76 q_8_76 qb_8_76 bit_8_76 bitb_8_76 word8_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_76 q_9_76 qb_9_76 bit_9_76 bitb_9_76 word9_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_76 q_10_76 qb_10_76 bit_10_76 bitb_10_76 word10_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_76 q_11_76 qb_11_76 bit_11_76 bitb_11_76 word11_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_76 q_12_76 qb_12_76 bit_12_76 bitb_12_76 word12_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_76 q_13_76 qb_13_76 bit_13_76 bitb_13_76 word13_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_76 q_14_76 qb_14_76 bit_14_76 bitb_14_76 word14_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_76 q_15_76 qb_15_76 bit_15_76 bitb_15_76 word15_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_76 q_16_76 qb_16_76 bit_16_76 bitb_16_76 word16_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_76 q_17_76 qb_17_76 bit_17_76 bitb_17_76 word17_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_76 q_18_76 qb_18_76 bit_18_76 bitb_18_76 word18_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_76 q_19_76 qb_19_76 bit_19_76 bitb_19_76 word19_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_76 q_20_76 qb_20_76 bit_20_76 bitb_20_76 word20_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_76 q_21_76 qb_21_76 bit_21_76 bitb_21_76 word21_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_76 q_22_76 qb_22_76 bit_22_76 bitb_22_76 word22_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_76 q_23_76 qb_23_76 bit_23_76 bitb_23_76 word23_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_76 q_24_76 qb_24_76 bit_24_76 bitb_24_76 word24_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_76 q_25_76 qb_25_76 bit_25_76 bitb_25_76 word25_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_76 q_26_76 qb_26_76 bit_26_76 bitb_26_76 word26_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_76 q_27_76 qb_27_76 bit_27_76 bitb_27_76 word27_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_76 q_28_76 qb_28_76 bit_28_76 bitb_28_76 word28_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_76 q_29_76 qb_29_76 bit_29_76 bitb_29_76 word29_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_76 q_30_76 qb_30_76 bit_30_76 bitb_30_76 word30_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_76 q_31_76 qb_31_76 bit_31_76 bitb_31_76 word31_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_76 q_32_76 qb_32_76 bit_32_76 bitb_32_76 word32_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_76 q_33_76 qb_33_76 bit_33_76 bitb_33_76 word33_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_76 q_34_76 qb_34_76 bit_34_76 bitb_34_76 word34_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_76 q_35_76 qb_35_76 bit_35_76 bitb_35_76 word35_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_76 q_36_76 qb_36_76 bit_36_76 bitb_36_76 word36_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_76 q_37_76 qb_37_76 bit_37_76 bitb_37_76 word37_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_76 q_38_76 qb_38_76 bit_38_76 bitb_38_76 word38_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_76 q_39_76 qb_39_76 bit_39_76 bitb_39_76 word39_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_76 q_40_76 qb_40_76 bit_40_76 bitb_40_76 word40_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_76 q_41_76 qb_41_76 bit_41_76 bitb_41_76 word41_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_76 q_42_76 qb_42_76 bit_42_76 bitb_42_76 word42_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_76 q_43_76 qb_43_76 bit_43_76 bitb_43_76 word43_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_76 q_44_76 qb_44_76 bit_44_76 bitb_44_76 word44_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_76 q_45_76 qb_45_76 bit_45_76 bitb_45_76 word45_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_76 q_46_76 qb_46_76 bit_46_76 bitb_46_76 word46_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_76 q_47_76 qb_47_76 bit_47_76 bitb_47_76 word47_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_76 q_48_76 qb_48_76 bit_48_76 bitb_48_76 word48_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_76 q_49_76 qb_49_76 bit_49_76 bitb_49_76 word49_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_76 q_50_76 qb_50_76 bit_50_76 bitb_50_76 word50_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_76 q_51_76 qb_51_76 bit_51_76 bitb_51_76 word51_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_76 q_52_76 qb_52_76 bit_52_76 bitb_52_76 word52_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_76 q_53_76 qb_53_76 bit_53_76 bitb_53_76 word53_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_76 q_54_76 qb_54_76 bit_54_76 bitb_54_76 word54_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_76 q_55_76 qb_55_76 bit_55_76 bitb_55_76 word55_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_76 q_56_76 qb_56_76 bit_56_76 bitb_56_76 word56_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_76 q_57_76 qb_57_76 bit_57_76 bitb_57_76 word57_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_76 q_58_76 qb_58_76 bit_58_76 bitb_58_76 word58_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_76 q_59_76 qb_59_76 bit_59_76 bitb_59_76 word59_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_76 q_60_76 qb_60_76 bit_60_76 bitb_60_76 word60_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_76 q_61_76 qb_61_76 bit_61_76 bitb_61_76 word61_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_76 q_62_76 qb_62_76 bit_62_76 bitb_62_76 word62_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_76 q_63_76 qb_63_76 bit_63_76 bitb_63_76 word63_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_76 q_64_76 qb_64_76 bit_64_76 bitb_64_76 word64_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_76 q_65_76 qb_65_76 bit_65_76 bitb_65_76 word65_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_76 q_66_76 qb_66_76 bit_66_76 bitb_66_76 word66_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_76 q_67_76 qb_67_76 bit_67_76 bitb_67_76 word67_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_76 q_68_76 qb_68_76 bit_68_76 bitb_68_76 word68_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_76 q_69_76 qb_69_76 bit_69_76 bitb_69_76 word69_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_76 q_70_76 qb_70_76 bit_70_76 bitb_70_76 word70_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_76 q_71_76 qb_71_76 bit_71_76 bitb_71_76 word71_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_76 q_72_76 qb_72_76 bit_72_76 bitb_72_76 word72_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_76 q_73_76 qb_73_76 bit_73_76 bitb_73_76 word73_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_76 q_74_76 qb_74_76 bit_74_76 bitb_74_76 word74_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_76 q_75_76 qb_75_76 bit_75_76 bitb_75_76 word75_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_76 q_76_76 qb_76_76 bit_76_76 bitb_76_76 word76_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_76 q_77_76 qb_77_76 bit_77_76 bitb_77_76 word77_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_76 q_78_76 qb_78_76 bit_78_76 bitb_78_76 word78_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_76 q_79_76 qb_79_76 bit_79_76 bitb_79_76 word79_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_76 q_80_76 qb_80_76 bit_80_76 bitb_80_76 word80_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_76 q_81_76 qb_81_76 bit_81_76 bitb_81_76 word81_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_76 q_82_76 qb_82_76 bit_82_76 bitb_82_76 word82_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_76 q_83_76 qb_83_76 bit_83_76 bitb_83_76 word83_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_76 q_84_76 qb_84_76 bit_84_76 bitb_84_76 word84_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_76 q_85_76 qb_85_76 bit_85_76 bitb_85_76 word85_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_76 q_86_76 qb_86_76 bit_86_76 bitb_86_76 word86_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_76 q_87_76 qb_87_76 bit_87_76 bitb_87_76 word87_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_76 q_88_76 qb_88_76 bit_88_76 bitb_88_76 word88_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_76 q_89_76 qb_89_76 bit_89_76 bitb_89_76 word89_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_76 q_90_76 qb_90_76 bit_90_76 bitb_90_76 word90_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_76 q_91_76 qb_91_76 bit_91_76 bitb_91_76 word91_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_76 q_92_76 qb_92_76 bit_92_76 bitb_92_76 word92_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_76 q_93_76 qb_93_76 bit_93_76 bitb_93_76 word93_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_76 q_94_76 qb_94_76 bit_94_76 bitb_94_76 word94_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_76 q_95_76 qb_95_76 bit_95_76 bitb_95_76 word95_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_76 q_96_76 qb_96_76 bit_96_76 bitb_96_76 word96_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_76 q_97_76 qb_97_76 bit_97_76 bitb_97_76 word97_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_76 q_98_76 qb_98_76 bit_98_76 bitb_98_76 word98_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_76 q_99_76 qb_99_76 bit_99_76 bitb_99_76 word99_76 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_77 q_0_77 qb_0_77 bit_0_77 bitb_0_77 word0_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_77 q_1_77 qb_1_77 bit_1_77 bitb_1_77 word1_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_77 q_2_77 qb_2_77 bit_2_77 bitb_2_77 word2_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_77 q_3_77 qb_3_77 bit_3_77 bitb_3_77 word3_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_77 q_4_77 qb_4_77 bit_4_77 bitb_4_77 word4_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_77 q_5_77 qb_5_77 bit_5_77 bitb_5_77 word5_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_77 q_6_77 qb_6_77 bit_6_77 bitb_6_77 word6_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_77 q_7_77 qb_7_77 bit_7_77 bitb_7_77 word7_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_77 q_8_77 qb_8_77 bit_8_77 bitb_8_77 word8_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_77 q_9_77 qb_9_77 bit_9_77 bitb_9_77 word9_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_77 q_10_77 qb_10_77 bit_10_77 bitb_10_77 word10_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_77 q_11_77 qb_11_77 bit_11_77 bitb_11_77 word11_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_77 q_12_77 qb_12_77 bit_12_77 bitb_12_77 word12_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_77 q_13_77 qb_13_77 bit_13_77 bitb_13_77 word13_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_77 q_14_77 qb_14_77 bit_14_77 bitb_14_77 word14_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_77 q_15_77 qb_15_77 bit_15_77 bitb_15_77 word15_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_77 q_16_77 qb_16_77 bit_16_77 bitb_16_77 word16_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_77 q_17_77 qb_17_77 bit_17_77 bitb_17_77 word17_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_77 q_18_77 qb_18_77 bit_18_77 bitb_18_77 word18_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_77 q_19_77 qb_19_77 bit_19_77 bitb_19_77 word19_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_77 q_20_77 qb_20_77 bit_20_77 bitb_20_77 word20_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_77 q_21_77 qb_21_77 bit_21_77 bitb_21_77 word21_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_77 q_22_77 qb_22_77 bit_22_77 bitb_22_77 word22_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_77 q_23_77 qb_23_77 bit_23_77 bitb_23_77 word23_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_77 q_24_77 qb_24_77 bit_24_77 bitb_24_77 word24_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_77 q_25_77 qb_25_77 bit_25_77 bitb_25_77 word25_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_77 q_26_77 qb_26_77 bit_26_77 bitb_26_77 word26_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_77 q_27_77 qb_27_77 bit_27_77 bitb_27_77 word27_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_77 q_28_77 qb_28_77 bit_28_77 bitb_28_77 word28_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_77 q_29_77 qb_29_77 bit_29_77 bitb_29_77 word29_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_77 q_30_77 qb_30_77 bit_30_77 bitb_30_77 word30_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_77 q_31_77 qb_31_77 bit_31_77 bitb_31_77 word31_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_77 q_32_77 qb_32_77 bit_32_77 bitb_32_77 word32_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_77 q_33_77 qb_33_77 bit_33_77 bitb_33_77 word33_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_77 q_34_77 qb_34_77 bit_34_77 bitb_34_77 word34_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_77 q_35_77 qb_35_77 bit_35_77 bitb_35_77 word35_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_77 q_36_77 qb_36_77 bit_36_77 bitb_36_77 word36_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_77 q_37_77 qb_37_77 bit_37_77 bitb_37_77 word37_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_77 q_38_77 qb_38_77 bit_38_77 bitb_38_77 word38_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_77 q_39_77 qb_39_77 bit_39_77 bitb_39_77 word39_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_77 q_40_77 qb_40_77 bit_40_77 bitb_40_77 word40_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_77 q_41_77 qb_41_77 bit_41_77 bitb_41_77 word41_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_77 q_42_77 qb_42_77 bit_42_77 bitb_42_77 word42_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_77 q_43_77 qb_43_77 bit_43_77 bitb_43_77 word43_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_77 q_44_77 qb_44_77 bit_44_77 bitb_44_77 word44_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_77 q_45_77 qb_45_77 bit_45_77 bitb_45_77 word45_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_77 q_46_77 qb_46_77 bit_46_77 bitb_46_77 word46_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_77 q_47_77 qb_47_77 bit_47_77 bitb_47_77 word47_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_77 q_48_77 qb_48_77 bit_48_77 bitb_48_77 word48_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_77 q_49_77 qb_49_77 bit_49_77 bitb_49_77 word49_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_77 q_50_77 qb_50_77 bit_50_77 bitb_50_77 word50_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_77 q_51_77 qb_51_77 bit_51_77 bitb_51_77 word51_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_77 q_52_77 qb_52_77 bit_52_77 bitb_52_77 word52_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_77 q_53_77 qb_53_77 bit_53_77 bitb_53_77 word53_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_77 q_54_77 qb_54_77 bit_54_77 bitb_54_77 word54_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_77 q_55_77 qb_55_77 bit_55_77 bitb_55_77 word55_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_77 q_56_77 qb_56_77 bit_56_77 bitb_56_77 word56_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_77 q_57_77 qb_57_77 bit_57_77 bitb_57_77 word57_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_77 q_58_77 qb_58_77 bit_58_77 bitb_58_77 word58_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_77 q_59_77 qb_59_77 bit_59_77 bitb_59_77 word59_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_77 q_60_77 qb_60_77 bit_60_77 bitb_60_77 word60_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_77 q_61_77 qb_61_77 bit_61_77 bitb_61_77 word61_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_77 q_62_77 qb_62_77 bit_62_77 bitb_62_77 word62_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_77 q_63_77 qb_63_77 bit_63_77 bitb_63_77 word63_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_77 q_64_77 qb_64_77 bit_64_77 bitb_64_77 word64_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_77 q_65_77 qb_65_77 bit_65_77 bitb_65_77 word65_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_77 q_66_77 qb_66_77 bit_66_77 bitb_66_77 word66_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_77 q_67_77 qb_67_77 bit_67_77 bitb_67_77 word67_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_77 q_68_77 qb_68_77 bit_68_77 bitb_68_77 word68_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_77 q_69_77 qb_69_77 bit_69_77 bitb_69_77 word69_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_77 q_70_77 qb_70_77 bit_70_77 bitb_70_77 word70_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_77 q_71_77 qb_71_77 bit_71_77 bitb_71_77 word71_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_77 q_72_77 qb_72_77 bit_72_77 bitb_72_77 word72_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_77 q_73_77 qb_73_77 bit_73_77 bitb_73_77 word73_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_77 q_74_77 qb_74_77 bit_74_77 bitb_74_77 word74_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_77 q_75_77 qb_75_77 bit_75_77 bitb_75_77 word75_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_77 q_76_77 qb_76_77 bit_76_77 bitb_76_77 word76_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_77 q_77_77 qb_77_77 bit_77_77 bitb_77_77 word77_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_77 q_78_77 qb_78_77 bit_78_77 bitb_78_77 word78_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_77 q_79_77 qb_79_77 bit_79_77 bitb_79_77 word79_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_77 q_80_77 qb_80_77 bit_80_77 bitb_80_77 word80_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_77 q_81_77 qb_81_77 bit_81_77 bitb_81_77 word81_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_77 q_82_77 qb_82_77 bit_82_77 bitb_82_77 word82_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_77 q_83_77 qb_83_77 bit_83_77 bitb_83_77 word83_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_77 q_84_77 qb_84_77 bit_84_77 bitb_84_77 word84_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_77 q_85_77 qb_85_77 bit_85_77 bitb_85_77 word85_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_77 q_86_77 qb_86_77 bit_86_77 bitb_86_77 word86_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_77 q_87_77 qb_87_77 bit_87_77 bitb_87_77 word87_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_77 q_88_77 qb_88_77 bit_88_77 bitb_88_77 word88_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_77 q_89_77 qb_89_77 bit_89_77 bitb_89_77 word89_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_77 q_90_77 qb_90_77 bit_90_77 bitb_90_77 word90_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_77 q_91_77 qb_91_77 bit_91_77 bitb_91_77 word91_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_77 q_92_77 qb_92_77 bit_92_77 bitb_92_77 word92_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_77 q_93_77 qb_93_77 bit_93_77 bitb_93_77 word93_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_77 q_94_77 qb_94_77 bit_94_77 bitb_94_77 word94_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_77 q_95_77 qb_95_77 bit_95_77 bitb_95_77 word95_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_77 q_96_77 qb_96_77 bit_96_77 bitb_96_77 word96_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_77 q_97_77 qb_97_77 bit_97_77 bitb_97_77 word97_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_77 q_98_77 qb_98_77 bit_98_77 bitb_98_77 word98_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_77 q_99_77 qb_99_77 bit_99_77 bitb_99_77 word99_77 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_78 q_0_78 qb_0_78 bit_0_78 bitb_0_78 word0_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_78 q_1_78 qb_1_78 bit_1_78 bitb_1_78 word1_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_78 q_2_78 qb_2_78 bit_2_78 bitb_2_78 word2_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_78 q_3_78 qb_3_78 bit_3_78 bitb_3_78 word3_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_78 q_4_78 qb_4_78 bit_4_78 bitb_4_78 word4_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_78 q_5_78 qb_5_78 bit_5_78 bitb_5_78 word5_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_78 q_6_78 qb_6_78 bit_6_78 bitb_6_78 word6_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_78 q_7_78 qb_7_78 bit_7_78 bitb_7_78 word7_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_78 q_8_78 qb_8_78 bit_8_78 bitb_8_78 word8_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_78 q_9_78 qb_9_78 bit_9_78 bitb_9_78 word9_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_78 q_10_78 qb_10_78 bit_10_78 bitb_10_78 word10_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_78 q_11_78 qb_11_78 bit_11_78 bitb_11_78 word11_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_78 q_12_78 qb_12_78 bit_12_78 bitb_12_78 word12_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_78 q_13_78 qb_13_78 bit_13_78 bitb_13_78 word13_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_78 q_14_78 qb_14_78 bit_14_78 bitb_14_78 word14_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_78 q_15_78 qb_15_78 bit_15_78 bitb_15_78 word15_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_78 q_16_78 qb_16_78 bit_16_78 bitb_16_78 word16_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_78 q_17_78 qb_17_78 bit_17_78 bitb_17_78 word17_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_78 q_18_78 qb_18_78 bit_18_78 bitb_18_78 word18_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_78 q_19_78 qb_19_78 bit_19_78 bitb_19_78 word19_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_78 q_20_78 qb_20_78 bit_20_78 bitb_20_78 word20_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_78 q_21_78 qb_21_78 bit_21_78 bitb_21_78 word21_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_78 q_22_78 qb_22_78 bit_22_78 bitb_22_78 word22_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_78 q_23_78 qb_23_78 bit_23_78 bitb_23_78 word23_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_78 q_24_78 qb_24_78 bit_24_78 bitb_24_78 word24_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_78 q_25_78 qb_25_78 bit_25_78 bitb_25_78 word25_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_78 q_26_78 qb_26_78 bit_26_78 bitb_26_78 word26_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_78 q_27_78 qb_27_78 bit_27_78 bitb_27_78 word27_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_78 q_28_78 qb_28_78 bit_28_78 bitb_28_78 word28_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_78 q_29_78 qb_29_78 bit_29_78 bitb_29_78 word29_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_78 q_30_78 qb_30_78 bit_30_78 bitb_30_78 word30_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_78 q_31_78 qb_31_78 bit_31_78 bitb_31_78 word31_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_78 q_32_78 qb_32_78 bit_32_78 bitb_32_78 word32_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_78 q_33_78 qb_33_78 bit_33_78 bitb_33_78 word33_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_78 q_34_78 qb_34_78 bit_34_78 bitb_34_78 word34_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_78 q_35_78 qb_35_78 bit_35_78 bitb_35_78 word35_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_78 q_36_78 qb_36_78 bit_36_78 bitb_36_78 word36_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_78 q_37_78 qb_37_78 bit_37_78 bitb_37_78 word37_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_78 q_38_78 qb_38_78 bit_38_78 bitb_38_78 word38_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_78 q_39_78 qb_39_78 bit_39_78 bitb_39_78 word39_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_78 q_40_78 qb_40_78 bit_40_78 bitb_40_78 word40_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_78 q_41_78 qb_41_78 bit_41_78 bitb_41_78 word41_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_78 q_42_78 qb_42_78 bit_42_78 bitb_42_78 word42_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_78 q_43_78 qb_43_78 bit_43_78 bitb_43_78 word43_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_78 q_44_78 qb_44_78 bit_44_78 bitb_44_78 word44_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_78 q_45_78 qb_45_78 bit_45_78 bitb_45_78 word45_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_78 q_46_78 qb_46_78 bit_46_78 bitb_46_78 word46_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_78 q_47_78 qb_47_78 bit_47_78 bitb_47_78 word47_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_78 q_48_78 qb_48_78 bit_48_78 bitb_48_78 word48_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_78 q_49_78 qb_49_78 bit_49_78 bitb_49_78 word49_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_78 q_50_78 qb_50_78 bit_50_78 bitb_50_78 word50_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_78 q_51_78 qb_51_78 bit_51_78 bitb_51_78 word51_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_78 q_52_78 qb_52_78 bit_52_78 bitb_52_78 word52_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_78 q_53_78 qb_53_78 bit_53_78 bitb_53_78 word53_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_78 q_54_78 qb_54_78 bit_54_78 bitb_54_78 word54_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_78 q_55_78 qb_55_78 bit_55_78 bitb_55_78 word55_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_78 q_56_78 qb_56_78 bit_56_78 bitb_56_78 word56_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_78 q_57_78 qb_57_78 bit_57_78 bitb_57_78 word57_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_78 q_58_78 qb_58_78 bit_58_78 bitb_58_78 word58_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_78 q_59_78 qb_59_78 bit_59_78 bitb_59_78 word59_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_78 q_60_78 qb_60_78 bit_60_78 bitb_60_78 word60_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_78 q_61_78 qb_61_78 bit_61_78 bitb_61_78 word61_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_78 q_62_78 qb_62_78 bit_62_78 bitb_62_78 word62_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_78 q_63_78 qb_63_78 bit_63_78 bitb_63_78 word63_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_78 q_64_78 qb_64_78 bit_64_78 bitb_64_78 word64_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_78 q_65_78 qb_65_78 bit_65_78 bitb_65_78 word65_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_78 q_66_78 qb_66_78 bit_66_78 bitb_66_78 word66_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_78 q_67_78 qb_67_78 bit_67_78 bitb_67_78 word67_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_78 q_68_78 qb_68_78 bit_68_78 bitb_68_78 word68_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_78 q_69_78 qb_69_78 bit_69_78 bitb_69_78 word69_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_78 q_70_78 qb_70_78 bit_70_78 bitb_70_78 word70_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_78 q_71_78 qb_71_78 bit_71_78 bitb_71_78 word71_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_78 q_72_78 qb_72_78 bit_72_78 bitb_72_78 word72_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_78 q_73_78 qb_73_78 bit_73_78 bitb_73_78 word73_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_78 q_74_78 qb_74_78 bit_74_78 bitb_74_78 word74_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_78 q_75_78 qb_75_78 bit_75_78 bitb_75_78 word75_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_78 q_76_78 qb_76_78 bit_76_78 bitb_76_78 word76_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_78 q_77_78 qb_77_78 bit_77_78 bitb_77_78 word77_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_78 q_78_78 qb_78_78 bit_78_78 bitb_78_78 word78_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_78 q_79_78 qb_79_78 bit_79_78 bitb_79_78 word79_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_78 q_80_78 qb_80_78 bit_80_78 bitb_80_78 word80_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_78 q_81_78 qb_81_78 bit_81_78 bitb_81_78 word81_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_78 q_82_78 qb_82_78 bit_82_78 bitb_82_78 word82_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_78 q_83_78 qb_83_78 bit_83_78 bitb_83_78 word83_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_78 q_84_78 qb_84_78 bit_84_78 bitb_84_78 word84_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_78 q_85_78 qb_85_78 bit_85_78 bitb_85_78 word85_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_78 q_86_78 qb_86_78 bit_86_78 bitb_86_78 word86_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_78 q_87_78 qb_87_78 bit_87_78 bitb_87_78 word87_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_78 q_88_78 qb_88_78 bit_88_78 bitb_88_78 word88_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_78 q_89_78 qb_89_78 bit_89_78 bitb_89_78 word89_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_78 q_90_78 qb_90_78 bit_90_78 bitb_90_78 word90_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_78 q_91_78 qb_91_78 bit_91_78 bitb_91_78 word91_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_78 q_92_78 qb_92_78 bit_92_78 bitb_92_78 word92_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_78 q_93_78 qb_93_78 bit_93_78 bitb_93_78 word93_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_78 q_94_78 qb_94_78 bit_94_78 bitb_94_78 word94_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_78 q_95_78 qb_95_78 bit_95_78 bitb_95_78 word95_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_78 q_96_78 qb_96_78 bit_96_78 bitb_96_78 word96_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_78 q_97_78 qb_97_78 bit_97_78 bitb_97_78 word97_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_78 q_98_78 qb_98_78 bit_98_78 bitb_98_78 word98_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_78 q_99_78 qb_99_78 bit_99_78 bitb_99_78 word99_78 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_79 q_0_79 qb_0_79 bit_0_79 bitb_0_79 word0_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_79 q_1_79 qb_1_79 bit_1_79 bitb_1_79 word1_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_79 q_2_79 qb_2_79 bit_2_79 bitb_2_79 word2_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_79 q_3_79 qb_3_79 bit_3_79 bitb_3_79 word3_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_79 q_4_79 qb_4_79 bit_4_79 bitb_4_79 word4_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_79 q_5_79 qb_5_79 bit_5_79 bitb_5_79 word5_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_79 q_6_79 qb_6_79 bit_6_79 bitb_6_79 word6_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_79 q_7_79 qb_7_79 bit_7_79 bitb_7_79 word7_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_79 q_8_79 qb_8_79 bit_8_79 bitb_8_79 word8_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_79 q_9_79 qb_9_79 bit_9_79 bitb_9_79 word9_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_79 q_10_79 qb_10_79 bit_10_79 bitb_10_79 word10_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_79 q_11_79 qb_11_79 bit_11_79 bitb_11_79 word11_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_79 q_12_79 qb_12_79 bit_12_79 bitb_12_79 word12_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_79 q_13_79 qb_13_79 bit_13_79 bitb_13_79 word13_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_79 q_14_79 qb_14_79 bit_14_79 bitb_14_79 word14_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_79 q_15_79 qb_15_79 bit_15_79 bitb_15_79 word15_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_79 q_16_79 qb_16_79 bit_16_79 bitb_16_79 word16_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_79 q_17_79 qb_17_79 bit_17_79 bitb_17_79 word17_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_79 q_18_79 qb_18_79 bit_18_79 bitb_18_79 word18_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_79 q_19_79 qb_19_79 bit_19_79 bitb_19_79 word19_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_79 q_20_79 qb_20_79 bit_20_79 bitb_20_79 word20_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_79 q_21_79 qb_21_79 bit_21_79 bitb_21_79 word21_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_79 q_22_79 qb_22_79 bit_22_79 bitb_22_79 word22_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_79 q_23_79 qb_23_79 bit_23_79 bitb_23_79 word23_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_79 q_24_79 qb_24_79 bit_24_79 bitb_24_79 word24_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_79 q_25_79 qb_25_79 bit_25_79 bitb_25_79 word25_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_79 q_26_79 qb_26_79 bit_26_79 bitb_26_79 word26_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_79 q_27_79 qb_27_79 bit_27_79 bitb_27_79 word27_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_79 q_28_79 qb_28_79 bit_28_79 bitb_28_79 word28_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_79 q_29_79 qb_29_79 bit_29_79 bitb_29_79 word29_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_79 q_30_79 qb_30_79 bit_30_79 bitb_30_79 word30_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_79 q_31_79 qb_31_79 bit_31_79 bitb_31_79 word31_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_79 q_32_79 qb_32_79 bit_32_79 bitb_32_79 word32_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_79 q_33_79 qb_33_79 bit_33_79 bitb_33_79 word33_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_79 q_34_79 qb_34_79 bit_34_79 bitb_34_79 word34_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_79 q_35_79 qb_35_79 bit_35_79 bitb_35_79 word35_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_79 q_36_79 qb_36_79 bit_36_79 bitb_36_79 word36_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_79 q_37_79 qb_37_79 bit_37_79 bitb_37_79 word37_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_79 q_38_79 qb_38_79 bit_38_79 bitb_38_79 word38_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_79 q_39_79 qb_39_79 bit_39_79 bitb_39_79 word39_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_79 q_40_79 qb_40_79 bit_40_79 bitb_40_79 word40_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_79 q_41_79 qb_41_79 bit_41_79 bitb_41_79 word41_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_79 q_42_79 qb_42_79 bit_42_79 bitb_42_79 word42_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_79 q_43_79 qb_43_79 bit_43_79 bitb_43_79 word43_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_79 q_44_79 qb_44_79 bit_44_79 bitb_44_79 word44_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_79 q_45_79 qb_45_79 bit_45_79 bitb_45_79 word45_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_79 q_46_79 qb_46_79 bit_46_79 bitb_46_79 word46_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_79 q_47_79 qb_47_79 bit_47_79 bitb_47_79 word47_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_79 q_48_79 qb_48_79 bit_48_79 bitb_48_79 word48_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_79 q_49_79 qb_49_79 bit_49_79 bitb_49_79 word49_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_79 q_50_79 qb_50_79 bit_50_79 bitb_50_79 word50_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_79 q_51_79 qb_51_79 bit_51_79 bitb_51_79 word51_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_79 q_52_79 qb_52_79 bit_52_79 bitb_52_79 word52_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_79 q_53_79 qb_53_79 bit_53_79 bitb_53_79 word53_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_79 q_54_79 qb_54_79 bit_54_79 bitb_54_79 word54_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_79 q_55_79 qb_55_79 bit_55_79 bitb_55_79 word55_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_79 q_56_79 qb_56_79 bit_56_79 bitb_56_79 word56_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_79 q_57_79 qb_57_79 bit_57_79 bitb_57_79 word57_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_79 q_58_79 qb_58_79 bit_58_79 bitb_58_79 word58_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_79 q_59_79 qb_59_79 bit_59_79 bitb_59_79 word59_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_79 q_60_79 qb_60_79 bit_60_79 bitb_60_79 word60_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_79 q_61_79 qb_61_79 bit_61_79 bitb_61_79 word61_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_79 q_62_79 qb_62_79 bit_62_79 bitb_62_79 word62_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_79 q_63_79 qb_63_79 bit_63_79 bitb_63_79 word63_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_79 q_64_79 qb_64_79 bit_64_79 bitb_64_79 word64_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_79 q_65_79 qb_65_79 bit_65_79 bitb_65_79 word65_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_79 q_66_79 qb_66_79 bit_66_79 bitb_66_79 word66_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_79 q_67_79 qb_67_79 bit_67_79 bitb_67_79 word67_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_79 q_68_79 qb_68_79 bit_68_79 bitb_68_79 word68_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_79 q_69_79 qb_69_79 bit_69_79 bitb_69_79 word69_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_79 q_70_79 qb_70_79 bit_70_79 bitb_70_79 word70_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_79 q_71_79 qb_71_79 bit_71_79 bitb_71_79 word71_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_79 q_72_79 qb_72_79 bit_72_79 bitb_72_79 word72_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_79 q_73_79 qb_73_79 bit_73_79 bitb_73_79 word73_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_79 q_74_79 qb_74_79 bit_74_79 bitb_74_79 word74_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_79 q_75_79 qb_75_79 bit_75_79 bitb_75_79 word75_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_79 q_76_79 qb_76_79 bit_76_79 bitb_76_79 word76_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_79 q_77_79 qb_77_79 bit_77_79 bitb_77_79 word77_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_79 q_78_79 qb_78_79 bit_78_79 bitb_78_79 word78_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_79 q_79_79 qb_79_79 bit_79_79 bitb_79_79 word79_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_79 q_80_79 qb_80_79 bit_80_79 bitb_80_79 word80_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_79 q_81_79 qb_81_79 bit_81_79 bitb_81_79 word81_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_79 q_82_79 qb_82_79 bit_82_79 bitb_82_79 word82_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_79 q_83_79 qb_83_79 bit_83_79 bitb_83_79 word83_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_79 q_84_79 qb_84_79 bit_84_79 bitb_84_79 word84_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_79 q_85_79 qb_85_79 bit_85_79 bitb_85_79 word85_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_79 q_86_79 qb_86_79 bit_86_79 bitb_86_79 word86_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_79 q_87_79 qb_87_79 bit_87_79 bitb_87_79 word87_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_79 q_88_79 qb_88_79 bit_88_79 bitb_88_79 word88_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_79 q_89_79 qb_89_79 bit_89_79 bitb_89_79 word89_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_79 q_90_79 qb_90_79 bit_90_79 bitb_90_79 word90_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_79 q_91_79 qb_91_79 bit_91_79 bitb_91_79 word91_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_79 q_92_79 qb_92_79 bit_92_79 bitb_92_79 word92_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_79 q_93_79 qb_93_79 bit_93_79 bitb_93_79 word93_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_79 q_94_79 qb_94_79 bit_94_79 bitb_94_79 word94_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_79 q_95_79 qb_95_79 bit_95_79 bitb_95_79 word95_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_79 q_96_79 qb_96_79 bit_96_79 bitb_96_79 word96_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_79 q_97_79 qb_97_79 bit_97_79 bitb_97_79 word97_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_79 q_98_79 qb_98_79 bit_98_79 bitb_98_79 word98_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_79 q_99_79 qb_99_79 bit_99_79 bitb_99_79 word99_79 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_80 q_0_80 qb_0_80 bit_0_80 bitb_0_80 word0_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_80 q_1_80 qb_1_80 bit_1_80 bitb_1_80 word1_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_80 q_2_80 qb_2_80 bit_2_80 bitb_2_80 word2_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_80 q_3_80 qb_3_80 bit_3_80 bitb_3_80 word3_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_80 q_4_80 qb_4_80 bit_4_80 bitb_4_80 word4_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_80 q_5_80 qb_5_80 bit_5_80 bitb_5_80 word5_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_80 q_6_80 qb_6_80 bit_6_80 bitb_6_80 word6_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_80 q_7_80 qb_7_80 bit_7_80 bitb_7_80 word7_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_80 q_8_80 qb_8_80 bit_8_80 bitb_8_80 word8_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_80 q_9_80 qb_9_80 bit_9_80 bitb_9_80 word9_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_80 q_10_80 qb_10_80 bit_10_80 bitb_10_80 word10_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_80 q_11_80 qb_11_80 bit_11_80 bitb_11_80 word11_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_80 q_12_80 qb_12_80 bit_12_80 bitb_12_80 word12_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_80 q_13_80 qb_13_80 bit_13_80 bitb_13_80 word13_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_80 q_14_80 qb_14_80 bit_14_80 bitb_14_80 word14_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_80 q_15_80 qb_15_80 bit_15_80 bitb_15_80 word15_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_80 q_16_80 qb_16_80 bit_16_80 bitb_16_80 word16_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_80 q_17_80 qb_17_80 bit_17_80 bitb_17_80 word17_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_80 q_18_80 qb_18_80 bit_18_80 bitb_18_80 word18_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_80 q_19_80 qb_19_80 bit_19_80 bitb_19_80 word19_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_80 q_20_80 qb_20_80 bit_20_80 bitb_20_80 word20_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_80 q_21_80 qb_21_80 bit_21_80 bitb_21_80 word21_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_80 q_22_80 qb_22_80 bit_22_80 bitb_22_80 word22_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_80 q_23_80 qb_23_80 bit_23_80 bitb_23_80 word23_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_80 q_24_80 qb_24_80 bit_24_80 bitb_24_80 word24_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_80 q_25_80 qb_25_80 bit_25_80 bitb_25_80 word25_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_80 q_26_80 qb_26_80 bit_26_80 bitb_26_80 word26_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_80 q_27_80 qb_27_80 bit_27_80 bitb_27_80 word27_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_80 q_28_80 qb_28_80 bit_28_80 bitb_28_80 word28_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_80 q_29_80 qb_29_80 bit_29_80 bitb_29_80 word29_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_80 q_30_80 qb_30_80 bit_30_80 bitb_30_80 word30_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_80 q_31_80 qb_31_80 bit_31_80 bitb_31_80 word31_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_80 q_32_80 qb_32_80 bit_32_80 bitb_32_80 word32_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_80 q_33_80 qb_33_80 bit_33_80 bitb_33_80 word33_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_80 q_34_80 qb_34_80 bit_34_80 bitb_34_80 word34_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_80 q_35_80 qb_35_80 bit_35_80 bitb_35_80 word35_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_80 q_36_80 qb_36_80 bit_36_80 bitb_36_80 word36_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_80 q_37_80 qb_37_80 bit_37_80 bitb_37_80 word37_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_80 q_38_80 qb_38_80 bit_38_80 bitb_38_80 word38_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_80 q_39_80 qb_39_80 bit_39_80 bitb_39_80 word39_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_80 q_40_80 qb_40_80 bit_40_80 bitb_40_80 word40_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_80 q_41_80 qb_41_80 bit_41_80 bitb_41_80 word41_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_80 q_42_80 qb_42_80 bit_42_80 bitb_42_80 word42_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_80 q_43_80 qb_43_80 bit_43_80 bitb_43_80 word43_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_80 q_44_80 qb_44_80 bit_44_80 bitb_44_80 word44_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_80 q_45_80 qb_45_80 bit_45_80 bitb_45_80 word45_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_80 q_46_80 qb_46_80 bit_46_80 bitb_46_80 word46_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_80 q_47_80 qb_47_80 bit_47_80 bitb_47_80 word47_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_80 q_48_80 qb_48_80 bit_48_80 bitb_48_80 word48_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_80 q_49_80 qb_49_80 bit_49_80 bitb_49_80 word49_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_80 q_50_80 qb_50_80 bit_50_80 bitb_50_80 word50_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_80 q_51_80 qb_51_80 bit_51_80 bitb_51_80 word51_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_80 q_52_80 qb_52_80 bit_52_80 bitb_52_80 word52_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_80 q_53_80 qb_53_80 bit_53_80 bitb_53_80 word53_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_80 q_54_80 qb_54_80 bit_54_80 bitb_54_80 word54_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_80 q_55_80 qb_55_80 bit_55_80 bitb_55_80 word55_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_80 q_56_80 qb_56_80 bit_56_80 bitb_56_80 word56_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_80 q_57_80 qb_57_80 bit_57_80 bitb_57_80 word57_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_80 q_58_80 qb_58_80 bit_58_80 bitb_58_80 word58_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_80 q_59_80 qb_59_80 bit_59_80 bitb_59_80 word59_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_80 q_60_80 qb_60_80 bit_60_80 bitb_60_80 word60_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_80 q_61_80 qb_61_80 bit_61_80 bitb_61_80 word61_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_80 q_62_80 qb_62_80 bit_62_80 bitb_62_80 word62_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_80 q_63_80 qb_63_80 bit_63_80 bitb_63_80 word63_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_80 q_64_80 qb_64_80 bit_64_80 bitb_64_80 word64_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_80 q_65_80 qb_65_80 bit_65_80 bitb_65_80 word65_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_80 q_66_80 qb_66_80 bit_66_80 bitb_66_80 word66_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_80 q_67_80 qb_67_80 bit_67_80 bitb_67_80 word67_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_80 q_68_80 qb_68_80 bit_68_80 bitb_68_80 word68_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_80 q_69_80 qb_69_80 bit_69_80 bitb_69_80 word69_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_80 q_70_80 qb_70_80 bit_70_80 bitb_70_80 word70_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_80 q_71_80 qb_71_80 bit_71_80 bitb_71_80 word71_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_80 q_72_80 qb_72_80 bit_72_80 bitb_72_80 word72_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_80 q_73_80 qb_73_80 bit_73_80 bitb_73_80 word73_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_80 q_74_80 qb_74_80 bit_74_80 bitb_74_80 word74_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_80 q_75_80 qb_75_80 bit_75_80 bitb_75_80 word75_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_80 q_76_80 qb_76_80 bit_76_80 bitb_76_80 word76_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_80 q_77_80 qb_77_80 bit_77_80 bitb_77_80 word77_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_80 q_78_80 qb_78_80 bit_78_80 bitb_78_80 word78_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_80 q_79_80 qb_79_80 bit_79_80 bitb_79_80 word79_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_80 q_80_80 qb_80_80 bit_80_80 bitb_80_80 word80_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_80 q_81_80 qb_81_80 bit_81_80 bitb_81_80 word81_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_80 q_82_80 qb_82_80 bit_82_80 bitb_82_80 word82_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_80 q_83_80 qb_83_80 bit_83_80 bitb_83_80 word83_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_80 q_84_80 qb_84_80 bit_84_80 bitb_84_80 word84_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_80 q_85_80 qb_85_80 bit_85_80 bitb_85_80 word85_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_80 q_86_80 qb_86_80 bit_86_80 bitb_86_80 word86_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_80 q_87_80 qb_87_80 bit_87_80 bitb_87_80 word87_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_80 q_88_80 qb_88_80 bit_88_80 bitb_88_80 word88_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_80 q_89_80 qb_89_80 bit_89_80 bitb_89_80 word89_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_80 q_90_80 qb_90_80 bit_90_80 bitb_90_80 word90_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_80 q_91_80 qb_91_80 bit_91_80 bitb_91_80 word91_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_80 q_92_80 qb_92_80 bit_92_80 bitb_92_80 word92_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_80 q_93_80 qb_93_80 bit_93_80 bitb_93_80 word93_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_80 q_94_80 qb_94_80 bit_94_80 bitb_94_80 word94_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_80 q_95_80 qb_95_80 bit_95_80 bitb_95_80 word95_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_80 q_96_80 qb_96_80 bit_96_80 bitb_96_80 word96_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_80 q_97_80 qb_97_80 bit_97_80 bitb_97_80 word97_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_80 q_98_80 qb_98_80 bit_98_80 bitb_98_80 word98_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_80 q_99_80 qb_99_80 bit_99_80 bitb_99_80 word99_80 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_81 q_0_81 qb_0_81 bit_0_81 bitb_0_81 word0_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_81 q_1_81 qb_1_81 bit_1_81 bitb_1_81 word1_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_81 q_2_81 qb_2_81 bit_2_81 bitb_2_81 word2_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_81 q_3_81 qb_3_81 bit_3_81 bitb_3_81 word3_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_81 q_4_81 qb_4_81 bit_4_81 bitb_4_81 word4_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_81 q_5_81 qb_5_81 bit_5_81 bitb_5_81 word5_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_81 q_6_81 qb_6_81 bit_6_81 bitb_6_81 word6_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_81 q_7_81 qb_7_81 bit_7_81 bitb_7_81 word7_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_81 q_8_81 qb_8_81 bit_8_81 bitb_8_81 word8_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_81 q_9_81 qb_9_81 bit_9_81 bitb_9_81 word9_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_81 q_10_81 qb_10_81 bit_10_81 bitb_10_81 word10_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_81 q_11_81 qb_11_81 bit_11_81 bitb_11_81 word11_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_81 q_12_81 qb_12_81 bit_12_81 bitb_12_81 word12_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_81 q_13_81 qb_13_81 bit_13_81 bitb_13_81 word13_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_81 q_14_81 qb_14_81 bit_14_81 bitb_14_81 word14_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_81 q_15_81 qb_15_81 bit_15_81 bitb_15_81 word15_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_81 q_16_81 qb_16_81 bit_16_81 bitb_16_81 word16_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_81 q_17_81 qb_17_81 bit_17_81 bitb_17_81 word17_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_81 q_18_81 qb_18_81 bit_18_81 bitb_18_81 word18_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_81 q_19_81 qb_19_81 bit_19_81 bitb_19_81 word19_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_81 q_20_81 qb_20_81 bit_20_81 bitb_20_81 word20_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_81 q_21_81 qb_21_81 bit_21_81 bitb_21_81 word21_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_81 q_22_81 qb_22_81 bit_22_81 bitb_22_81 word22_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_81 q_23_81 qb_23_81 bit_23_81 bitb_23_81 word23_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_81 q_24_81 qb_24_81 bit_24_81 bitb_24_81 word24_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_81 q_25_81 qb_25_81 bit_25_81 bitb_25_81 word25_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_81 q_26_81 qb_26_81 bit_26_81 bitb_26_81 word26_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_81 q_27_81 qb_27_81 bit_27_81 bitb_27_81 word27_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_81 q_28_81 qb_28_81 bit_28_81 bitb_28_81 word28_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_81 q_29_81 qb_29_81 bit_29_81 bitb_29_81 word29_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_81 q_30_81 qb_30_81 bit_30_81 bitb_30_81 word30_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_81 q_31_81 qb_31_81 bit_31_81 bitb_31_81 word31_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_81 q_32_81 qb_32_81 bit_32_81 bitb_32_81 word32_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_81 q_33_81 qb_33_81 bit_33_81 bitb_33_81 word33_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_81 q_34_81 qb_34_81 bit_34_81 bitb_34_81 word34_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_81 q_35_81 qb_35_81 bit_35_81 bitb_35_81 word35_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_81 q_36_81 qb_36_81 bit_36_81 bitb_36_81 word36_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_81 q_37_81 qb_37_81 bit_37_81 bitb_37_81 word37_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_81 q_38_81 qb_38_81 bit_38_81 bitb_38_81 word38_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_81 q_39_81 qb_39_81 bit_39_81 bitb_39_81 word39_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_81 q_40_81 qb_40_81 bit_40_81 bitb_40_81 word40_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_81 q_41_81 qb_41_81 bit_41_81 bitb_41_81 word41_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_81 q_42_81 qb_42_81 bit_42_81 bitb_42_81 word42_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_81 q_43_81 qb_43_81 bit_43_81 bitb_43_81 word43_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_81 q_44_81 qb_44_81 bit_44_81 bitb_44_81 word44_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_81 q_45_81 qb_45_81 bit_45_81 bitb_45_81 word45_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_81 q_46_81 qb_46_81 bit_46_81 bitb_46_81 word46_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_81 q_47_81 qb_47_81 bit_47_81 bitb_47_81 word47_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_81 q_48_81 qb_48_81 bit_48_81 bitb_48_81 word48_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_81 q_49_81 qb_49_81 bit_49_81 bitb_49_81 word49_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_81 q_50_81 qb_50_81 bit_50_81 bitb_50_81 word50_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_81 q_51_81 qb_51_81 bit_51_81 bitb_51_81 word51_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_81 q_52_81 qb_52_81 bit_52_81 bitb_52_81 word52_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_81 q_53_81 qb_53_81 bit_53_81 bitb_53_81 word53_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_81 q_54_81 qb_54_81 bit_54_81 bitb_54_81 word54_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_81 q_55_81 qb_55_81 bit_55_81 bitb_55_81 word55_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_81 q_56_81 qb_56_81 bit_56_81 bitb_56_81 word56_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_81 q_57_81 qb_57_81 bit_57_81 bitb_57_81 word57_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_81 q_58_81 qb_58_81 bit_58_81 bitb_58_81 word58_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_81 q_59_81 qb_59_81 bit_59_81 bitb_59_81 word59_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_81 q_60_81 qb_60_81 bit_60_81 bitb_60_81 word60_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_81 q_61_81 qb_61_81 bit_61_81 bitb_61_81 word61_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_81 q_62_81 qb_62_81 bit_62_81 bitb_62_81 word62_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_81 q_63_81 qb_63_81 bit_63_81 bitb_63_81 word63_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_81 q_64_81 qb_64_81 bit_64_81 bitb_64_81 word64_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_81 q_65_81 qb_65_81 bit_65_81 bitb_65_81 word65_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_81 q_66_81 qb_66_81 bit_66_81 bitb_66_81 word66_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_81 q_67_81 qb_67_81 bit_67_81 bitb_67_81 word67_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_81 q_68_81 qb_68_81 bit_68_81 bitb_68_81 word68_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_81 q_69_81 qb_69_81 bit_69_81 bitb_69_81 word69_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_81 q_70_81 qb_70_81 bit_70_81 bitb_70_81 word70_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_81 q_71_81 qb_71_81 bit_71_81 bitb_71_81 word71_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_81 q_72_81 qb_72_81 bit_72_81 bitb_72_81 word72_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_81 q_73_81 qb_73_81 bit_73_81 bitb_73_81 word73_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_81 q_74_81 qb_74_81 bit_74_81 bitb_74_81 word74_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_81 q_75_81 qb_75_81 bit_75_81 bitb_75_81 word75_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_81 q_76_81 qb_76_81 bit_76_81 bitb_76_81 word76_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_81 q_77_81 qb_77_81 bit_77_81 bitb_77_81 word77_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_81 q_78_81 qb_78_81 bit_78_81 bitb_78_81 word78_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_81 q_79_81 qb_79_81 bit_79_81 bitb_79_81 word79_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_81 q_80_81 qb_80_81 bit_80_81 bitb_80_81 word80_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_81 q_81_81 qb_81_81 bit_81_81 bitb_81_81 word81_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_81 q_82_81 qb_82_81 bit_82_81 bitb_82_81 word82_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_81 q_83_81 qb_83_81 bit_83_81 bitb_83_81 word83_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_81 q_84_81 qb_84_81 bit_84_81 bitb_84_81 word84_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_81 q_85_81 qb_85_81 bit_85_81 bitb_85_81 word85_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_81 q_86_81 qb_86_81 bit_86_81 bitb_86_81 word86_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_81 q_87_81 qb_87_81 bit_87_81 bitb_87_81 word87_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_81 q_88_81 qb_88_81 bit_88_81 bitb_88_81 word88_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_81 q_89_81 qb_89_81 bit_89_81 bitb_89_81 word89_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_81 q_90_81 qb_90_81 bit_90_81 bitb_90_81 word90_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_81 q_91_81 qb_91_81 bit_91_81 bitb_91_81 word91_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_81 q_92_81 qb_92_81 bit_92_81 bitb_92_81 word92_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_81 q_93_81 qb_93_81 bit_93_81 bitb_93_81 word93_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_81 q_94_81 qb_94_81 bit_94_81 bitb_94_81 word94_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_81 q_95_81 qb_95_81 bit_95_81 bitb_95_81 word95_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_81 q_96_81 qb_96_81 bit_96_81 bitb_96_81 word96_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_81 q_97_81 qb_97_81 bit_97_81 bitb_97_81 word97_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_81 q_98_81 qb_98_81 bit_98_81 bitb_98_81 word98_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_81 q_99_81 qb_99_81 bit_99_81 bitb_99_81 word99_81 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_82 q_0_82 qb_0_82 bit_0_82 bitb_0_82 word0_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_82 q_1_82 qb_1_82 bit_1_82 bitb_1_82 word1_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_82 q_2_82 qb_2_82 bit_2_82 bitb_2_82 word2_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_82 q_3_82 qb_3_82 bit_3_82 bitb_3_82 word3_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_82 q_4_82 qb_4_82 bit_4_82 bitb_4_82 word4_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_82 q_5_82 qb_5_82 bit_5_82 bitb_5_82 word5_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_82 q_6_82 qb_6_82 bit_6_82 bitb_6_82 word6_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_82 q_7_82 qb_7_82 bit_7_82 bitb_7_82 word7_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_82 q_8_82 qb_8_82 bit_8_82 bitb_8_82 word8_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_82 q_9_82 qb_9_82 bit_9_82 bitb_9_82 word9_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_82 q_10_82 qb_10_82 bit_10_82 bitb_10_82 word10_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_82 q_11_82 qb_11_82 bit_11_82 bitb_11_82 word11_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_82 q_12_82 qb_12_82 bit_12_82 bitb_12_82 word12_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_82 q_13_82 qb_13_82 bit_13_82 bitb_13_82 word13_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_82 q_14_82 qb_14_82 bit_14_82 bitb_14_82 word14_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_82 q_15_82 qb_15_82 bit_15_82 bitb_15_82 word15_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_82 q_16_82 qb_16_82 bit_16_82 bitb_16_82 word16_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_82 q_17_82 qb_17_82 bit_17_82 bitb_17_82 word17_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_82 q_18_82 qb_18_82 bit_18_82 bitb_18_82 word18_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_82 q_19_82 qb_19_82 bit_19_82 bitb_19_82 word19_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_82 q_20_82 qb_20_82 bit_20_82 bitb_20_82 word20_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_82 q_21_82 qb_21_82 bit_21_82 bitb_21_82 word21_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_82 q_22_82 qb_22_82 bit_22_82 bitb_22_82 word22_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_82 q_23_82 qb_23_82 bit_23_82 bitb_23_82 word23_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_82 q_24_82 qb_24_82 bit_24_82 bitb_24_82 word24_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_82 q_25_82 qb_25_82 bit_25_82 bitb_25_82 word25_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_82 q_26_82 qb_26_82 bit_26_82 bitb_26_82 word26_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_82 q_27_82 qb_27_82 bit_27_82 bitb_27_82 word27_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_82 q_28_82 qb_28_82 bit_28_82 bitb_28_82 word28_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_82 q_29_82 qb_29_82 bit_29_82 bitb_29_82 word29_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_82 q_30_82 qb_30_82 bit_30_82 bitb_30_82 word30_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_82 q_31_82 qb_31_82 bit_31_82 bitb_31_82 word31_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_82 q_32_82 qb_32_82 bit_32_82 bitb_32_82 word32_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_82 q_33_82 qb_33_82 bit_33_82 bitb_33_82 word33_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_82 q_34_82 qb_34_82 bit_34_82 bitb_34_82 word34_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_82 q_35_82 qb_35_82 bit_35_82 bitb_35_82 word35_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_82 q_36_82 qb_36_82 bit_36_82 bitb_36_82 word36_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_82 q_37_82 qb_37_82 bit_37_82 bitb_37_82 word37_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_82 q_38_82 qb_38_82 bit_38_82 bitb_38_82 word38_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_82 q_39_82 qb_39_82 bit_39_82 bitb_39_82 word39_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_82 q_40_82 qb_40_82 bit_40_82 bitb_40_82 word40_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_82 q_41_82 qb_41_82 bit_41_82 bitb_41_82 word41_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_82 q_42_82 qb_42_82 bit_42_82 bitb_42_82 word42_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_82 q_43_82 qb_43_82 bit_43_82 bitb_43_82 word43_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_82 q_44_82 qb_44_82 bit_44_82 bitb_44_82 word44_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_82 q_45_82 qb_45_82 bit_45_82 bitb_45_82 word45_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_82 q_46_82 qb_46_82 bit_46_82 bitb_46_82 word46_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_82 q_47_82 qb_47_82 bit_47_82 bitb_47_82 word47_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_82 q_48_82 qb_48_82 bit_48_82 bitb_48_82 word48_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_82 q_49_82 qb_49_82 bit_49_82 bitb_49_82 word49_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_82 q_50_82 qb_50_82 bit_50_82 bitb_50_82 word50_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_82 q_51_82 qb_51_82 bit_51_82 bitb_51_82 word51_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_82 q_52_82 qb_52_82 bit_52_82 bitb_52_82 word52_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_82 q_53_82 qb_53_82 bit_53_82 bitb_53_82 word53_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_82 q_54_82 qb_54_82 bit_54_82 bitb_54_82 word54_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_82 q_55_82 qb_55_82 bit_55_82 bitb_55_82 word55_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_82 q_56_82 qb_56_82 bit_56_82 bitb_56_82 word56_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_82 q_57_82 qb_57_82 bit_57_82 bitb_57_82 word57_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_82 q_58_82 qb_58_82 bit_58_82 bitb_58_82 word58_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_82 q_59_82 qb_59_82 bit_59_82 bitb_59_82 word59_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_82 q_60_82 qb_60_82 bit_60_82 bitb_60_82 word60_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_82 q_61_82 qb_61_82 bit_61_82 bitb_61_82 word61_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_82 q_62_82 qb_62_82 bit_62_82 bitb_62_82 word62_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_82 q_63_82 qb_63_82 bit_63_82 bitb_63_82 word63_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_82 q_64_82 qb_64_82 bit_64_82 bitb_64_82 word64_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_82 q_65_82 qb_65_82 bit_65_82 bitb_65_82 word65_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_82 q_66_82 qb_66_82 bit_66_82 bitb_66_82 word66_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_82 q_67_82 qb_67_82 bit_67_82 bitb_67_82 word67_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_82 q_68_82 qb_68_82 bit_68_82 bitb_68_82 word68_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_82 q_69_82 qb_69_82 bit_69_82 bitb_69_82 word69_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_82 q_70_82 qb_70_82 bit_70_82 bitb_70_82 word70_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_82 q_71_82 qb_71_82 bit_71_82 bitb_71_82 word71_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_82 q_72_82 qb_72_82 bit_72_82 bitb_72_82 word72_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_82 q_73_82 qb_73_82 bit_73_82 bitb_73_82 word73_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_82 q_74_82 qb_74_82 bit_74_82 bitb_74_82 word74_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_82 q_75_82 qb_75_82 bit_75_82 bitb_75_82 word75_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_82 q_76_82 qb_76_82 bit_76_82 bitb_76_82 word76_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_82 q_77_82 qb_77_82 bit_77_82 bitb_77_82 word77_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_82 q_78_82 qb_78_82 bit_78_82 bitb_78_82 word78_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_82 q_79_82 qb_79_82 bit_79_82 bitb_79_82 word79_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_82 q_80_82 qb_80_82 bit_80_82 bitb_80_82 word80_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_82 q_81_82 qb_81_82 bit_81_82 bitb_81_82 word81_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_82 q_82_82 qb_82_82 bit_82_82 bitb_82_82 word82_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_82 q_83_82 qb_83_82 bit_83_82 bitb_83_82 word83_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_82 q_84_82 qb_84_82 bit_84_82 bitb_84_82 word84_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_82 q_85_82 qb_85_82 bit_85_82 bitb_85_82 word85_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_82 q_86_82 qb_86_82 bit_86_82 bitb_86_82 word86_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_82 q_87_82 qb_87_82 bit_87_82 bitb_87_82 word87_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_82 q_88_82 qb_88_82 bit_88_82 bitb_88_82 word88_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_82 q_89_82 qb_89_82 bit_89_82 bitb_89_82 word89_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_82 q_90_82 qb_90_82 bit_90_82 bitb_90_82 word90_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_82 q_91_82 qb_91_82 bit_91_82 bitb_91_82 word91_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_82 q_92_82 qb_92_82 bit_92_82 bitb_92_82 word92_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_82 q_93_82 qb_93_82 bit_93_82 bitb_93_82 word93_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_82 q_94_82 qb_94_82 bit_94_82 bitb_94_82 word94_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_82 q_95_82 qb_95_82 bit_95_82 bitb_95_82 word95_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_82 q_96_82 qb_96_82 bit_96_82 bitb_96_82 word96_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_82 q_97_82 qb_97_82 bit_97_82 bitb_97_82 word97_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_82 q_98_82 qb_98_82 bit_98_82 bitb_98_82 word98_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_82 q_99_82 qb_99_82 bit_99_82 bitb_99_82 word99_82 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_83 q_0_83 qb_0_83 bit_0_83 bitb_0_83 word0_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_83 q_1_83 qb_1_83 bit_1_83 bitb_1_83 word1_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_83 q_2_83 qb_2_83 bit_2_83 bitb_2_83 word2_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_83 q_3_83 qb_3_83 bit_3_83 bitb_3_83 word3_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_83 q_4_83 qb_4_83 bit_4_83 bitb_4_83 word4_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_83 q_5_83 qb_5_83 bit_5_83 bitb_5_83 word5_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_83 q_6_83 qb_6_83 bit_6_83 bitb_6_83 word6_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_83 q_7_83 qb_7_83 bit_7_83 bitb_7_83 word7_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_83 q_8_83 qb_8_83 bit_8_83 bitb_8_83 word8_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_83 q_9_83 qb_9_83 bit_9_83 bitb_9_83 word9_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_83 q_10_83 qb_10_83 bit_10_83 bitb_10_83 word10_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_83 q_11_83 qb_11_83 bit_11_83 bitb_11_83 word11_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_83 q_12_83 qb_12_83 bit_12_83 bitb_12_83 word12_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_83 q_13_83 qb_13_83 bit_13_83 bitb_13_83 word13_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_83 q_14_83 qb_14_83 bit_14_83 bitb_14_83 word14_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_83 q_15_83 qb_15_83 bit_15_83 bitb_15_83 word15_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_83 q_16_83 qb_16_83 bit_16_83 bitb_16_83 word16_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_83 q_17_83 qb_17_83 bit_17_83 bitb_17_83 word17_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_83 q_18_83 qb_18_83 bit_18_83 bitb_18_83 word18_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_83 q_19_83 qb_19_83 bit_19_83 bitb_19_83 word19_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_83 q_20_83 qb_20_83 bit_20_83 bitb_20_83 word20_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_83 q_21_83 qb_21_83 bit_21_83 bitb_21_83 word21_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_83 q_22_83 qb_22_83 bit_22_83 bitb_22_83 word22_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_83 q_23_83 qb_23_83 bit_23_83 bitb_23_83 word23_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_83 q_24_83 qb_24_83 bit_24_83 bitb_24_83 word24_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_83 q_25_83 qb_25_83 bit_25_83 bitb_25_83 word25_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_83 q_26_83 qb_26_83 bit_26_83 bitb_26_83 word26_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_83 q_27_83 qb_27_83 bit_27_83 bitb_27_83 word27_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_83 q_28_83 qb_28_83 bit_28_83 bitb_28_83 word28_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_83 q_29_83 qb_29_83 bit_29_83 bitb_29_83 word29_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_83 q_30_83 qb_30_83 bit_30_83 bitb_30_83 word30_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_83 q_31_83 qb_31_83 bit_31_83 bitb_31_83 word31_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_83 q_32_83 qb_32_83 bit_32_83 bitb_32_83 word32_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_83 q_33_83 qb_33_83 bit_33_83 bitb_33_83 word33_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_83 q_34_83 qb_34_83 bit_34_83 bitb_34_83 word34_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_83 q_35_83 qb_35_83 bit_35_83 bitb_35_83 word35_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_83 q_36_83 qb_36_83 bit_36_83 bitb_36_83 word36_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_83 q_37_83 qb_37_83 bit_37_83 bitb_37_83 word37_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_83 q_38_83 qb_38_83 bit_38_83 bitb_38_83 word38_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_83 q_39_83 qb_39_83 bit_39_83 bitb_39_83 word39_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_83 q_40_83 qb_40_83 bit_40_83 bitb_40_83 word40_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_83 q_41_83 qb_41_83 bit_41_83 bitb_41_83 word41_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_83 q_42_83 qb_42_83 bit_42_83 bitb_42_83 word42_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_83 q_43_83 qb_43_83 bit_43_83 bitb_43_83 word43_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_83 q_44_83 qb_44_83 bit_44_83 bitb_44_83 word44_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_83 q_45_83 qb_45_83 bit_45_83 bitb_45_83 word45_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_83 q_46_83 qb_46_83 bit_46_83 bitb_46_83 word46_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_83 q_47_83 qb_47_83 bit_47_83 bitb_47_83 word47_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_83 q_48_83 qb_48_83 bit_48_83 bitb_48_83 word48_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_83 q_49_83 qb_49_83 bit_49_83 bitb_49_83 word49_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_83 q_50_83 qb_50_83 bit_50_83 bitb_50_83 word50_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_83 q_51_83 qb_51_83 bit_51_83 bitb_51_83 word51_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_83 q_52_83 qb_52_83 bit_52_83 bitb_52_83 word52_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_83 q_53_83 qb_53_83 bit_53_83 bitb_53_83 word53_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_83 q_54_83 qb_54_83 bit_54_83 bitb_54_83 word54_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_83 q_55_83 qb_55_83 bit_55_83 bitb_55_83 word55_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_83 q_56_83 qb_56_83 bit_56_83 bitb_56_83 word56_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_83 q_57_83 qb_57_83 bit_57_83 bitb_57_83 word57_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_83 q_58_83 qb_58_83 bit_58_83 bitb_58_83 word58_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_83 q_59_83 qb_59_83 bit_59_83 bitb_59_83 word59_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_83 q_60_83 qb_60_83 bit_60_83 bitb_60_83 word60_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_83 q_61_83 qb_61_83 bit_61_83 bitb_61_83 word61_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_83 q_62_83 qb_62_83 bit_62_83 bitb_62_83 word62_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_83 q_63_83 qb_63_83 bit_63_83 bitb_63_83 word63_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_83 q_64_83 qb_64_83 bit_64_83 bitb_64_83 word64_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_83 q_65_83 qb_65_83 bit_65_83 bitb_65_83 word65_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_83 q_66_83 qb_66_83 bit_66_83 bitb_66_83 word66_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_83 q_67_83 qb_67_83 bit_67_83 bitb_67_83 word67_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_83 q_68_83 qb_68_83 bit_68_83 bitb_68_83 word68_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_83 q_69_83 qb_69_83 bit_69_83 bitb_69_83 word69_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_83 q_70_83 qb_70_83 bit_70_83 bitb_70_83 word70_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_83 q_71_83 qb_71_83 bit_71_83 bitb_71_83 word71_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_83 q_72_83 qb_72_83 bit_72_83 bitb_72_83 word72_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_83 q_73_83 qb_73_83 bit_73_83 bitb_73_83 word73_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_83 q_74_83 qb_74_83 bit_74_83 bitb_74_83 word74_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_83 q_75_83 qb_75_83 bit_75_83 bitb_75_83 word75_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_83 q_76_83 qb_76_83 bit_76_83 bitb_76_83 word76_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_83 q_77_83 qb_77_83 bit_77_83 bitb_77_83 word77_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_83 q_78_83 qb_78_83 bit_78_83 bitb_78_83 word78_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_83 q_79_83 qb_79_83 bit_79_83 bitb_79_83 word79_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_83 q_80_83 qb_80_83 bit_80_83 bitb_80_83 word80_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_83 q_81_83 qb_81_83 bit_81_83 bitb_81_83 word81_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_83 q_82_83 qb_82_83 bit_82_83 bitb_82_83 word82_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_83 q_83_83 qb_83_83 bit_83_83 bitb_83_83 word83_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_83 q_84_83 qb_84_83 bit_84_83 bitb_84_83 word84_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_83 q_85_83 qb_85_83 bit_85_83 bitb_85_83 word85_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_83 q_86_83 qb_86_83 bit_86_83 bitb_86_83 word86_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_83 q_87_83 qb_87_83 bit_87_83 bitb_87_83 word87_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_83 q_88_83 qb_88_83 bit_88_83 bitb_88_83 word88_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_83 q_89_83 qb_89_83 bit_89_83 bitb_89_83 word89_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_83 q_90_83 qb_90_83 bit_90_83 bitb_90_83 word90_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_83 q_91_83 qb_91_83 bit_91_83 bitb_91_83 word91_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_83 q_92_83 qb_92_83 bit_92_83 bitb_92_83 word92_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_83 q_93_83 qb_93_83 bit_93_83 bitb_93_83 word93_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_83 q_94_83 qb_94_83 bit_94_83 bitb_94_83 word94_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_83 q_95_83 qb_95_83 bit_95_83 bitb_95_83 word95_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_83 q_96_83 qb_96_83 bit_96_83 bitb_96_83 word96_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_83 q_97_83 qb_97_83 bit_97_83 bitb_97_83 word97_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_83 q_98_83 qb_98_83 bit_98_83 bitb_98_83 word98_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_83 q_99_83 qb_99_83 bit_99_83 bitb_99_83 word99_83 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_84 q_0_84 qb_0_84 bit_0_84 bitb_0_84 word0_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_84 q_1_84 qb_1_84 bit_1_84 bitb_1_84 word1_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_84 q_2_84 qb_2_84 bit_2_84 bitb_2_84 word2_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_84 q_3_84 qb_3_84 bit_3_84 bitb_3_84 word3_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_84 q_4_84 qb_4_84 bit_4_84 bitb_4_84 word4_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_84 q_5_84 qb_5_84 bit_5_84 bitb_5_84 word5_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_84 q_6_84 qb_6_84 bit_6_84 bitb_6_84 word6_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_84 q_7_84 qb_7_84 bit_7_84 bitb_7_84 word7_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_84 q_8_84 qb_8_84 bit_8_84 bitb_8_84 word8_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_84 q_9_84 qb_9_84 bit_9_84 bitb_9_84 word9_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_84 q_10_84 qb_10_84 bit_10_84 bitb_10_84 word10_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_84 q_11_84 qb_11_84 bit_11_84 bitb_11_84 word11_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_84 q_12_84 qb_12_84 bit_12_84 bitb_12_84 word12_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_84 q_13_84 qb_13_84 bit_13_84 bitb_13_84 word13_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_84 q_14_84 qb_14_84 bit_14_84 bitb_14_84 word14_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_84 q_15_84 qb_15_84 bit_15_84 bitb_15_84 word15_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_84 q_16_84 qb_16_84 bit_16_84 bitb_16_84 word16_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_84 q_17_84 qb_17_84 bit_17_84 bitb_17_84 word17_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_84 q_18_84 qb_18_84 bit_18_84 bitb_18_84 word18_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_84 q_19_84 qb_19_84 bit_19_84 bitb_19_84 word19_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_84 q_20_84 qb_20_84 bit_20_84 bitb_20_84 word20_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_84 q_21_84 qb_21_84 bit_21_84 bitb_21_84 word21_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_84 q_22_84 qb_22_84 bit_22_84 bitb_22_84 word22_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_84 q_23_84 qb_23_84 bit_23_84 bitb_23_84 word23_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_84 q_24_84 qb_24_84 bit_24_84 bitb_24_84 word24_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_84 q_25_84 qb_25_84 bit_25_84 bitb_25_84 word25_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_84 q_26_84 qb_26_84 bit_26_84 bitb_26_84 word26_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_84 q_27_84 qb_27_84 bit_27_84 bitb_27_84 word27_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_84 q_28_84 qb_28_84 bit_28_84 bitb_28_84 word28_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_84 q_29_84 qb_29_84 bit_29_84 bitb_29_84 word29_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_84 q_30_84 qb_30_84 bit_30_84 bitb_30_84 word30_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_84 q_31_84 qb_31_84 bit_31_84 bitb_31_84 word31_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_84 q_32_84 qb_32_84 bit_32_84 bitb_32_84 word32_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_84 q_33_84 qb_33_84 bit_33_84 bitb_33_84 word33_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_84 q_34_84 qb_34_84 bit_34_84 bitb_34_84 word34_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_84 q_35_84 qb_35_84 bit_35_84 bitb_35_84 word35_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_84 q_36_84 qb_36_84 bit_36_84 bitb_36_84 word36_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_84 q_37_84 qb_37_84 bit_37_84 bitb_37_84 word37_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_84 q_38_84 qb_38_84 bit_38_84 bitb_38_84 word38_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_84 q_39_84 qb_39_84 bit_39_84 bitb_39_84 word39_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_84 q_40_84 qb_40_84 bit_40_84 bitb_40_84 word40_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_84 q_41_84 qb_41_84 bit_41_84 bitb_41_84 word41_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_84 q_42_84 qb_42_84 bit_42_84 bitb_42_84 word42_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_84 q_43_84 qb_43_84 bit_43_84 bitb_43_84 word43_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_84 q_44_84 qb_44_84 bit_44_84 bitb_44_84 word44_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_84 q_45_84 qb_45_84 bit_45_84 bitb_45_84 word45_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_84 q_46_84 qb_46_84 bit_46_84 bitb_46_84 word46_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_84 q_47_84 qb_47_84 bit_47_84 bitb_47_84 word47_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_84 q_48_84 qb_48_84 bit_48_84 bitb_48_84 word48_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_84 q_49_84 qb_49_84 bit_49_84 bitb_49_84 word49_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_84 q_50_84 qb_50_84 bit_50_84 bitb_50_84 word50_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_84 q_51_84 qb_51_84 bit_51_84 bitb_51_84 word51_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_84 q_52_84 qb_52_84 bit_52_84 bitb_52_84 word52_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_84 q_53_84 qb_53_84 bit_53_84 bitb_53_84 word53_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_84 q_54_84 qb_54_84 bit_54_84 bitb_54_84 word54_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_84 q_55_84 qb_55_84 bit_55_84 bitb_55_84 word55_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_84 q_56_84 qb_56_84 bit_56_84 bitb_56_84 word56_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_84 q_57_84 qb_57_84 bit_57_84 bitb_57_84 word57_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_84 q_58_84 qb_58_84 bit_58_84 bitb_58_84 word58_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_84 q_59_84 qb_59_84 bit_59_84 bitb_59_84 word59_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_84 q_60_84 qb_60_84 bit_60_84 bitb_60_84 word60_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_84 q_61_84 qb_61_84 bit_61_84 bitb_61_84 word61_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_84 q_62_84 qb_62_84 bit_62_84 bitb_62_84 word62_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_84 q_63_84 qb_63_84 bit_63_84 bitb_63_84 word63_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_84 q_64_84 qb_64_84 bit_64_84 bitb_64_84 word64_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_84 q_65_84 qb_65_84 bit_65_84 bitb_65_84 word65_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_84 q_66_84 qb_66_84 bit_66_84 bitb_66_84 word66_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_84 q_67_84 qb_67_84 bit_67_84 bitb_67_84 word67_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_84 q_68_84 qb_68_84 bit_68_84 bitb_68_84 word68_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_84 q_69_84 qb_69_84 bit_69_84 bitb_69_84 word69_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_84 q_70_84 qb_70_84 bit_70_84 bitb_70_84 word70_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_84 q_71_84 qb_71_84 bit_71_84 bitb_71_84 word71_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_84 q_72_84 qb_72_84 bit_72_84 bitb_72_84 word72_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_84 q_73_84 qb_73_84 bit_73_84 bitb_73_84 word73_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_84 q_74_84 qb_74_84 bit_74_84 bitb_74_84 word74_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_84 q_75_84 qb_75_84 bit_75_84 bitb_75_84 word75_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_84 q_76_84 qb_76_84 bit_76_84 bitb_76_84 word76_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_84 q_77_84 qb_77_84 bit_77_84 bitb_77_84 word77_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_84 q_78_84 qb_78_84 bit_78_84 bitb_78_84 word78_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_84 q_79_84 qb_79_84 bit_79_84 bitb_79_84 word79_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_84 q_80_84 qb_80_84 bit_80_84 bitb_80_84 word80_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_84 q_81_84 qb_81_84 bit_81_84 bitb_81_84 word81_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_84 q_82_84 qb_82_84 bit_82_84 bitb_82_84 word82_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_84 q_83_84 qb_83_84 bit_83_84 bitb_83_84 word83_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_84 q_84_84 qb_84_84 bit_84_84 bitb_84_84 word84_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_84 q_85_84 qb_85_84 bit_85_84 bitb_85_84 word85_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_84 q_86_84 qb_86_84 bit_86_84 bitb_86_84 word86_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_84 q_87_84 qb_87_84 bit_87_84 bitb_87_84 word87_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_84 q_88_84 qb_88_84 bit_88_84 bitb_88_84 word88_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_84 q_89_84 qb_89_84 bit_89_84 bitb_89_84 word89_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_84 q_90_84 qb_90_84 bit_90_84 bitb_90_84 word90_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_84 q_91_84 qb_91_84 bit_91_84 bitb_91_84 word91_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_84 q_92_84 qb_92_84 bit_92_84 bitb_92_84 word92_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_84 q_93_84 qb_93_84 bit_93_84 bitb_93_84 word93_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_84 q_94_84 qb_94_84 bit_94_84 bitb_94_84 word94_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_84 q_95_84 qb_95_84 bit_95_84 bitb_95_84 word95_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_84 q_96_84 qb_96_84 bit_96_84 bitb_96_84 word96_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_84 q_97_84 qb_97_84 bit_97_84 bitb_97_84 word97_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_84 q_98_84 qb_98_84 bit_98_84 bitb_98_84 word98_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_84 q_99_84 qb_99_84 bit_99_84 bitb_99_84 word99_84 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_85 q_0_85 qb_0_85 bit_0_85 bitb_0_85 word0_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_85 q_1_85 qb_1_85 bit_1_85 bitb_1_85 word1_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_85 q_2_85 qb_2_85 bit_2_85 bitb_2_85 word2_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_85 q_3_85 qb_3_85 bit_3_85 bitb_3_85 word3_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_85 q_4_85 qb_4_85 bit_4_85 bitb_4_85 word4_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_85 q_5_85 qb_5_85 bit_5_85 bitb_5_85 word5_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_85 q_6_85 qb_6_85 bit_6_85 bitb_6_85 word6_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_85 q_7_85 qb_7_85 bit_7_85 bitb_7_85 word7_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_85 q_8_85 qb_8_85 bit_8_85 bitb_8_85 word8_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_85 q_9_85 qb_9_85 bit_9_85 bitb_9_85 word9_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_85 q_10_85 qb_10_85 bit_10_85 bitb_10_85 word10_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_85 q_11_85 qb_11_85 bit_11_85 bitb_11_85 word11_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_85 q_12_85 qb_12_85 bit_12_85 bitb_12_85 word12_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_85 q_13_85 qb_13_85 bit_13_85 bitb_13_85 word13_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_85 q_14_85 qb_14_85 bit_14_85 bitb_14_85 word14_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_85 q_15_85 qb_15_85 bit_15_85 bitb_15_85 word15_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_85 q_16_85 qb_16_85 bit_16_85 bitb_16_85 word16_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_85 q_17_85 qb_17_85 bit_17_85 bitb_17_85 word17_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_85 q_18_85 qb_18_85 bit_18_85 bitb_18_85 word18_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_85 q_19_85 qb_19_85 bit_19_85 bitb_19_85 word19_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_85 q_20_85 qb_20_85 bit_20_85 bitb_20_85 word20_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_85 q_21_85 qb_21_85 bit_21_85 bitb_21_85 word21_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_85 q_22_85 qb_22_85 bit_22_85 bitb_22_85 word22_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_85 q_23_85 qb_23_85 bit_23_85 bitb_23_85 word23_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_85 q_24_85 qb_24_85 bit_24_85 bitb_24_85 word24_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_85 q_25_85 qb_25_85 bit_25_85 bitb_25_85 word25_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_85 q_26_85 qb_26_85 bit_26_85 bitb_26_85 word26_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_85 q_27_85 qb_27_85 bit_27_85 bitb_27_85 word27_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_85 q_28_85 qb_28_85 bit_28_85 bitb_28_85 word28_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_85 q_29_85 qb_29_85 bit_29_85 bitb_29_85 word29_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_85 q_30_85 qb_30_85 bit_30_85 bitb_30_85 word30_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_85 q_31_85 qb_31_85 bit_31_85 bitb_31_85 word31_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_85 q_32_85 qb_32_85 bit_32_85 bitb_32_85 word32_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_85 q_33_85 qb_33_85 bit_33_85 bitb_33_85 word33_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_85 q_34_85 qb_34_85 bit_34_85 bitb_34_85 word34_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_85 q_35_85 qb_35_85 bit_35_85 bitb_35_85 word35_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_85 q_36_85 qb_36_85 bit_36_85 bitb_36_85 word36_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_85 q_37_85 qb_37_85 bit_37_85 bitb_37_85 word37_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_85 q_38_85 qb_38_85 bit_38_85 bitb_38_85 word38_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_85 q_39_85 qb_39_85 bit_39_85 bitb_39_85 word39_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_85 q_40_85 qb_40_85 bit_40_85 bitb_40_85 word40_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_85 q_41_85 qb_41_85 bit_41_85 bitb_41_85 word41_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_85 q_42_85 qb_42_85 bit_42_85 bitb_42_85 word42_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_85 q_43_85 qb_43_85 bit_43_85 bitb_43_85 word43_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_85 q_44_85 qb_44_85 bit_44_85 bitb_44_85 word44_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_85 q_45_85 qb_45_85 bit_45_85 bitb_45_85 word45_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_85 q_46_85 qb_46_85 bit_46_85 bitb_46_85 word46_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_85 q_47_85 qb_47_85 bit_47_85 bitb_47_85 word47_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_85 q_48_85 qb_48_85 bit_48_85 bitb_48_85 word48_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_85 q_49_85 qb_49_85 bit_49_85 bitb_49_85 word49_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_85 q_50_85 qb_50_85 bit_50_85 bitb_50_85 word50_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_85 q_51_85 qb_51_85 bit_51_85 bitb_51_85 word51_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_85 q_52_85 qb_52_85 bit_52_85 bitb_52_85 word52_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_85 q_53_85 qb_53_85 bit_53_85 bitb_53_85 word53_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_85 q_54_85 qb_54_85 bit_54_85 bitb_54_85 word54_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_85 q_55_85 qb_55_85 bit_55_85 bitb_55_85 word55_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_85 q_56_85 qb_56_85 bit_56_85 bitb_56_85 word56_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_85 q_57_85 qb_57_85 bit_57_85 bitb_57_85 word57_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_85 q_58_85 qb_58_85 bit_58_85 bitb_58_85 word58_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_85 q_59_85 qb_59_85 bit_59_85 bitb_59_85 word59_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_85 q_60_85 qb_60_85 bit_60_85 bitb_60_85 word60_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_85 q_61_85 qb_61_85 bit_61_85 bitb_61_85 word61_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_85 q_62_85 qb_62_85 bit_62_85 bitb_62_85 word62_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_85 q_63_85 qb_63_85 bit_63_85 bitb_63_85 word63_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_85 q_64_85 qb_64_85 bit_64_85 bitb_64_85 word64_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_85 q_65_85 qb_65_85 bit_65_85 bitb_65_85 word65_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_85 q_66_85 qb_66_85 bit_66_85 bitb_66_85 word66_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_85 q_67_85 qb_67_85 bit_67_85 bitb_67_85 word67_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_85 q_68_85 qb_68_85 bit_68_85 bitb_68_85 word68_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_85 q_69_85 qb_69_85 bit_69_85 bitb_69_85 word69_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_85 q_70_85 qb_70_85 bit_70_85 bitb_70_85 word70_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_85 q_71_85 qb_71_85 bit_71_85 bitb_71_85 word71_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_85 q_72_85 qb_72_85 bit_72_85 bitb_72_85 word72_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_85 q_73_85 qb_73_85 bit_73_85 bitb_73_85 word73_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_85 q_74_85 qb_74_85 bit_74_85 bitb_74_85 word74_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_85 q_75_85 qb_75_85 bit_75_85 bitb_75_85 word75_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_85 q_76_85 qb_76_85 bit_76_85 bitb_76_85 word76_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_85 q_77_85 qb_77_85 bit_77_85 bitb_77_85 word77_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_85 q_78_85 qb_78_85 bit_78_85 bitb_78_85 word78_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_85 q_79_85 qb_79_85 bit_79_85 bitb_79_85 word79_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_85 q_80_85 qb_80_85 bit_80_85 bitb_80_85 word80_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_85 q_81_85 qb_81_85 bit_81_85 bitb_81_85 word81_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_85 q_82_85 qb_82_85 bit_82_85 bitb_82_85 word82_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_85 q_83_85 qb_83_85 bit_83_85 bitb_83_85 word83_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_85 q_84_85 qb_84_85 bit_84_85 bitb_84_85 word84_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_85 q_85_85 qb_85_85 bit_85_85 bitb_85_85 word85_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_85 q_86_85 qb_86_85 bit_86_85 bitb_86_85 word86_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_85 q_87_85 qb_87_85 bit_87_85 bitb_87_85 word87_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_85 q_88_85 qb_88_85 bit_88_85 bitb_88_85 word88_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_85 q_89_85 qb_89_85 bit_89_85 bitb_89_85 word89_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_85 q_90_85 qb_90_85 bit_90_85 bitb_90_85 word90_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_85 q_91_85 qb_91_85 bit_91_85 bitb_91_85 word91_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_85 q_92_85 qb_92_85 bit_92_85 bitb_92_85 word92_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_85 q_93_85 qb_93_85 bit_93_85 bitb_93_85 word93_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_85 q_94_85 qb_94_85 bit_94_85 bitb_94_85 word94_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_85 q_95_85 qb_95_85 bit_95_85 bitb_95_85 word95_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_85 q_96_85 qb_96_85 bit_96_85 bitb_96_85 word96_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_85 q_97_85 qb_97_85 bit_97_85 bitb_97_85 word97_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_85 q_98_85 qb_98_85 bit_98_85 bitb_98_85 word98_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_85 q_99_85 qb_99_85 bit_99_85 bitb_99_85 word99_85 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_86 q_0_86 qb_0_86 bit_0_86 bitb_0_86 word0_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_86 q_1_86 qb_1_86 bit_1_86 bitb_1_86 word1_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_86 q_2_86 qb_2_86 bit_2_86 bitb_2_86 word2_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_86 q_3_86 qb_3_86 bit_3_86 bitb_3_86 word3_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_86 q_4_86 qb_4_86 bit_4_86 bitb_4_86 word4_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_86 q_5_86 qb_5_86 bit_5_86 bitb_5_86 word5_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_86 q_6_86 qb_6_86 bit_6_86 bitb_6_86 word6_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_86 q_7_86 qb_7_86 bit_7_86 bitb_7_86 word7_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_86 q_8_86 qb_8_86 bit_8_86 bitb_8_86 word8_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_86 q_9_86 qb_9_86 bit_9_86 bitb_9_86 word9_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_86 q_10_86 qb_10_86 bit_10_86 bitb_10_86 word10_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_86 q_11_86 qb_11_86 bit_11_86 bitb_11_86 word11_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_86 q_12_86 qb_12_86 bit_12_86 bitb_12_86 word12_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_86 q_13_86 qb_13_86 bit_13_86 bitb_13_86 word13_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_86 q_14_86 qb_14_86 bit_14_86 bitb_14_86 word14_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_86 q_15_86 qb_15_86 bit_15_86 bitb_15_86 word15_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_86 q_16_86 qb_16_86 bit_16_86 bitb_16_86 word16_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_86 q_17_86 qb_17_86 bit_17_86 bitb_17_86 word17_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_86 q_18_86 qb_18_86 bit_18_86 bitb_18_86 word18_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_86 q_19_86 qb_19_86 bit_19_86 bitb_19_86 word19_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_86 q_20_86 qb_20_86 bit_20_86 bitb_20_86 word20_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_86 q_21_86 qb_21_86 bit_21_86 bitb_21_86 word21_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_86 q_22_86 qb_22_86 bit_22_86 bitb_22_86 word22_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_86 q_23_86 qb_23_86 bit_23_86 bitb_23_86 word23_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_86 q_24_86 qb_24_86 bit_24_86 bitb_24_86 word24_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_86 q_25_86 qb_25_86 bit_25_86 bitb_25_86 word25_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_86 q_26_86 qb_26_86 bit_26_86 bitb_26_86 word26_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_86 q_27_86 qb_27_86 bit_27_86 bitb_27_86 word27_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_86 q_28_86 qb_28_86 bit_28_86 bitb_28_86 word28_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_86 q_29_86 qb_29_86 bit_29_86 bitb_29_86 word29_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_86 q_30_86 qb_30_86 bit_30_86 bitb_30_86 word30_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_86 q_31_86 qb_31_86 bit_31_86 bitb_31_86 word31_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_86 q_32_86 qb_32_86 bit_32_86 bitb_32_86 word32_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_86 q_33_86 qb_33_86 bit_33_86 bitb_33_86 word33_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_86 q_34_86 qb_34_86 bit_34_86 bitb_34_86 word34_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_86 q_35_86 qb_35_86 bit_35_86 bitb_35_86 word35_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_86 q_36_86 qb_36_86 bit_36_86 bitb_36_86 word36_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_86 q_37_86 qb_37_86 bit_37_86 bitb_37_86 word37_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_86 q_38_86 qb_38_86 bit_38_86 bitb_38_86 word38_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_86 q_39_86 qb_39_86 bit_39_86 bitb_39_86 word39_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_86 q_40_86 qb_40_86 bit_40_86 bitb_40_86 word40_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_86 q_41_86 qb_41_86 bit_41_86 bitb_41_86 word41_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_86 q_42_86 qb_42_86 bit_42_86 bitb_42_86 word42_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_86 q_43_86 qb_43_86 bit_43_86 bitb_43_86 word43_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_86 q_44_86 qb_44_86 bit_44_86 bitb_44_86 word44_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_86 q_45_86 qb_45_86 bit_45_86 bitb_45_86 word45_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_86 q_46_86 qb_46_86 bit_46_86 bitb_46_86 word46_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_86 q_47_86 qb_47_86 bit_47_86 bitb_47_86 word47_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_86 q_48_86 qb_48_86 bit_48_86 bitb_48_86 word48_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_86 q_49_86 qb_49_86 bit_49_86 bitb_49_86 word49_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_86 q_50_86 qb_50_86 bit_50_86 bitb_50_86 word50_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_86 q_51_86 qb_51_86 bit_51_86 bitb_51_86 word51_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_86 q_52_86 qb_52_86 bit_52_86 bitb_52_86 word52_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_86 q_53_86 qb_53_86 bit_53_86 bitb_53_86 word53_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_86 q_54_86 qb_54_86 bit_54_86 bitb_54_86 word54_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_86 q_55_86 qb_55_86 bit_55_86 bitb_55_86 word55_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_86 q_56_86 qb_56_86 bit_56_86 bitb_56_86 word56_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_86 q_57_86 qb_57_86 bit_57_86 bitb_57_86 word57_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_86 q_58_86 qb_58_86 bit_58_86 bitb_58_86 word58_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_86 q_59_86 qb_59_86 bit_59_86 bitb_59_86 word59_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_86 q_60_86 qb_60_86 bit_60_86 bitb_60_86 word60_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_86 q_61_86 qb_61_86 bit_61_86 bitb_61_86 word61_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_86 q_62_86 qb_62_86 bit_62_86 bitb_62_86 word62_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_86 q_63_86 qb_63_86 bit_63_86 bitb_63_86 word63_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_86 q_64_86 qb_64_86 bit_64_86 bitb_64_86 word64_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_86 q_65_86 qb_65_86 bit_65_86 bitb_65_86 word65_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_86 q_66_86 qb_66_86 bit_66_86 bitb_66_86 word66_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_86 q_67_86 qb_67_86 bit_67_86 bitb_67_86 word67_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_86 q_68_86 qb_68_86 bit_68_86 bitb_68_86 word68_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_86 q_69_86 qb_69_86 bit_69_86 bitb_69_86 word69_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_86 q_70_86 qb_70_86 bit_70_86 bitb_70_86 word70_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_86 q_71_86 qb_71_86 bit_71_86 bitb_71_86 word71_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_86 q_72_86 qb_72_86 bit_72_86 bitb_72_86 word72_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_86 q_73_86 qb_73_86 bit_73_86 bitb_73_86 word73_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_86 q_74_86 qb_74_86 bit_74_86 bitb_74_86 word74_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_86 q_75_86 qb_75_86 bit_75_86 bitb_75_86 word75_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_86 q_76_86 qb_76_86 bit_76_86 bitb_76_86 word76_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_86 q_77_86 qb_77_86 bit_77_86 bitb_77_86 word77_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_86 q_78_86 qb_78_86 bit_78_86 bitb_78_86 word78_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_86 q_79_86 qb_79_86 bit_79_86 bitb_79_86 word79_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_86 q_80_86 qb_80_86 bit_80_86 bitb_80_86 word80_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_86 q_81_86 qb_81_86 bit_81_86 bitb_81_86 word81_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_86 q_82_86 qb_82_86 bit_82_86 bitb_82_86 word82_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_86 q_83_86 qb_83_86 bit_83_86 bitb_83_86 word83_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_86 q_84_86 qb_84_86 bit_84_86 bitb_84_86 word84_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_86 q_85_86 qb_85_86 bit_85_86 bitb_85_86 word85_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_86 q_86_86 qb_86_86 bit_86_86 bitb_86_86 word86_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_86 q_87_86 qb_87_86 bit_87_86 bitb_87_86 word87_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_86 q_88_86 qb_88_86 bit_88_86 bitb_88_86 word88_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_86 q_89_86 qb_89_86 bit_89_86 bitb_89_86 word89_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_86 q_90_86 qb_90_86 bit_90_86 bitb_90_86 word90_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_86 q_91_86 qb_91_86 bit_91_86 bitb_91_86 word91_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_86 q_92_86 qb_92_86 bit_92_86 bitb_92_86 word92_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_86 q_93_86 qb_93_86 bit_93_86 bitb_93_86 word93_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_86 q_94_86 qb_94_86 bit_94_86 bitb_94_86 word94_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_86 q_95_86 qb_95_86 bit_95_86 bitb_95_86 word95_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_86 q_96_86 qb_96_86 bit_96_86 bitb_96_86 word96_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_86 q_97_86 qb_97_86 bit_97_86 bitb_97_86 word97_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_86 q_98_86 qb_98_86 bit_98_86 bitb_98_86 word98_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_86 q_99_86 qb_99_86 bit_99_86 bitb_99_86 word99_86 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_87 q_0_87 qb_0_87 bit_0_87 bitb_0_87 word0_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_87 q_1_87 qb_1_87 bit_1_87 bitb_1_87 word1_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_87 q_2_87 qb_2_87 bit_2_87 bitb_2_87 word2_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_87 q_3_87 qb_3_87 bit_3_87 bitb_3_87 word3_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_87 q_4_87 qb_4_87 bit_4_87 bitb_4_87 word4_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_87 q_5_87 qb_5_87 bit_5_87 bitb_5_87 word5_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_87 q_6_87 qb_6_87 bit_6_87 bitb_6_87 word6_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_87 q_7_87 qb_7_87 bit_7_87 bitb_7_87 word7_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_87 q_8_87 qb_8_87 bit_8_87 bitb_8_87 word8_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_87 q_9_87 qb_9_87 bit_9_87 bitb_9_87 word9_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_87 q_10_87 qb_10_87 bit_10_87 bitb_10_87 word10_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_87 q_11_87 qb_11_87 bit_11_87 bitb_11_87 word11_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_87 q_12_87 qb_12_87 bit_12_87 bitb_12_87 word12_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_87 q_13_87 qb_13_87 bit_13_87 bitb_13_87 word13_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_87 q_14_87 qb_14_87 bit_14_87 bitb_14_87 word14_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_87 q_15_87 qb_15_87 bit_15_87 bitb_15_87 word15_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_87 q_16_87 qb_16_87 bit_16_87 bitb_16_87 word16_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_87 q_17_87 qb_17_87 bit_17_87 bitb_17_87 word17_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_87 q_18_87 qb_18_87 bit_18_87 bitb_18_87 word18_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_87 q_19_87 qb_19_87 bit_19_87 bitb_19_87 word19_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_87 q_20_87 qb_20_87 bit_20_87 bitb_20_87 word20_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_87 q_21_87 qb_21_87 bit_21_87 bitb_21_87 word21_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_87 q_22_87 qb_22_87 bit_22_87 bitb_22_87 word22_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_87 q_23_87 qb_23_87 bit_23_87 bitb_23_87 word23_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_87 q_24_87 qb_24_87 bit_24_87 bitb_24_87 word24_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_87 q_25_87 qb_25_87 bit_25_87 bitb_25_87 word25_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_87 q_26_87 qb_26_87 bit_26_87 bitb_26_87 word26_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_87 q_27_87 qb_27_87 bit_27_87 bitb_27_87 word27_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_87 q_28_87 qb_28_87 bit_28_87 bitb_28_87 word28_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_87 q_29_87 qb_29_87 bit_29_87 bitb_29_87 word29_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_87 q_30_87 qb_30_87 bit_30_87 bitb_30_87 word30_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_87 q_31_87 qb_31_87 bit_31_87 bitb_31_87 word31_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_87 q_32_87 qb_32_87 bit_32_87 bitb_32_87 word32_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_87 q_33_87 qb_33_87 bit_33_87 bitb_33_87 word33_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_87 q_34_87 qb_34_87 bit_34_87 bitb_34_87 word34_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_87 q_35_87 qb_35_87 bit_35_87 bitb_35_87 word35_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_87 q_36_87 qb_36_87 bit_36_87 bitb_36_87 word36_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_87 q_37_87 qb_37_87 bit_37_87 bitb_37_87 word37_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_87 q_38_87 qb_38_87 bit_38_87 bitb_38_87 word38_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_87 q_39_87 qb_39_87 bit_39_87 bitb_39_87 word39_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_87 q_40_87 qb_40_87 bit_40_87 bitb_40_87 word40_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_87 q_41_87 qb_41_87 bit_41_87 bitb_41_87 word41_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_87 q_42_87 qb_42_87 bit_42_87 bitb_42_87 word42_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_87 q_43_87 qb_43_87 bit_43_87 bitb_43_87 word43_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_87 q_44_87 qb_44_87 bit_44_87 bitb_44_87 word44_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_87 q_45_87 qb_45_87 bit_45_87 bitb_45_87 word45_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_87 q_46_87 qb_46_87 bit_46_87 bitb_46_87 word46_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_87 q_47_87 qb_47_87 bit_47_87 bitb_47_87 word47_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_87 q_48_87 qb_48_87 bit_48_87 bitb_48_87 word48_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_87 q_49_87 qb_49_87 bit_49_87 bitb_49_87 word49_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_87 q_50_87 qb_50_87 bit_50_87 bitb_50_87 word50_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_87 q_51_87 qb_51_87 bit_51_87 bitb_51_87 word51_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_87 q_52_87 qb_52_87 bit_52_87 bitb_52_87 word52_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_87 q_53_87 qb_53_87 bit_53_87 bitb_53_87 word53_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_87 q_54_87 qb_54_87 bit_54_87 bitb_54_87 word54_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_87 q_55_87 qb_55_87 bit_55_87 bitb_55_87 word55_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_87 q_56_87 qb_56_87 bit_56_87 bitb_56_87 word56_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_87 q_57_87 qb_57_87 bit_57_87 bitb_57_87 word57_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_87 q_58_87 qb_58_87 bit_58_87 bitb_58_87 word58_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_87 q_59_87 qb_59_87 bit_59_87 bitb_59_87 word59_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_87 q_60_87 qb_60_87 bit_60_87 bitb_60_87 word60_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_87 q_61_87 qb_61_87 bit_61_87 bitb_61_87 word61_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_87 q_62_87 qb_62_87 bit_62_87 bitb_62_87 word62_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_87 q_63_87 qb_63_87 bit_63_87 bitb_63_87 word63_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_87 q_64_87 qb_64_87 bit_64_87 bitb_64_87 word64_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_87 q_65_87 qb_65_87 bit_65_87 bitb_65_87 word65_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_87 q_66_87 qb_66_87 bit_66_87 bitb_66_87 word66_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_87 q_67_87 qb_67_87 bit_67_87 bitb_67_87 word67_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_87 q_68_87 qb_68_87 bit_68_87 bitb_68_87 word68_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_87 q_69_87 qb_69_87 bit_69_87 bitb_69_87 word69_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_87 q_70_87 qb_70_87 bit_70_87 bitb_70_87 word70_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_87 q_71_87 qb_71_87 bit_71_87 bitb_71_87 word71_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_87 q_72_87 qb_72_87 bit_72_87 bitb_72_87 word72_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_87 q_73_87 qb_73_87 bit_73_87 bitb_73_87 word73_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_87 q_74_87 qb_74_87 bit_74_87 bitb_74_87 word74_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_87 q_75_87 qb_75_87 bit_75_87 bitb_75_87 word75_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_87 q_76_87 qb_76_87 bit_76_87 bitb_76_87 word76_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_87 q_77_87 qb_77_87 bit_77_87 bitb_77_87 word77_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_87 q_78_87 qb_78_87 bit_78_87 bitb_78_87 word78_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_87 q_79_87 qb_79_87 bit_79_87 bitb_79_87 word79_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_87 q_80_87 qb_80_87 bit_80_87 bitb_80_87 word80_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_87 q_81_87 qb_81_87 bit_81_87 bitb_81_87 word81_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_87 q_82_87 qb_82_87 bit_82_87 bitb_82_87 word82_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_87 q_83_87 qb_83_87 bit_83_87 bitb_83_87 word83_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_87 q_84_87 qb_84_87 bit_84_87 bitb_84_87 word84_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_87 q_85_87 qb_85_87 bit_85_87 bitb_85_87 word85_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_87 q_86_87 qb_86_87 bit_86_87 bitb_86_87 word86_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_87 q_87_87 qb_87_87 bit_87_87 bitb_87_87 word87_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_87 q_88_87 qb_88_87 bit_88_87 bitb_88_87 word88_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_87 q_89_87 qb_89_87 bit_89_87 bitb_89_87 word89_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_87 q_90_87 qb_90_87 bit_90_87 bitb_90_87 word90_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_87 q_91_87 qb_91_87 bit_91_87 bitb_91_87 word91_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_87 q_92_87 qb_92_87 bit_92_87 bitb_92_87 word92_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_87 q_93_87 qb_93_87 bit_93_87 bitb_93_87 word93_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_87 q_94_87 qb_94_87 bit_94_87 bitb_94_87 word94_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_87 q_95_87 qb_95_87 bit_95_87 bitb_95_87 word95_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_87 q_96_87 qb_96_87 bit_96_87 bitb_96_87 word96_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_87 q_97_87 qb_97_87 bit_97_87 bitb_97_87 word97_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_87 q_98_87 qb_98_87 bit_98_87 bitb_98_87 word98_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_87 q_99_87 qb_99_87 bit_99_87 bitb_99_87 word99_87 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_88 q_0_88 qb_0_88 bit_0_88 bitb_0_88 word0_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_88 q_1_88 qb_1_88 bit_1_88 bitb_1_88 word1_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_88 q_2_88 qb_2_88 bit_2_88 bitb_2_88 word2_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_88 q_3_88 qb_3_88 bit_3_88 bitb_3_88 word3_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_88 q_4_88 qb_4_88 bit_4_88 bitb_4_88 word4_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_88 q_5_88 qb_5_88 bit_5_88 bitb_5_88 word5_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_88 q_6_88 qb_6_88 bit_6_88 bitb_6_88 word6_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_88 q_7_88 qb_7_88 bit_7_88 bitb_7_88 word7_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_88 q_8_88 qb_8_88 bit_8_88 bitb_8_88 word8_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_88 q_9_88 qb_9_88 bit_9_88 bitb_9_88 word9_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_88 q_10_88 qb_10_88 bit_10_88 bitb_10_88 word10_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_88 q_11_88 qb_11_88 bit_11_88 bitb_11_88 word11_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_88 q_12_88 qb_12_88 bit_12_88 bitb_12_88 word12_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_88 q_13_88 qb_13_88 bit_13_88 bitb_13_88 word13_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_88 q_14_88 qb_14_88 bit_14_88 bitb_14_88 word14_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_88 q_15_88 qb_15_88 bit_15_88 bitb_15_88 word15_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_88 q_16_88 qb_16_88 bit_16_88 bitb_16_88 word16_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_88 q_17_88 qb_17_88 bit_17_88 bitb_17_88 word17_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_88 q_18_88 qb_18_88 bit_18_88 bitb_18_88 word18_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_88 q_19_88 qb_19_88 bit_19_88 bitb_19_88 word19_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_88 q_20_88 qb_20_88 bit_20_88 bitb_20_88 word20_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_88 q_21_88 qb_21_88 bit_21_88 bitb_21_88 word21_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_88 q_22_88 qb_22_88 bit_22_88 bitb_22_88 word22_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_88 q_23_88 qb_23_88 bit_23_88 bitb_23_88 word23_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_88 q_24_88 qb_24_88 bit_24_88 bitb_24_88 word24_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_88 q_25_88 qb_25_88 bit_25_88 bitb_25_88 word25_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_88 q_26_88 qb_26_88 bit_26_88 bitb_26_88 word26_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_88 q_27_88 qb_27_88 bit_27_88 bitb_27_88 word27_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_88 q_28_88 qb_28_88 bit_28_88 bitb_28_88 word28_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_88 q_29_88 qb_29_88 bit_29_88 bitb_29_88 word29_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_88 q_30_88 qb_30_88 bit_30_88 bitb_30_88 word30_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_88 q_31_88 qb_31_88 bit_31_88 bitb_31_88 word31_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_88 q_32_88 qb_32_88 bit_32_88 bitb_32_88 word32_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_88 q_33_88 qb_33_88 bit_33_88 bitb_33_88 word33_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_88 q_34_88 qb_34_88 bit_34_88 bitb_34_88 word34_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_88 q_35_88 qb_35_88 bit_35_88 bitb_35_88 word35_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_88 q_36_88 qb_36_88 bit_36_88 bitb_36_88 word36_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_88 q_37_88 qb_37_88 bit_37_88 bitb_37_88 word37_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_88 q_38_88 qb_38_88 bit_38_88 bitb_38_88 word38_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_88 q_39_88 qb_39_88 bit_39_88 bitb_39_88 word39_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_88 q_40_88 qb_40_88 bit_40_88 bitb_40_88 word40_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_88 q_41_88 qb_41_88 bit_41_88 bitb_41_88 word41_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_88 q_42_88 qb_42_88 bit_42_88 bitb_42_88 word42_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_88 q_43_88 qb_43_88 bit_43_88 bitb_43_88 word43_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_88 q_44_88 qb_44_88 bit_44_88 bitb_44_88 word44_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_88 q_45_88 qb_45_88 bit_45_88 bitb_45_88 word45_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_88 q_46_88 qb_46_88 bit_46_88 bitb_46_88 word46_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_88 q_47_88 qb_47_88 bit_47_88 bitb_47_88 word47_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_88 q_48_88 qb_48_88 bit_48_88 bitb_48_88 word48_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_88 q_49_88 qb_49_88 bit_49_88 bitb_49_88 word49_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_88 q_50_88 qb_50_88 bit_50_88 bitb_50_88 word50_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_88 q_51_88 qb_51_88 bit_51_88 bitb_51_88 word51_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_88 q_52_88 qb_52_88 bit_52_88 bitb_52_88 word52_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_88 q_53_88 qb_53_88 bit_53_88 bitb_53_88 word53_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_88 q_54_88 qb_54_88 bit_54_88 bitb_54_88 word54_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_88 q_55_88 qb_55_88 bit_55_88 bitb_55_88 word55_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_88 q_56_88 qb_56_88 bit_56_88 bitb_56_88 word56_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_88 q_57_88 qb_57_88 bit_57_88 bitb_57_88 word57_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_88 q_58_88 qb_58_88 bit_58_88 bitb_58_88 word58_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_88 q_59_88 qb_59_88 bit_59_88 bitb_59_88 word59_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_88 q_60_88 qb_60_88 bit_60_88 bitb_60_88 word60_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_88 q_61_88 qb_61_88 bit_61_88 bitb_61_88 word61_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_88 q_62_88 qb_62_88 bit_62_88 bitb_62_88 word62_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_88 q_63_88 qb_63_88 bit_63_88 bitb_63_88 word63_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_88 q_64_88 qb_64_88 bit_64_88 bitb_64_88 word64_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_88 q_65_88 qb_65_88 bit_65_88 bitb_65_88 word65_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_88 q_66_88 qb_66_88 bit_66_88 bitb_66_88 word66_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_88 q_67_88 qb_67_88 bit_67_88 bitb_67_88 word67_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_88 q_68_88 qb_68_88 bit_68_88 bitb_68_88 word68_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_88 q_69_88 qb_69_88 bit_69_88 bitb_69_88 word69_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_88 q_70_88 qb_70_88 bit_70_88 bitb_70_88 word70_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_88 q_71_88 qb_71_88 bit_71_88 bitb_71_88 word71_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_88 q_72_88 qb_72_88 bit_72_88 bitb_72_88 word72_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_88 q_73_88 qb_73_88 bit_73_88 bitb_73_88 word73_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_88 q_74_88 qb_74_88 bit_74_88 bitb_74_88 word74_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_88 q_75_88 qb_75_88 bit_75_88 bitb_75_88 word75_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_88 q_76_88 qb_76_88 bit_76_88 bitb_76_88 word76_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_88 q_77_88 qb_77_88 bit_77_88 bitb_77_88 word77_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_88 q_78_88 qb_78_88 bit_78_88 bitb_78_88 word78_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_88 q_79_88 qb_79_88 bit_79_88 bitb_79_88 word79_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_88 q_80_88 qb_80_88 bit_80_88 bitb_80_88 word80_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_88 q_81_88 qb_81_88 bit_81_88 bitb_81_88 word81_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_88 q_82_88 qb_82_88 bit_82_88 bitb_82_88 word82_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_88 q_83_88 qb_83_88 bit_83_88 bitb_83_88 word83_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_88 q_84_88 qb_84_88 bit_84_88 bitb_84_88 word84_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_88 q_85_88 qb_85_88 bit_85_88 bitb_85_88 word85_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_88 q_86_88 qb_86_88 bit_86_88 bitb_86_88 word86_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_88 q_87_88 qb_87_88 bit_87_88 bitb_87_88 word87_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_88 q_88_88 qb_88_88 bit_88_88 bitb_88_88 word88_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_88 q_89_88 qb_89_88 bit_89_88 bitb_89_88 word89_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_88 q_90_88 qb_90_88 bit_90_88 bitb_90_88 word90_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_88 q_91_88 qb_91_88 bit_91_88 bitb_91_88 word91_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_88 q_92_88 qb_92_88 bit_92_88 bitb_92_88 word92_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_88 q_93_88 qb_93_88 bit_93_88 bitb_93_88 word93_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_88 q_94_88 qb_94_88 bit_94_88 bitb_94_88 word94_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_88 q_95_88 qb_95_88 bit_95_88 bitb_95_88 word95_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_88 q_96_88 qb_96_88 bit_96_88 bitb_96_88 word96_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_88 q_97_88 qb_97_88 bit_97_88 bitb_97_88 word97_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_88 q_98_88 qb_98_88 bit_98_88 bitb_98_88 word98_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_88 q_99_88 qb_99_88 bit_99_88 bitb_99_88 word99_88 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_89 q_0_89 qb_0_89 bit_0_89 bitb_0_89 word0_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_89 q_1_89 qb_1_89 bit_1_89 bitb_1_89 word1_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_89 q_2_89 qb_2_89 bit_2_89 bitb_2_89 word2_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_89 q_3_89 qb_3_89 bit_3_89 bitb_3_89 word3_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_89 q_4_89 qb_4_89 bit_4_89 bitb_4_89 word4_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_89 q_5_89 qb_5_89 bit_5_89 bitb_5_89 word5_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_89 q_6_89 qb_6_89 bit_6_89 bitb_6_89 word6_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_89 q_7_89 qb_7_89 bit_7_89 bitb_7_89 word7_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_89 q_8_89 qb_8_89 bit_8_89 bitb_8_89 word8_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_89 q_9_89 qb_9_89 bit_9_89 bitb_9_89 word9_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_89 q_10_89 qb_10_89 bit_10_89 bitb_10_89 word10_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_89 q_11_89 qb_11_89 bit_11_89 bitb_11_89 word11_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_89 q_12_89 qb_12_89 bit_12_89 bitb_12_89 word12_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_89 q_13_89 qb_13_89 bit_13_89 bitb_13_89 word13_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_89 q_14_89 qb_14_89 bit_14_89 bitb_14_89 word14_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_89 q_15_89 qb_15_89 bit_15_89 bitb_15_89 word15_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_89 q_16_89 qb_16_89 bit_16_89 bitb_16_89 word16_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_89 q_17_89 qb_17_89 bit_17_89 bitb_17_89 word17_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_89 q_18_89 qb_18_89 bit_18_89 bitb_18_89 word18_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_89 q_19_89 qb_19_89 bit_19_89 bitb_19_89 word19_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_89 q_20_89 qb_20_89 bit_20_89 bitb_20_89 word20_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_89 q_21_89 qb_21_89 bit_21_89 bitb_21_89 word21_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_89 q_22_89 qb_22_89 bit_22_89 bitb_22_89 word22_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_89 q_23_89 qb_23_89 bit_23_89 bitb_23_89 word23_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_89 q_24_89 qb_24_89 bit_24_89 bitb_24_89 word24_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_89 q_25_89 qb_25_89 bit_25_89 bitb_25_89 word25_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_89 q_26_89 qb_26_89 bit_26_89 bitb_26_89 word26_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_89 q_27_89 qb_27_89 bit_27_89 bitb_27_89 word27_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_89 q_28_89 qb_28_89 bit_28_89 bitb_28_89 word28_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_89 q_29_89 qb_29_89 bit_29_89 bitb_29_89 word29_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_89 q_30_89 qb_30_89 bit_30_89 bitb_30_89 word30_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_89 q_31_89 qb_31_89 bit_31_89 bitb_31_89 word31_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_89 q_32_89 qb_32_89 bit_32_89 bitb_32_89 word32_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_89 q_33_89 qb_33_89 bit_33_89 bitb_33_89 word33_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_89 q_34_89 qb_34_89 bit_34_89 bitb_34_89 word34_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_89 q_35_89 qb_35_89 bit_35_89 bitb_35_89 word35_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_89 q_36_89 qb_36_89 bit_36_89 bitb_36_89 word36_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_89 q_37_89 qb_37_89 bit_37_89 bitb_37_89 word37_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_89 q_38_89 qb_38_89 bit_38_89 bitb_38_89 word38_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_89 q_39_89 qb_39_89 bit_39_89 bitb_39_89 word39_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_89 q_40_89 qb_40_89 bit_40_89 bitb_40_89 word40_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_89 q_41_89 qb_41_89 bit_41_89 bitb_41_89 word41_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_89 q_42_89 qb_42_89 bit_42_89 bitb_42_89 word42_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_89 q_43_89 qb_43_89 bit_43_89 bitb_43_89 word43_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_89 q_44_89 qb_44_89 bit_44_89 bitb_44_89 word44_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_89 q_45_89 qb_45_89 bit_45_89 bitb_45_89 word45_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_89 q_46_89 qb_46_89 bit_46_89 bitb_46_89 word46_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_89 q_47_89 qb_47_89 bit_47_89 bitb_47_89 word47_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_89 q_48_89 qb_48_89 bit_48_89 bitb_48_89 word48_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_89 q_49_89 qb_49_89 bit_49_89 bitb_49_89 word49_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_89 q_50_89 qb_50_89 bit_50_89 bitb_50_89 word50_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_89 q_51_89 qb_51_89 bit_51_89 bitb_51_89 word51_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_89 q_52_89 qb_52_89 bit_52_89 bitb_52_89 word52_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_89 q_53_89 qb_53_89 bit_53_89 bitb_53_89 word53_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_89 q_54_89 qb_54_89 bit_54_89 bitb_54_89 word54_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_89 q_55_89 qb_55_89 bit_55_89 bitb_55_89 word55_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_89 q_56_89 qb_56_89 bit_56_89 bitb_56_89 word56_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_89 q_57_89 qb_57_89 bit_57_89 bitb_57_89 word57_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_89 q_58_89 qb_58_89 bit_58_89 bitb_58_89 word58_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_89 q_59_89 qb_59_89 bit_59_89 bitb_59_89 word59_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_89 q_60_89 qb_60_89 bit_60_89 bitb_60_89 word60_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_89 q_61_89 qb_61_89 bit_61_89 bitb_61_89 word61_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_89 q_62_89 qb_62_89 bit_62_89 bitb_62_89 word62_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_89 q_63_89 qb_63_89 bit_63_89 bitb_63_89 word63_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_89 q_64_89 qb_64_89 bit_64_89 bitb_64_89 word64_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_89 q_65_89 qb_65_89 bit_65_89 bitb_65_89 word65_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_89 q_66_89 qb_66_89 bit_66_89 bitb_66_89 word66_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_89 q_67_89 qb_67_89 bit_67_89 bitb_67_89 word67_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_89 q_68_89 qb_68_89 bit_68_89 bitb_68_89 word68_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_89 q_69_89 qb_69_89 bit_69_89 bitb_69_89 word69_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_89 q_70_89 qb_70_89 bit_70_89 bitb_70_89 word70_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_89 q_71_89 qb_71_89 bit_71_89 bitb_71_89 word71_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_89 q_72_89 qb_72_89 bit_72_89 bitb_72_89 word72_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_89 q_73_89 qb_73_89 bit_73_89 bitb_73_89 word73_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_89 q_74_89 qb_74_89 bit_74_89 bitb_74_89 word74_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_89 q_75_89 qb_75_89 bit_75_89 bitb_75_89 word75_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_89 q_76_89 qb_76_89 bit_76_89 bitb_76_89 word76_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_89 q_77_89 qb_77_89 bit_77_89 bitb_77_89 word77_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_89 q_78_89 qb_78_89 bit_78_89 bitb_78_89 word78_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_89 q_79_89 qb_79_89 bit_79_89 bitb_79_89 word79_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_89 q_80_89 qb_80_89 bit_80_89 bitb_80_89 word80_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_89 q_81_89 qb_81_89 bit_81_89 bitb_81_89 word81_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_89 q_82_89 qb_82_89 bit_82_89 bitb_82_89 word82_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_89 q_83_89 qb_83_89 bit_83_89 bitb_83_89 word83_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_89 q_84_89 qb_84_89 bit_84_89 bitb_84_89 word84_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_89 q_85_89 qb_85_89 bit_85_89 bitb_85_89 word85_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_89 q_86_89 qb_86_89 bit_86_89 bitb_86_89 word86_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_89 q_87_89 qb_87_89 bit_87_89 bitb_87_89 word87_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_89 q_88_89 qb_88_89 bit_88_89 bitb_88_89 word88_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_89 q_89_89 qb_89_89 bit_89_89 bitb_89_89 word89_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_89 q_90_89 qb_90_89 bit_90_89 bitb_90_89 word90_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_89 q_91_89 qb_91_89 bit_91_89 bitb_91_89 word91_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_89 q_92_89 qb_92_89 bit_92_89 bitb_92_89 word92_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_89 q_93_89 qb_93_89 bit_93_89 bitb_93_89 word93_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_89 q_94_89 qb_94_89 bit_94_89 bitb_94_89 word94_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_89 q_95_89 qb_95_89 bit_95_89 bitb_95_89 word95_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_89 q_96_89 qb_96_89 bit_96_89 bitb_96_89 word96_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_89 q_97_89 qb_97_89 bit_97_89 bitb_97_89 word97_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_89 q_98_89 qb_98_89 bit_98_89 bitb_98_89 word98_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_89 q_99_89 qb_99_89 bit_99_89 bitb_99_89 word99_89 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_90 q_0_90 qb_0_90 bit_0_90 bitb_0_90 word0_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_90 q_1_90 qb_1_90 bit_1_90 bitb_1_90 word1_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_90 q_2_90 qb_2_90 bit_2_90 bitb_2_90 word2_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_90 q_3_90 qb_3_90 bit_3_90 bitb_3_90 word3_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_90 q_4_90 qb_4_90 bit_4_90 bitb_4_90 word4_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_90 q_5_90 qb_5_90 bit_5_90 bitb_5_90 word5_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_90 q_6_90 qb_6_90 bit_6_90 bitb_6_90 word6_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_90 q_7_90 qb_7_90 bit_7_90 bitb_7_90 word7_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_90 q_8_90 qb_8_90 bit_8_90 bitb_8_90 word8_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_90 q_9_90 qb_9_90 bit_9_90 bitb_9_90 word9_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_90 q_10_90 qb_10_90 bit_10_90 bitb_10_90 word10_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_90 q_11_90 qb_11_90 bit_11_90 bitb_11_90 word11_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_90 q_12_90 qb_12_90 bit_12_90 bitb_12_90 word12_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_90 q_13_90 qb_13_90 bit_13_90 bitb_13_90 word13_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_90 q_14_90 qb_14_90 bit_14_90 bitb_14_90 word14_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_90 q_15_90 qb_15_90 bit_15_90 bitb_15_90 word15_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_90 q_16_90 qb_16_90 bit_16_90 bitb_16_90 word16_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_90 q_17_90 qb_17_90 bit_17_90 bitb_17_90 word17_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_90 q_18_90 qb_18_90 bit_18_90 bitb_18_90 word18_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_90 q_19_90 qb_19_90 bit_19_90 bitb_19_90 word19_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_90 q_20_90 qb_20_90 bit_20_90 bitb_20_90 word20_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_90 q_21_90 qb_21_90 bit_21_90 bitb_21_90 word21_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_90 q_22_90 qb_22_90 bit_22_90 bitb_22_90 word22_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_90 q_23_90 qb_23_90 bit_23_90 bitb_23_90 word23_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_90 q_24_90 qb_24_90 bit_24_90 bitb_24_90 word24_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_90 q_25_90 qb_25_90 bit_25_90 bitb_25_90 word25_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_90 q_26_90 qb_26_90 bit_26_90 bitb_26_90 word26_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_90 q_27_90 qb_27_90 bit_27_90 bitb_27_90 word27_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_90 q_28_90 qb_28_90 bit_28_90 bitb_28_90 word28_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_90 q_29_90 qb_29_90 bit_29_90 bitb_29_90 word29_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_90 q_30_90 qb_30_90 bit_30_90 bitb_30_90 word30_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_90 q_31_90 qb_31_90 bit_31_90 bitb_31_90 word31_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_90 q_32_90 qb_32_90 bit_32_90 bitb_32_90 word32_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_90 q_33_90 qb_33_90 bit_33_90 bitb_33_90 word33_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_90 q_34_90 qb_34_90 bit_34_90 bitb_34_90 word34_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_90 q_35_90 qb_35_90 bit_35_90 bitb_35_90 word35_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_90 q_36_90 qb_36_90 bit_36_90 bitb_36_90 word36_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_90 q_37_90 qb_37_90 bit_37_90 bitb_37_90 word37_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_90 q_38_90 qb_38_90 bit_38_90 bitb_38_90 word38_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_90 q_39_90 qb_39_90 bit_39_90 bitb_39_90 word39_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_90 q_40_90 qb_40_90 bit_40_90 bitb_40_90 word40_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_90 q_41_90 qb_41_90 bit_41_90 bitb_41_90 word41_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_90 q_42_90 qb_42_90 bit_42_90 bitb_42_90 word42_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_90 q_43_90 qb_43_90 bit_43_90 bitb_43_90 word43_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_90 q_44_90 qb_44_90 bit_44_90 bitb_44_90 word44_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_90 q_45_90 qb_45_90 bit_45_90 bitb_45_90 word45_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_90 q_46_90 qb_46_90 bit_46_90 bitb_46_90 word46_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_90 q_47_90 qb_47_90 bit_47_90 bitb_47_90 word47_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_90 q_48_90 qb_48_90 bit_48_90 bitb_48_90 word48_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_90 q_49_90 qb_49_90 bit_49_90 bitb_49_90 word49_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_90 q_50_90 qb_50_90 bit_50_90 bitb_50_90 word50_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_90 q_51_90 qb_51_90 bit_51_90 bitb_51_90 word51_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_90 q_52_90 qb_52_90 bit_52_90 bitb_52_90 word52_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_90 q_53_90 qb_53_90 bit_53_90 bitb_53_90 word53_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_90 q_54_90 qb_54_90 bit_54_90 bitb_54_90 word54_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_90 q_55_90 qb_55_90 bit_55_90 bitb_55_90 word55_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_90 q_56_90 qb_56_90 bit_56_90 bitb_56_90 word56_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_90 q_57_90 qb_57_90 bit_57_90 bitb_57_90 word57_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_90 q_58_90 qb_58_90 bit_58_90 bitb_58_90 word58_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_90 q_59_90 qb_59_90 bit_59_90 bitb_59_90 word59_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_90 q_60_90 qb_60_90 bit_60_90 bitb_60_90 word60_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_90 q_61_90 qb_61_90 bit_61_90 bitb_61_90 word61_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_90 q_62_90 qb_62_90 bit_62_90 bitb_62_90 word62_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_90 q_63_90 qb_63_90 bit_63_90 bitb_63_90 word63_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_90 q_64_90 qb_64_90 bit_64_90 bitb_64_90 word64_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_90 q_65_90 qb_65_90 bit_65_90 bitb_65_90 word65_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_90 q_66_90 qb_66_90 bit_66_90 bitb_66_90 word66_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_90 q_67_90 qb_67_90 bit_67_90 bitb_67_90 word67_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_90 q_68_90 qb_68_90 bit_68_90 bitb_68_90 word68_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_90 q_69_90 qb_69_90 bit_69_90 bitb_69_90 word69_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_90 q_70_90 qb_70_90 bit_70_90 bitb_70_90 word70_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_90 q_71_90 qb_71_90 bit_71_90 bitb_71_90 word71_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_90 q_72_90 qb_72_90 bit_72_90 bitb_72_90 word72_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_90 q_73_90 qb_73_90 bit_73_90 bitb_73_90 word73_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_90 q_74_90 qb_74_90 bit_74_90 bitb_74_90 word74_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_90 q_75_90 qb_75_90 bit_75_90 bitb_75_90 word75_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_90 q_76_90 qb_76_90 bit_76_90 bitb_76_90 word76_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_90 q_77_90 qb_77_90 bit_77_90 bitb_77_90 word77_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_90 q_78_90 qb_78_90 bit_78_90 bitb_78_90 word78_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_90 q_79_90 qb_79_90 bit_79_90 bitb_79_90 word79_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_90 q_80_90 qb_80_90 bit_80_90 bitb_80_90 word80_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_90 q_81_90 qb_81_90 bit_81_90 bitb_81_90 word81_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_90 q_82_90 qb_82_90 bit_82_90 bitb_82_90 word82_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_90 q_83_90 qb_83_90 bit_83_90 bitb_83_90 word83_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_90 q_84_90 qb_84_90 bit_84_90 bitb_84_90 word84_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_90 q_85_90 qb_85_90 bit_85_90 bitb_85_90 word85_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_90 q_86_90 qb_86_90 bit_86_90 bitb_86_90 word86_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_90 q_87_90 qb_87_90 bit_87_90 bitb_87_90 word87_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_90 q_88_90 qb_88_90 bit_88_90 bitb_88_90 word88_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_90 q_89_90 qb_89_90 bit_89_90 bitb_89_90 word89_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_90 q_90_90 qb_90_90 bit_90_90 bitb_90_90 word90_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_90 q_91_90 qb_91_90 bit_91_90 bitb_91_90 word91_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_90 q_92_90 qb_92_90 bit_92_90 bitb_92_90 word92_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_90 q_93_90 qb_93_90 bit_93_90 bitb_93_90 word93_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_90 q_94_90 qb_94_90 bit_94_90 bitb_94_90 word94_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_90 q_95_90 qb_95_90 bit_95_90 bitb_95_90 word95_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_90 q_96_90 qb_96_90 bit_96_90 bitb_96_90 word96_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_90 q_97_90 qb_97_90 bit_97_90 bitb_97_90 word97_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_90 q_98_90 qb_98_90 bit_98_90 bitb_98_90 word98_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_90 q_99_90 qb_99_90 bit_99_90 bitb_99_90 word99_90 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_91 q_0_91 qb_0_91 bit_0_91 bitb_0_91 word0_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_91 q_1_91 qb_1_91 bit_1_91 bitb_1_91 word1_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_91 q_2_91 qb_2_91 bit_2_91 bitb_2_91 word2_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_91 q_3_91 qb_3_91 bit_3_91 bitb_3_91 word3_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_91 q_4_91 qb_4_91 bit_4_91 bitb_4_91 word4_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_91 q_5_91 qb_5_91 bit_5_91 bitb_5_91 word5_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_91 q_6_91 qb_6_91 bit_6_91 bitb_6_91 word6_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_91 q_7_91 qb_7_91 bit_7_91 bitb_7_91 word7_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_91 q_8_91 qb_8_91 bit_8_91 bitb_8_91 word8_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_91 q_9_91 qb_9_91 bit_9_91 bitb_9_91 word9_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_91 q_10_91 qb_10_91 bit_10_91 bitb_10_91 word10_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_91 q_11_91 qb_11_91 bit_11_91 bitb_11_91 word11_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_91 q_12_91 qb_12_91 bit_12_91 bitb_12_91 word12_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_91 q_13_91 qb_13_91 bit_13_91 bitb_13_91 word13_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_91 q_14_91 qb_14_91 bit_14_91 bitb_14_91 word14_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_91 q_15_91 qb_15_91 bit_15_91 bitb_15_91 word15_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_91 q_16_91 qb_16_91 bit_16_91 bitb_16_91 word16_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_91 q_17_91 qb_17_91 bit_17_91 bitb_17_91 word17_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_91 q_18_91 qb_18_91 bit_18_91 bitb_18_91 word18_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_91 q_19_91 qb_19_91 bit_19_91 bitb_19_91 word19_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_91 q_20_91 qb_20_91 bit_20_91 bitb_20_91 word20_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_91 q_21_91 qb_21_91 bit_21_91 bitb_21_91 word21_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_91 q_22_91 qb_22_91 bit_22_91 bitb_22_91 word22_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_91 q_23_91 qb_23_91 bit_23_91 bitb_23_91 word23_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_91 q_24_91 qb_24_91 bit_24_91 bitb_24_91 word24_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_91 q_25_91 qb_25_91 bit_25_91 bitb_25_91 word25_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_91 q_26_91 qb_26_91 bit_26_91 bitb_26_91 word26_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_91 q_27_91 qb_27_91 bit_27_91 bitb_27_91 word27_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_91 q_28_91 qb_28_91 bit_28_91 bitb_28_91 word28_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_91 q_29_91 qb_29_91 bit_29_91 bitb_29_91 word29_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_91 q_30_91 qb_30_91 bit_30_91 bitb_30_91 word30_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_91 q_31_91 qb_31_91 bit_31_91 bitb_31_91 word31_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_91 q_32_91 qb_32_91 bit_32_91 bitb_32_91 word32_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_91 q_33_91 qb_33_91 bit_33_91 bitb_33_91 word33_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_91 q_34_91 qb_34_91 bit_34_91 bitb_34_91 word34_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_91 q_35_91 qb_35_91 bit_35_91 bitb_35_91 word35_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_91 q_36_91 qb_36_91 bit_36_91 bitb_36_91 word36_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_91 q_37_91 qb_37_91 bit_37_91 bitb_37_91 word37_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_91 q_38_91 qb_38_91 bit_38_91 bitb_38_91 word38_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_91 q_39_91 qb_39_91 bit_39_91 bitb_39_91 word39_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_91 q_40_91 qb_40_91 bit_40_91 bitb_40_91 word40_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_91 q_41_91 qb_41_91 bit_41_91 bitb_41_91 word41_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_91 q_42_91 qb_42_91 bit_42_91 bitb_42_91 word42_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_91 q_43_91 qb_43_91 bit_43_91 bitb_43_91 word43_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_91 q_44_91 qb_44_91 bit_44_91 bitb_44_91 word44_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_91 q_45_91 qb_45_91 bit_45_91 bitb_45_91 word45_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_91 q_46_91 qb_46_91 bit_46_91 bitb_46_91 word46_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_91 q_47_91 qb_47_91 bit_47_91 bitb_47_91 word47_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_91 q_48_91 qb_48_91 bit_48_91 bitb_48_91 word48_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_91 q_49_91 qb_49_91 bit_49_91 bitb_49_91 word49_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_91 q_50_91 qb_50_91 bit_50_91 bitb_50_91 word50_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_91 q_51_91 qb_51_91 bit_51_91 bitb_51_91 word51_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_91 q_52_91 qb_52_91 bit_52_91 bitb_52_91 word52_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_91 q_53_91 qb_53_91 bit_53_91 bitb_53_91 word53_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_91 q_54_91 qb_54_91 bit_54_91 bitb_54_91 word54_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_91 q_55_91 qb_55_91 bit_55_91 bitb_55_91 word55_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_91 q_56_91 qb_56_91 bit_56_91 bitb_56_91 word56_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_91 q_57_91 qb_57_91 bit_57_91 bitb_57_91 word57_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_91 q_58_91 qb_58_91 bit_58_91 bitb_58_91 word58_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_91 q_59_91 qb_59_91 bit_59_91 bitb_59_91 word59_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_91 q_60_91 qb_60_91 bit_60_91 bitb_60_91 word60_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_91 q_61_91 qb_61_91 bit_61_91 bitb_61_91 word61_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_91 q_62_91 qb_62_91 bit_62_91 bitb_62_91 word62_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_91 q_63_91 qb_63_91 bit_63_91 bitb_63_91 word63_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_91 q_64_91 qb_64_91 bit_64_91 bitb_64_91 word64_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_91 q_65_91 qb_65_91 bit_65_91 bitb_65_91 word65_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_91 q_66_91 qb_66_91 bit_66_91 bitb_66_91 word66_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_91 q_67_91 qb_67_91 bit_67_91 bitb_67_91 word67_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_91 q_68_91 qb_68_91 bit_68_91 bitb_68_91 word68_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_91 q_69_91 qb_69_91 bit_69_91 bitb_69_91 word69_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_91 q_70_91 qb_70_91 bit_70_91 bitb_70_91 word70_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_91 q_71_91 qb_71_91 bit_71_91 bitb_71_91 word71_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_91 q_72_91 qb_72_91 bit_72_91 bitb_72_91 word72_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_91 q_73_91 qb_73_91 bit_73_91 bitb_73_91 word73_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_91 q_74_91 qb_74_91 bit_74_91 bitb_74_91 word74_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_91 q_75_91 qb_75_91 bit_75_91 bitb_75_91 word75_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_91 q_76_91 qb_76_91 bit_76_91 bitb_76_91 word76_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_91 q_77_91 qb_77_91 bit_77_91 bitb_77_91 word77_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_91 q_78_91 qb_78_91 bit_78_91 bitb_78_91 word78_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_91 q_79_91 qb_79_91 bit_79_91 bitb_79_91 word79_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_91 q_80_91 qb_80_91 bit_80_91 bitb_80_91 word80_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_91 q_81_91 qb_81_91 bit_81_91 bitb_81_91 word81_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_91 q_82_91 qb_82_91 bit_82_91 bitb_82_91 word82_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_91 q_83_91 qb_83_91 bit_83_91 bitb_83_91 word83_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_91 q_84_91 qb_84_91 bit_84_91 bitb_84_91 word84_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_91 q_85_91 qb_85_91 bit_85_91 bitb_85_91 word85_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_91 q_86_91 qb_86_91 bit_86_91 bitb_86_91 word86_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_91 q_87_91 qb_87_91 bit_87_91 bitb_87_91 word87_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_91 q_88_91 qb_88_91 bit_88_91 bitb_88_91 word88_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_91 q_89_91 qb_89_91 bit_89_91 bitb_89_91 word89_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_91 q_90_91 qb_90_91 bit_90_91 bitb_90_91 word90_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_91 q_91_91 qb_91_91 bit_91_91 bitb_91_91 word91_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_91 q_92_91 qb_92_91 bit_92_91 bitb_92_91 word92_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_91 q_93_91 qb_93_91 bit_93_91 bitb_93_91 word93_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_91 q_94_91 qb_94_91 bit_94_91 bitb_94_91 word94_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_91 q_95_91 qb_95_91 bit_95_91 bitb_95_91 word95_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_91 q_96_91 qb_96_91 bit_96_91 bitb_96_91 word96_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_91 q_97_91 qb_97_91 bit_97_91 bitb_97_91 word97_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_91 q_98_91 qb_98_91 bit_98_91 bitb_98_91 word98_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_91 q_99_91 qb_99_91 bit_99_91 bitb_99_91 word99_91 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_92 q_0_92 qb_0_92 bit_0_92 bitb_0_92 word0_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_92 q_1_92 qb_1_92 bit_1_92 bitb_1_92 word1_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_92 q_2_92 qb_2_92 bit_2_92 bitb_2_92 word2_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_92 q_3_92 qb_3_92 bit_3_92 bitb_3_92 word3_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_92 q_4_92 qb_4_92 bit_4_92 bitb_4_92 word4_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_92 q_5_92 qb_5_92 bit_5_92 bitb_5_92 word5_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_92 q_6_92 qb_6_92 bit_6_92 bitb_6_92 word6_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_92 q_7_92 qb_7_92 bit_7_92 bitb_7_92 word7_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_92 q_8_92 qb_8_92 bit_8_92 bitb_8_92 word8_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_92 q_9_92 qb_9_92 bit_9_92 bitb_9_92 word9_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_92 q_10_92 qb_10_92 bit_10_92 bitb_10_92 word10_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_92 q_11_92 qb_11_92 bit_11_92 bitb_11_92 word11_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_92 q_12_92 qb_12_92 bit_12_92 bitb_12_92 word12_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_92 q_13_92 qb_13_92 bit_13_92 bitb_13_92 word13_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_92 q_14_92 qb_14_92 bit_14_92 bitb_14_92 word14_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_92 q_15_92 qb_15_92 bit_15_92 bitb_15_92 word15_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_92 q_16_92 qb_16_92 bit_16_92 bitb_16_92 word16_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_92 q_17_92 qb_17_92 bit_17_92 bitb_17_92 word17_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_92 q_18_92 qb_18_92 bit_18_92 bitb_18_92 word18_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_92 q_19_92 qb_19_92 bit_19_92 bitb_19_92 word19_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_92 q_20_92 qb_20_92 bit_20_92 bitb_20_92 word20_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_92 q_21_92 qb_21_92 bit_21_92 bitb_21_92 word21_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_92 q_22_92 qb_22_92 bit_22_92 bitb_22_92 word22_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_92 q_23_92 qb_23_92 bit_23_92 bitb_23_92 word23_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_92 q_24_92 qb_24_92 bit_24_92 bitb_24_92 word24_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_92 q_25_92 qb_25_92 bit_25_92 bitb_25_92 word25_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_92 q_26_92 qb_26_92 bit_26_92 bitb_26_92 word26_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_92 q_27_92 qb_27_92 bit_27_92 bitb_27_92 word27_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_92 q_28_92 qb_28_92 bit_28_92 bitb_28_92 word28_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_92 q_29_92 qb_29_92 bit_29_92 bitb_29_92 word29_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_92 q_30_92 qb_30_92 bit_30_92 bitb_30_92 word30_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_92 q_31_92 qb_31_92 bit_31_92 bitb_31_92 word31_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_92 q_32_92 qb_32_92 bit_32_92 bitb_32_92 word32_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_92 q_33_92 qb_33_92 bit_33_92 bitb_33_92 word33_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_92 q_34_92 qb_34_92 bit_34_92 bitb_34_92 word34_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_92 q_35_92 qb_35_92 bit_35_92 bitb_35_92 word35_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_92 q_36_92 qb_36_92 bit_36_92 bitb_36_92 word36_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_92 q_37_92 qb_37_92 bit_37_92 bitb_37_92 word37_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_92 q_38_92 qb_38_92 bit_38_92 bitb_38_92 word38_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_92 q_39_92 qb_39_92 bit_39_92 bitb_39_92 word39_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_92 q_40_92 qb_40_92 bit_40_92 bitb_40_92 word40_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_92 q_41_92 qb_41_92 bit_41_92 bitb_41_92 word41_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_92 q_42_92 qb_42_92 bit_42_92 bitb_42_92 word42_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_92 q_43_92 qb_43_92 bit_43_92 bitb_43_92 word43_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_92 q_44_92 qb_44_92 bit_44_92 bitb_44_92 word44_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_92 q_45_92 qb_45_92 bit_45_92 bitb_45_92 word45_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_92 q_46_92 qb_46_92 bit_46_92 bitb_46_92 word46_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_92 q_47_92 qb_47_92 bit_47_92 bitb_47_92 word47_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_92 q_48_92 qb_48_92 bit_48_92 bitb_48_92 word48_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_92 q_49_92 qb_49_92 bit_49_92 bitb_49_92 word49_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_92 q_50_92 qb_50_92 bit_50_92 bitb_50_92 word50_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_92 q_51_92 qb_51_92 bit_51_92 bitb_51_92 word51_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_92 q_52_92 qb_52_92 bit_52_92 bitb_52_92 word52_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_92 q_53_92 qb_53_92 bit_53_92 bitb_53_92 word53_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_92 q_54_92 qb_54_92 bit_54_92 bitb_54_92 word54_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_92 q_55_92 qb_55_92 bit_55_92 bitb_55_92 word55_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_92 q_56_92 qb_56_92 bit_56_92 bitb_56_92 word56_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_92 q_57_92 qb_57_92 bit_57_92 bitb_57_92 word57_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_92 q_58_92 qb_58_92 bit_58_92 bitb_58_92 word58_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_92 q_59_92 qb_59_92 bit_59_92 bitb_59_92 word59_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_92 q_60_92 qb_60_92 bit_60_92 bitb_60_92 word60_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_92 q_61_92 qb_61_92 bit_61_92 bitb_61_92 word61_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_92 q_62_92 qb_62_92 bit_62_92 bitb_62_92 word62_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_92 q_63_92 qb_63_92 bit_63_92 bitb_63_92 word63_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_92 q_64_92 qb_64_92 bit_64_92 bitb_64_92 word64_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_92 q_65_92 qb_65_92 bit_65_92 bitb_65_92 word65_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_92 q_66_92 qb_66_92 bit_66_92 bitb_66_92 word66_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_92 q_67_92 qb_67_92 bit_67_92 bitb_67_92 word67_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_92 q_68_92 qb_68_92 bit_68_92 bitb_68_92 word68_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_92 q_69_92 qb_69_92 bit_69_92 bitb_69_92 word69_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_92 q_70_92 qb_70_92 bit_70_92 bitb_70_92 word70_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_92 q_71_92 qb_71_92 bit_71_92 bitb_71_92 word71_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_92 q_72_92 qb_72_92 bit_72_92 bitb_72_92 word72_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_92 q_73_92 qb_73_92 bit_73_92 bitb_73_92 word73_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_92 q_74_92 qb_74_92 bit_74_92 bitb_74_92 word74_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_92 q_75_92 qb_75_92 bit_75_92 bitb_75_92 word75_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_92 q_76_92 qb_76_92 bit_76_92 bitb_76_92 word76_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_92 q_77_92 qb_77_92 bit_77_92 bitb_77_92 word77_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_92 q_78_92 qb_78_92 bit_78_92 bitb_78_92 word78_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_92 q_79_92 qb_79_92 bit_79_92 bitb_79_92 word79_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_92 q_80_92 qb_80_92 bit_80_92 bitb_80_92 word80_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_92 q_81_92 qb_81_92 bit_81_92 bitb_81_92 word81_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_92 q_82_92 qb_82_92 bit_82_92 bitb_82_92 word82_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_92 q_83_92 qb_83_92 bit_83_92 bitb_83_92 word83_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_92 q_84_92 qb_84_92 bit_84_92 bitb_84_92 word84_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_92 q_85_92 qb_85_92 bit_85_92 bitb_85_92 word85_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_92 q_86_92 qb_86_92 bit_86_92 bitb_86_92 word86_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_92 q_87_92 qb_87_92 bit_87_92 bitb_87_92 word87_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_92 q_88_92 qb_88_92 bit_88_92 bitb_88_92 word88_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_92 q_89_92 qb_89_92 bit_89_92 bitb_89_92 word89_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_92 q_90_92 qb_90_92 bit_90_92 bitb_90_92 word90_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_92 q_91_92 qb_91_92 bit_91_92 bitb_91_92 word91_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_92 q_92_92 qb_92_92 bit_92_92 bitb_92_92 word92_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_92 q_93_92 qb_93_92 bit_93_92 bitb_93_92 word93_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_92 q_94_92 qb_94_92 bit_94_92 bitb_94_92 word94_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_92 q_95_92 qb_95_92 bit_95_92 bitb_95_92 word95_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_92 q_96_92 qb_96_92 bit_96_92 bitb_96_92 word96_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_92 q_97_92 qb_97_92 bit_97_92 bitb_97_92 word97_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_92 q_98_92 qb_98_92 bit_98_92 bitb_98_92 word98_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_92 q_99_92 qb_99_92 bit_99_92 bitb_99_92 word99_92 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_93 q_0_93 qb_0_93 bit_0_93 bitb_0_93 word0_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_93 q_1_93 qb_1_93 bit_1_93 bitb_1_93 word1_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_93 q_2_93 qb_2_93 bit_2_93 bitb_2_93 word2_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_93 q_3_93 qb_3_93 bit_3_93 bitb_3_93 word3_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_93 q_4_93 qb_4_93 bit_4_93 bitb_4_93 word4_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_93 q_5_93 qb_5_93 bit_5_93 bitb_5_93 word5_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_93 q_6_93 qb_6_93 bit_6_93 bitb_6_93 word6_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_93 q_7_93 qb_7_93 bit_7_93 bitb_7_93 word7_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_93 q_8_93 qb_8_93 bit_8_93 bitb_8_93 word8_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_93 q_9_93 qb_9_93 bit_9_93 bitb_9_93 word9_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_93 q_10_93 qb_10_93 bit_10_93 bitb_10_93 word10_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_93 q_11_93 qb_11_93 bit_11_93 bitb_11_93 word11_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_93 q_12_93 qb_12_93 bit_12_93 bitb_12_93 word12_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_93 q_13_93 qb_13_93 bit_13_93 bitb_13_93 word13_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_93 q_14_93 qb_14_93 bit_14_93 bitb_14_93 word14_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_93 q_15_93 qb_15_93 bit_15_93 bitb_15_93 word15_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_93 q_16_93 qb_16_93 bit_16_93 bitb_16_93 word16_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_93 q_17_93 qb_17_93 bit_17_93 bitb_17_93 word17_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_93 q_18_93 qb_18_93 bit_18_93 bitb_18_93 word18_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_93 q_19_93 qb_19_93 bit_19_93 bitb_19_93 word19_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_93 q_20_93 qb_20_93 bit_20_93 bitb_20_93 word20_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_93 q_21_93 qb_21_93 bit_21_93 bitb_21_93 word21_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_93 q_22_93 qb_22_93 bit_22_93 bitb_22_93 word22_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_93 q_23_93 qb_23_93 bit_23_93 bitb_23_93 word23_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_93 q_24_93 qb_24_93 bit_24_93 bitb_24_93 word24_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_93 q_25_93 qb_25_93 bit_25_93 bitb_25_93 word25_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_93 q_26_93 qb_26_93 bit_26_93 bitb_26_93 word26_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_93 q_27_93 qb_27_93 bit_27_93 bitb_27_93 word27_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_93 q_28_93 qb_28_93 bit_28_93 bitb_28_93 word28_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_93 q_29_93 qb_29_93 bit_29_93 bitb_29_93 word29_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_93 q_30_93 qb_30_93 bit_30_93 bitb_30_93 word30_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_93 q_31_93 qb_31_93 bit_31_93 bitb_31_93 word31_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_93 q_32_93 qb_32_93 bit_32_93 bitb_32_93 word32_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_93 q_33_93 qb_33_93 bit_33_93 bitb_33_93 word33_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_93 q_34_93 qb_34_93 bit_34_93 bitb_34_93 word34_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_93 q_35_93 qb_35_93 bit_35_93 bitb_35_93 word35_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_93 q_36_93 qb_36_93 bit_36_93 bitb_36_93 word36_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_93 q_37_93 qb_37_93 bit_37_93 bitb_37_93 word37_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_93 q_38_93 qb_38_93 bit_38_93 bitb_38_93 word38_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_93 q_39_93 qb_39_93 bit_39_93 bitb_39_93 word39_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_93 q_40_93 qb_40_93 bit_40_93 bitb_40_93 word40_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_93 q_41_93 qb_41_93 bit_41_93 bitb_41_93 word41_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_93 q_42_93 qb_42_93 bit_42_93 bitb_42_93 word42_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_93 q_43_93 qb_43_93 bit_43_93 bitb_43_93 word43_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_93 q_44_93 qb_44_93 bit_44_93 bitb_44_93 word44_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_93 q_45_93 qb_45_93 bit_45_93 bitb_45_93 word45_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_93 q_46_93 qb_46_93 bit_46_93 bitb_46_93 word46_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_93 q_47_93 qb_47_93 bit_47_93 bitb_47_93 word47_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_93 q_48_93 qb_48_93 bit_48_93 bitb_48_93 word48_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_93 q_49_93 qb_49_93 bit_49_93 bitb_49_93 word49_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_93 q_50_93 qb_50_93 bit_50_93 bitb_50_93 word50_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_93 q_51_93 qb_51_93 bit_51_93 bitb_51_93 word51_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_93 q_52_93 qb_52_93 bit_52_93 bitb_52_93 word52_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_93 q_53_93 qb_53_93 bit_53_93 bitb_53_93 word53_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_93 q_54_93 qb_54_93 bit_54_93 bitb_54_93 word54_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_93 q_55_93 qb_55_93 bit_55_93 bitb_55_93 word55_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_93 q_56_93 qb_56_93 bit_56_93 bitb_56_93 word56_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_93 q_57_93 qb_57_93 bit_57_93 bitb_57_93 word57_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_93 q_58_93 qb_58_93 bit_58_93 bitb_58_93 word58_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_93 q_59_93 qb_59_93 bit_59_93 bitb_59_93 word59_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_93 q_60_93 qb_60_93 bit_60_93 bitb_60_93 word60_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_93 q_61_93 qb_61_93 bit_61_93 bitb_61_93 word61_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_93 q_62_93 qb_62_93 bit_62_93 bitb_62_93 word62_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_93 q_63_93 qb_63_93 bit_63_93 bitb_63_93 word63_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_93 q_64_93 qb_64_93 bit_64_93 bitb_64_93 word64_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_93 q_65_93 qb_65_93 bit_65_93 bitb_65_93 word65_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_93 q_66_93 qb_66_93 bit_66_93 bitb_66_93 word66_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_93 q_67_93 qb_67_93 bit_67_93 bitb_67_93 word67_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_93 q_68_93 qb_68_93 bit_68_93 bitb_68_93 word68_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_93 q_69_93 qb_69_93 bit_69_93 bitb_69_93 word69_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_93 q_70_93 qb_70_93 bit_70_93 bitb_70_93 word70_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_93 q_71_93 qb_71_93 bit_71_93 bitb_71_93 word71_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_93 q_72_93 qb_72_93 bit_72_93 bitb_72_93 word72_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_93 q_73_93 qb_73_93 bit_73_93 bitb_73_93 word73_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_93 q_74_93 qb_74_93 bit_74_93 bitb_74_93 word74_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_93 q_75_93 qb_75_93 bit_75_93 bitb_75_93 word75_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_93 q_76_93 qb_76_93 bit_76_93 bitb_76_93 word76_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_93 q_77_93 qb_77_93 bit_77_93 bitb_77_93 word77_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_93 q_78_93 qb_78_93 bit_78_93 bitb_78_93 word78_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_93 q_79_93 qb_79_93 bit_79_93 bitb_79_93 word79_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_93 q_80_93 qb_80_93 bit_80_93 bitb_80_93 word80_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_93 q_81_93 qb_81_93 bit_81_93 bitb_81_93 word81_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_93 q_82_93 qb_82_93 bit_82_93 bitb_82_93 word82_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_93 q_83_93 qb_83_93 bit_83_93 bitb_83_93 word83_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_93 q_84_93 qb_84_93 bit_84_93 bitb_84_93 word84_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_93 q_85_93 qb_85_93 bit_85_93 bitb_85_93 word85_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_93 q_86_93 qb_86_93 bit_86_93 bitb_86_93 word86_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_93 q_87_93 qb_87_93 bit_87_93 bitb_87_93 word87_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_93 q_88_93 qb_88_93 bit_88_93 bitb_88_93 word88_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_93 q_89_93 qb_89_93 bit_89_93 bitb_89_93 word89_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_93 q_90_93 qb_90_93 bit_90_93 bitb_90_93 word90_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_93 q_91_93 qb_91_93 bit_91_93 bitb_91_93 word91_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_93 q_92_93 qb_92_93 bit_92_93 bitb_92_93 word92_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_93 q_93_93 qb_93_93 bit_93_93 bitb_93_93 word93_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_93 q_94_93 qb_94_93 bit_94_93 bitb_94_93 word94_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_93 q_95_93 qb_95_93 bit_95_93 bitb_95_93 word95_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_93 q_96_93 qb_96_93 bit_96_93 bitb_96_93 word96_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_93 q_97_93 qb_97_93 bit_97_93 bitb_97_93 word97_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_93 q_98_93 qb_98_93 bit_98_93 bitb_98_93 word98_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_93 q_99_93 qb_99_93 bit_99_93 bitb_99_93 word99_93 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_94 q_0_94 qb_0_94 bit_0_94 bitb_0_94 word0_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_94 q_1_94 qb_1_94 bit_1_94 bitb_1_94 word1_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_94 q_2_94 qb_2_94 bit_2_94 bitb_2_94 word2_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_94 q_3_94 qb_3_94 bit_3_94 bitb_3_94 word3_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_94 q_4_94 qb_4_94 bit_4_94 bitb_4_94 word4_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_94 q_5_94 qb_5_94 bit_5_94 bitb_5_94 word5_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_94 q_6_94 qb_6_94 bit_6_94 bitb_6_94 word6_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_94 q_7_94 qb_7_94 bit_7_94 bitb_7_94 word7_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_94 q_8_94 qb_8_94 bit_8_94 bitb_8_94 word8_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_94 q_9_94 qb_9_94 bit_9_94 bitb_9_94 word9_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_94 q_10_94 qb_10_94 bit_10_94 bitb_10_94 word10_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_94 q_11_94 qb_11_94 bit_11_94 bitb_11_94 word11_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_94 q_12_94 qb_12_94 bit_12_94 bitb_12_94 word12_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_94 q_13_94 qb_13_94 bit_13_94 bitb_13_94 word13_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_94 q_14_94 qb_14_94 bit_14_94 bitb_14_94 word14_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_94 q_15_94 qb_15_94 bit_15_94 bitb_15_94 word15_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_94 q_16_94 qb_16_94 bit_16_94 bitb_16_94 word16_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_94 q_17_94 qb_17_94 bit_17_94 bitb_17_94 word17_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_94 q_18_94 qb_18_94 bit_18_94 bitb_18_94 word18_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_94 q_19_94 qb_19_94 bit_19_94 bitb_19_94 word19_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_94 q_20_94 qb_20_94 bit_20_94 bitb_20_94 word20_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_94 q_21_94 qb_21_94 bit_21_94 bitb_21_94 word21_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_94 q_22_94 qb_22_94 bit_22_94 bitb_22_94 word22_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_94 q_23_94 qb_23_94 bit_23_94 bitb_23_94 word23_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_94 q_24_94 qb_24_94 bit_24_94 bitb_24_94 word24_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_94 q_25_94 qb_25_94 bit_25_94 bitb_25_94 word25_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_94 q_26_94 qb_26_94 bit_26_94 bitb_26_94 word26_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_94 q_27_94 qb_27_94 bit_27_94 bitb_27_94 word27_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_94 q_28_94 qb_28_94 bit_28_94 bitb_28_94 word28_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_94 q_29_94 qb_29_94 bit_29_94 bitb_29_94 word29_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_94 q_30_94 qb_30_94 bit_30_94 bitb_30_94 word30_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_94 q_31_94 qb_31_94 bit_31_94 bitb_31_94 word31_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_94 q_32_94 qb_32_94 bit_32_94 bitb_32_94 word32_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_94 q_33_94 qb_33_94 bit_33_94 bitb_33_94 word33_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_94 q_34_94 qb_34_94 bit_34_94 bitb_34_94 word34_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_94 q_35_94 qb_35_94 bit_35_94 bitb_35_94 word35_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_94 q_36_94 qb_36_94 bit_36_94 bitb_36_94 word36_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_94 q_37_94 qb_37_94 bit_37_94 bitb_37_94 word37_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_94 q_38_94 qb_38_94 bit_38_94 bitb_38_94 word38_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_94 q_39_94 qb_39_94 bit_39_94 bitb_39_94 word39_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_94 q_40_94 qb_40_94 bit_40_94 bitb_40_94 word40_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_94 q_41_94 qb_41_94 bit_41_94 bitb_41_94 word41_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_94 q_42_94 qb_42_94 bit_42_94 bitb_42_94 word42_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_94 q_43_94 qb_43_94 bit_43_94 bitb_43_94 word43_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_94 q_44_94 qb_44_94 bit_44_94 bitb_44_94 word44_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_94 q_45_94 qb_45_94 bit_45_94 bitb_45_94 word45_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_94 q_46_94 qb_46_94 bit_46_94 bitb_46_94 word46_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_94 q_47_94 qb_47_94 bit_47_94 bitb_47_94 word47_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_94 q_48_94 qb_48_94 bit_48_94 bitb_48_94 word48_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_94 q_49_94 qb_49_94 bit_49_94 bitb_49_94 word49_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_94 q_50_94 qb_50_94 bit_50_94 bitb_50_94 word50_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_94 q_51_94 qb_51_94 bit_51_94 bitb_51_94 word51_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_94 q_52_94 qb_52_94 bit_52_94 bitb_52_94 word52_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_94 q_53_94 qb_53_94 bit_53_94 bitb_53_94 word53_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_94 q_54_94 qb_54_94 bit_54_94 bitb_54_94 word54_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_94 q_55_94 qb_55_94 bit_55_94 bitb_55_94 word55_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_94 q_56_94 qb_56_94 bit_56_94 bitb_56_94 word56_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_94 q_57_94 qb_57_94 bit_57_94 bitb_57_94 word57_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_94 q_58_94 qb_58_94 bit_58_94 bitb_58_94 word58_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_94 q_59_94 qb_59_94 bit_59_94 bitb_59_94 word59_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_94 q_60_94 qb_60_94 bit_60_94 bitb_60_94 word60_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_94 q_61_94 qb_61_94 bit_61_94 bitb_61_94 word61_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_94 q_62_94 qb_62_94 bit_62_94 bitb_62_94 word62_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_94 q_63_94 qb_63_94 bit_63_94 bitb_63_94 word63_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_94 q_64_94 qb_64_94 bit_64_94 bitb_64_94 word64_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_94 q_65_94 qb_65_94 bit_65_94 bitb_65_94 word65_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_94 q_66_94 qb_66_94 bit_66_94 bitb_66_94 word66_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_94 q_67_94 qb_67_94 bit_67_94 bitb_67_94 word67_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_94 q_68_94 qb_68_94 bit_68_94 bitb_68_94 word68_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_94 q_69_94 qb_69_94 bit_69_94 bitb_69_94 word69_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_94 q_70_94 qb_70_94 bit_70_94 bitb_70_94 word70_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_94 q_71_94 qb_71_94 bit_71_94 bitb_71_94 word71_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_94 q_72_94 qb_72_94 bit_72_94 bitb_72_94 word72_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_94 q_73_94 qb_73_94 bit_73_94 bitb_73_94 word73_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_94 q_74_94 qb_74_94 bit_74_94 bitb_74_94 word74_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_94 q_75_94 qb_75_94 bit_75_94 bitb_75_94 word75_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_94 q_76_94 qb_76_94 bit_76_94 bitb_76_94 word76_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_94 q_77_94 qb_77_94 bit_77_94 bitb_77_94 word77_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_94 q_78_94 qb_78_94 bit_78_94 bitb_78_94 word78_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_94 q_79_94 qb_79_94 bit_79_94 bitb_79_94 word79_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_94 q_80_94 qb_80_94 bit_80_94 bitb_80_94 word80_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_94 q_81_94 qb_81_94 bit_81_94 bitb_81_94 word81_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_94 q_82_94 qb_82_94 bit_82_94 bitb_82_94 word82_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_94 q_83_94 qb_83_94 bit_83_94 bitb_83_94 word83_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_94 q_84_94 qb_84_94 bit_84_94 bitb_84_94 word84_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_94 q_85_94 qb_85_94 bit_85_94 bitb_85_94 word85_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_94 q_86_94 qb_86_94 bit_86_94 bitb_86_94 word86_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_94 q_87_94 qb_87_94 bit_87_94 bitb_87_94 word87_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_94 q_88_94 qb_88_94 bit_88_94 bitb_88_94 word88_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_94 q_89_94 qb_89_94 bit_89_94 bitb_89_94 word89_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_94 q_90_94 qb_90_94 bit_90_94 bitb_90_94 word90_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_94 q_91_94 qb_91_94 bit_91_94 bitb_91_94 word91_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_94 q_92_94 qb_92_94 bit_92_94 bitb_92_94 word92_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_94 q_93_94 qb_93_94 bit_93_94 bitb_93_94 word93_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_94 q_94_94 qb_94_94 bit_94_94 bitb_94_94 word94_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_94 q_95_94 qb_95_94 bit_95_94 bitb_95_94 word95_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_94 q_96_94 qb_96_94 bit_96_94 bitb_96_94 word96_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_94 q_97_94 qb_97_94 bit_97_94 bitb_97_94 word97_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_94 q_98_94 qb_98_94 bit_98_94 bitb_98_94 word98_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_94 q_99_94 qb_99_94 bit_99_94 bitb_99_94 word99_94 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_95 q_0_95 qb_0_95 bit_0_95 bitb_0_95 word0_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_95 q_1_95 qb_1_95 bit_1_95 bitb_1_95 word1_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_95 q_2_95 qb_2_95 bit_2_95 bitb_2_95 word2_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_95 q_3_95 qb_3_95 bit_3_95 bitb_3_95 word3_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_95 q_4_95 qb_4_95 bit_4_95 bitb_4_95 word4_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_95 q_5_95 qb_5_95 bit_5_95 bitb_5_95 word5_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_95 q_6_95 qb_6_95 bit_6_95 bitb_6_95 word6_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_95 q_7_95 qb_7_95 bit_7_95 bitb_7_95 word7_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_95 q_8_95 qb_8_95 bit_8_95 bitb_8_95 word8_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_95 q_9_95 qb_9_95 bit_9_95 bitb_9_95 word9_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_95 q_10_95 qb_10_95 bit_10_95 bitb_10_95 word10_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_95 q_11_95 qb_11_95 bit_11_95 bitb_11_95 word11_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_95 q_12_95 qb_12_95 bit_12_95 bitb_12_95 word12_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_95 q_13_95 qb_13_95 bit_13_95 bitb_13_95 word13_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_95 q_14_95 qb_14_95 bit_14_95 bitb_14_95 word14_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_95 q_15_95 qb_15_95 bit_15_95 bitb_15_95 word15_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_95 q_16_95 qb_16_95 bit_16_95 bitb_16_95 word16_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_95 q_17_95 qb_17_95 bit_17_95 bitb_17_95 word17_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_95 q_18_95 qb_18_95 bit_18_95 bitb_18_95 word18_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_95 q_19_95 qb_19_95 bit_19_95 bitb_19_95 word19_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_95 q_20_95 qb_20_95 bit_20_95 bitb_20_95 word20_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_95 q_21_95 qb_21_95 bit_21_95 bitb_21_95 word21_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_95 q_22_95 qb_22_95 bit_22_95 bitb_22_95 word22_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_95 q_23_95 qb_23_95 bit_23_95 bitb_23_95 word23_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_95 q_24_95 qb_24_95 bit_24_95 bitb_24_95 word24_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_95 q_25_95 qb_25_95 bit_25_95 bitb_25_95 word25_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_95 q_26_95 qb_26_95 bit_26_95 bitb_26_95 word26_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_95 q_27_95 qb_27_95 bit_27_95 bitb_27_95 word27_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_95 q_28_95 qb_28_95 bit_28_95 bitb_28_95 word28_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_95 q_29_95 qb_29_95 bit_29_95 bitb_29_95 word29_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_95 q_30_95 qb_30_95 bit_30_95 bitb_30_95 word30_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_95 q_31_95 qb_31_95 bit_31_95 bitb_31_95 word31_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_95 q_32_95 qb_32_95 bit_32_95 bitb_32_95 word32_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_95 q_33_95 qb_33_95 bit_33_95 bitb_33_95 word33_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_95 q_34_95 qb_34_95 bit_34_95 bitb_34_95 word34_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_95 q_35_95 qb_35_95 bit_35_95 bitb_35_95 word35_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_95 q_36_95 qb_36_95 bit_36_95 bitb_36_95 word36_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_95 q_37_95 qb_37_95 bit_37_95 bitb_37_95 word37_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_95 q_38_95 qb_38_95 bit_38_95 bitb_38_95 word38_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_95 q_39_95 qb_39_95 bit_39_95 bitb_39_95 word39_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_95 q_40_95 qb_40_95 bit_40_95 bitb_40_95 word40_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_95 q_41_95 qb_41_95 bit_41_95 bitb_41_95 word41_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_95 q_42_95 qb_42_95 bit_42_95 bitb_42_95 word42_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_95 q_43_95 qb_43_95 bit_43_95 bitb_43_95 word43_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_95 q_44_95 qb_44_95 bit_44_95 bitb_44_95 word44_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_95 q_45_95 qb_45_95 bit_45_95 bitb_45_95 word45_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_95 q_46_95 qb_46_95 bit_46_95 bitb_46_95 word46_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_95 q_47_95 qb_47_95 bit_47_95 bitb_47_95 word47_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_95 q_48_95 qb_48_95 bit_48_95 bitb_48_95 word48_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_95 q_49_95 qb_49_95 bit_49_95 bitb_49_95 word49_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_95 q_50_95 qb_50_95 bit_50_95 bitb_50_95 word50_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_95 q_51_95 qb_51_95 bit_51_95 bitb_51_95 word51_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_95 q_52_95 qb_52_95 bit_52_95 bitb_52_95 word52_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_95 q_53_95 qb_53_95 bit_53_95 bitb_53_95 word53_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_95 q_54_95 qb_54_95 bit_54_95 bitb_54_95 word54_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_95 q_55_95 qb_55_95 bit_55_95 bitb_55_95 word55_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_95 q_56_95 qb_56_95 bit_56_95 bitb_56_95 word56_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_95 q_57_95 qb_57_95 bit_57_95 bitb_57_95 word57_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_95 q_58_95 qb_58_95 bit_58_95 bitb_58_95 word58_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_95 q_59_95 qb_59_95 bit_59_95 bitb_59_95 word59_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_95 q_60_95 qb_60_95 bit_60_95 bitb_60_95 word60_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_95 q_61_95 qb_61_95 bit_61_95 bitb_61_95 word61_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_95 q_62_95 qb_62_95 bit_62_95 bitb_62_95 word62_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_95 q_63_95 qb_63_95 bit_63_95 bitb_63_95 word63_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_95 q_64_95 qb_64_95 bit_64_95 bitb_64_95 word64_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_95 q_65_95 qb_65_95 bit_65_95 bitb_65_95 word65_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_95 q_66_95 qb_66_95 bit_66_95 bitb_66_95 word66_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_95 q_67_95 qb_67_95 bit_67_95 bitb_67_95 word67_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_95 q_68_95 qb_68_95 bit_68_95 bitb_68_95 word68_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_95 q_69_95 qb_69_95 bit_69_95 bitb_69_95 word69_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_95 q_70_95 qb_70_95 bit_70_95 bitb_70_95 word70_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_95 q_71_95 qb_71_95 bit_71_95 bitb_71_95 word71_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_95 q_72_95 qb_72_95 bit_72_95 bitb_72_95 word72_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_95 q_73_95 qb_73_95 bit_73_95 bitb_73_95 word73_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_95 q_74_95 qb_74_95 bit_74_95 bitb_74_95 word74_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_95 q_75_95 qb_75_95 bit_75_95 bitb_75_95 word75_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_95 q_76_95 qb_76_95 bit_76_95 bitb_76_95 word76_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_95 q_77_95 qb_77_95 bit_77_95 bitb_77_95 word77_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_95 q_78_95 qb_78_95 bit_78_95 bitb_78_95 word78_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_95 q_79_95 qb_79_95 bit_79_95 bitb_79_95 word79_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_95 q_80_95 qb_80_95 bit_80_95 bitb_80_95 word80_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_95 q_81_95 qb_81_95 bit_81_95 bitb_81_95 word81_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_95 q_82_95 qb_82_95 bit_82_95 bitb_82_95 word82_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_95 q_83_95 qb_83_95 bit_83_95 bitb_83_95 word83_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_95 q_84_95 qb_84_95 bit_84_95 bitb_84_95 word84_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_95 q_85_95 qb_85_95 bit_85_95 bitb_85_95 word85_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_95 q_86_95 qb_86_95 bit_86_95 bitb_86_95 word86_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_95 q_87_95 qb_87_95 bit_87_95 bitb_87_95 word87_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_95 q_88_95 qb_88_95 bit_88_95 bitb_88_95 word88_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_95 q_89_95 qb_89_95 bit_89_95 bitb_89_95 word89_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_95 q_90_95 qb_90_95 bit_90_95 bitb_90_95 word90_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_95 q_91_95 qb_91_95 bit_91_95 bitb_91_95 word91_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_95 q_92_95 qb_92_95 bit_92_95 bitb_92_95 word92_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_95 q_93_95 qb_93_95 bit_93_95 bitb_93_95 word93_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_95 q_94_95 qb_94_95 bit_94_95 bitb_94_95 word94_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_95 q_95_95 qb_95_95 bit_95_95 bitb_95_95 word95_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_95 q_96_95 qb_96_95 bit_96_95 bitb_96_95 word96_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_95 q_97_95 qb_97_95 bit_97_95 bitb_97_95 word97_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_95 q_98_95 qb_98_95 bit_98_95 bitb_98_95 word98_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_95 q_99_95 qb_99_95 bit_99_95 bitb_99_95 word99_95 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_96 q_0_96 qb_0_96 bit_0_96 bitb_0_96 word0_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_96 q_1_96 qb_1_96 bit_1_96 bitb_1_96 word1_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_96 q_2_96 qb_2_96 bit_2_96 bitb_2_96 word2_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_96 q_3_96 qb_3_96 bit_3_96 bitb_3_96 word3_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_96 q_4_96 qb_4_96 bit_4_96 bitb_4_96 word4_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_96 q_5_96 qb_5_96 bit_5_96 bitb_5_96 word5_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_96 q_6_96 qb_6_96 bit_6_96 bitb_6_96 word6_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_96 q_7_96 qb_7_96 bit_7_96 bitb_7_96 word7_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_96 q_8_96 qb_8_96 bit_8_96 bitb_8_96 word8_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_96 q_9_96 qb_9_96 bit_9_96 bitb_9_96 word9_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_96 q_10_96 qb_10_96 bit_10_96 bitb_10_96 word10_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_96 q_11_96 qb_11_96 bit_11_96 bitb_11_96 word11_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_96 q_12_96 qb_12_96 bit_12_96 bitb_12_96 word12_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_96 q_13_96 qb_13_96 bit_13_96 bitb_13_96 word13_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_96 q_14_96 qb_14_96 bit_14_96 bitb_14_96 word14_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_96 q_15_96 qb_15_96 bit_15_96 bitb_15_96 word15_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_96 q_16_96 qb_16_96 bit_16_96 bitb_16_96 word16_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_96 q_17_96 qb_17_96 bit_17_96 bitb_17_96 word17_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_96 q_18_96 qb_18_96 bit_18_96 bitb_18_96 word18_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_96 q_19_96 qb_19_96 bit_19_96 bitb_19_96 word19_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_96 q_20_96 qb_20_96 bit_20_96 bitb_20_96 word20_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_96 q_21_96 qb_21_96 bit_21_96 bitb_21_96 word21_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_96 q_22_96 qb_22_96 bit_22_96 bitb_22_96 word22_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_96 q_23_96 qb_23_96 bit_23_96 bitb_23_96 word23_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_96 q_24_96 qb_24_96 bit_24_96 bitb_24_96 word24_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_96 q_25_96 qb_25_96 bit_25_96 bitb_25_96 word25_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_96 q_26_96 qb_26_96 bit_26_96 bitb_26_96 word26_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_96 q_27_96 qb_27_96 bit_27_96 bitb_27_96 word27_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_96 q_28_96 qb_28_96 bit_28_96 bitb_28_96 word28_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_96 q_29_96 qb_29_96 bit_29_96 bitb_29_96 word29_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_96 q_30_96 qb_30_96 bit_30_96 bitb_30_96 word30_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_96 q_31_96 qb_31_96 bit_31_96 bitb_31_96 word31_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_96 q_32_96 qb_32_96 bit_32_96 bitb_32_96 word32_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_96 q_33_96 qb_33_96 bit_33_96 bitb_33_96 word33_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_96 q_34_96 qb_34_96 bit_34_96 bitb_34_96 word34_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_96 q_35_96 qb_35_96 bit_35_96 bitb_35_96 word35_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_96 q_36_96 qb_36_96 bit_36_96 bitb_36_96 word36_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_96 q_37_96 qb_37_96 bit_37_96 bitb_37_96 word37_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_96 q_38_96 qb_38_96 bit_38_96 bitb_38_96 word38_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_96 q_39_96 qb_39_96 bit_39_96 bitb_39_96 word39_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_96 q_40_96 qb_40_96 bit_40_96 bitb_40_96 word40_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_96 q_41_96 qb_41_96 bit_41_96 bitb_41_96 word41_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_96 q_42_96 qb_42_96 bit_42_96 bitb_42_96 word42_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_96 q_43_96 qb_43_96 bit_43_96 bitb_43_96 word43_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_96 q_44_96 qb_44_96 bit_44_96 bitb_44_96 word44_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_96 q_45_96 qb_45_96 bit_45_96 bitb_45_96 word45_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_96 q_46_96 qb_46_96 bit_46_96 bitb_46_96 word46_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_96 q_47_96 qb_47_96 bit_47_96 bitb_47_96 word47_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_96 q_48_96 qb_48_96 bit_48_96 bitb_48_96 word48_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_96 q_49_96 qb_49_96 bit_49_96 bitb_49_96 word49_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_96 q_50_96 qb_50_96 bit_50_96 bitb_50_96 word50_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_96 q_51_96 qb_51_96 bit_51_96 bitb_51_96 word51_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_96 q_52_96 qb_52_96 bit_52_96 bitb_52_96 word52_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_96 q_53_96 qb_53_96 bit_53_96 bitb_53_96 word53_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_96 q_54_96 qb_54_96 bit_54_96 bitb_54_96 word54_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_96 q_55_96 qb_55_96 bit_55_96 bitb_55_96 word55_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_96 q_56_96 qb_56_96 bit_56_96 bitb_56_96 word56_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_96 q_57_96 qb_57_96 bit_57_96 bitb_57_96 word57_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_96 q_58_96 qb_58_96 bit_58_96 bitb_58_96 word58_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_96 q_59_96 qb_59_96 bit_59_96 bitb_59_96 word59_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_96 q_60_96 qb_60_96 bit_60_96 bitb_60_96 word60_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_96 q_61_96 qb_61_96 bit_61_96 bitb_61_96 word61_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_96 q_62_96 qb_62_96 bit_62_96 bitb_62_96 word62_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_96 q_63_96 qb_63_96 bit_63_96 bitb_63_96 word63_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_96 q_64_96 qb_64_96 bit_64_96 bitb_64_96 word64_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_96 q_65_96 qb_65_96 bit_65_96 bitb_65_96 word65_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_96 q_66_96 qb_66_96 bit_66_96 bitb_66_96 word66_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_96 q_67_96 qb_67_96 bit_67_96 bitb_67_96 word67_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_96 q_68_96 qb_68_96 bit_68_96 bitb_68_96 word68_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_96 q_69_96 qb_69_96 bit_69_96 bitb_69_96 word69_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_96 q_70_96 qb_70_96 bit_70_96 bitb_70_96 word70_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_96 q_71_96 qb_71_96 bit_71_96 bitb_71_96 word71_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_96 q_72_96 qb_72_96 bit_72_96 bitb_72_96 word72_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_96 q_73_96 qb_73_96 bit_73_96 bitb_73_96 word73_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_96 q_74_96 qb_74_96 bit_74_96 bitb_74_96 word74_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_96 q_75_96 qb_75_96 bit_75_96 bitb_75_96 word75_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_96 q_76_96 qb_76_96 bit_76_96 bitb_76_96 word76_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_96 q_77_96 qb_77_96 bit_77_96 bitb_77_96 word77_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_96 q_78_96 qb_78_96 bit_78_96 bitb_78_96 word78_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_96 q_79_96 qb_79_96 bit_79_96 bitb_79_96 word79_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_96 q_80_96 qb_80_96 bit_80_96 bitb_80_96 word80_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_96 q_81_96 qb_81_96 bit_81_96 bitb_81_96 word81_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_96 q_82_96 qb_82_96 bit_82_96 bitb_82_96 word82_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_96 q_83_96 qb_83_96 bit_83_96 bitb_83_96 word83_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_96 q_84_96 qb_84_96 bit_84_96 bitb_84_96 word84_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_96 q_85_96 qb_85_96 bit_85_96 bitb_85_96 word85_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_96 q_86_96 qb_86_96 bit_86_96 bitb_86_96 word86_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_96 q_87_96 qb_87_96 bit_87_96 bitb_87_96 word87_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_96 q_88_96 qb_88_96 bit_88_96 bitb_88_96 word88_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_96 q_89_96 qb_89_96 bit_89_96 bitb_89_96 word89_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_96 q_90_96 qb_90_96 bit_90_96 bitb_90_96 word90_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_96 q_91_96 qb_91_96 bit_91_96 bitb_91_96 word91_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_96 q_92_96 qb_92_96 bit_92_96 bitb_92_96 word92_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_96 q_93_96 qb_93_96 bit_93_96 bitb_93_96 word93_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_96 q_94_96 qb_94_96 bit_94_96 bitb_94_96 word94_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_96 q_95_96 qb_95_96 bit_95_96 bitb_95_96 word95_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_96 q_96_96 qb_96_96 bit_96_96 bitb_96_96 word96_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_96 q_97_96 qb_97_96 bit_97_96 bitb_97_96 word97_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_96 q_98_96 qb_98_96 bit_98_96 bitb_98_96 word98_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_96 q_99_96 qb_99_96 bit_99_96 bitb_99_96 word99_96 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_97 q_0_97 qb_0_97 bit_0_97 bitb_0_97 word0_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_97 q_1_97 qb_1_97 bit_1_97 bitb_1_97 word1_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_97 q_2_97 qb_2_97 bit_2_97 bitb_2_97 word2_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_97 q_3_97 qb_3_97 bit_3_97 bitb_3_97 word3_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_97 q_4_97 qb_4_97 bit_4_97 bitb_4_97 word4_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_97 q_5_97 qb_5_97 bit_5_97 bitb_5_97 word5_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_97 q_6_97 qb_6_97 bit_6_97 bitb_6_97 word6_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_97 q_7_97 qb_7_97 bit_7_97 bitb_7_97 word7_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_97 q_8_97 qb_8_97 bit_8_97 bitb_8_97 word8_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_97 q_9_97 qb_9_97 bit_9_97 bitb_9_97 word9_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_97 q_10_97 qb_10_97 bit_10_97 bitb_10_97 word10_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_97 q_11_97 qb_11_97 bit_11_97 bitb_11_97 word11_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_97 q_12_97 qb_12_97 bit_12_97 bitb_12_97 word12_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_97 q_13_97 qb_13_97 bit_13_97 bitb_13_97 word13_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_97 q_14_97 qb_14_97 bit_14_97 bitb_14_97 word14_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_97 q_15_97 qb_15_97 bit_15_97 bitb_15_97 word15_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_97 q_16_97 qb_16_97 bit_16_97 bitb_16_97 word16_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_97 q_17_97 qb_17_97 bit_17_97 bitb_17_97 word17_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_97 q_18_97 qb_18_97 bit_18_97 bitb_18_97 word18_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_97 q_19_97 qb_19_97 bit_19_97 bitb_19_97 word19_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_97 q_20_97 qb_20_97 bit_20_97 bitb_20_97 word20_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_97 q_21_97 qb_21_97 bit_21_97 bitb_21_97 word21_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_97 q_22_97 qb_22_97 bit_22_97 bitb_22_97 word22_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_97 q_23_97 qb_23_97 bit_23_97 bitb_23_97 word23_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_97 q_24_97 qb_24_97 bit_24_97 bitb_24_97 word24_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_97 q_25_97 qb_25_97 bit_25_97 bitb_25_97 word25_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_97 q_26_97 qb_26_97 bit_26_97 bitb_26_97 word26_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_97 q_27_97 qb_27_97 bit_27_97 bitb_27_97 word27_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_97 q_28_97 qb_28_97 bit_28_97 bitb_28_97 word28_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_97 q_29_97 qb_29_97 bit_29_97 bitb_29_97 word29_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_97 q_30_97 qb_30_97 bit_30_97 bitb_30_97 word30_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_97 q_31_97 qb_31_97 bit_31_97 bitb_31_97 word31_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_97 q_32_97 qb_32_97 bit_32_97 bitb_32_97 word32_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_97 q_33_97 qb_33_97 bit_33_97 bitb_33_97 word33_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_97 q_34_97 qb_34_97 bit_34_97 bitb_34_97 word34_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_97 q_35_97 qb_35_97 bit_35_97 bitb_35_97 word35_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_97 q_36_97 qb_36_97 bit_36_97 bitb_36_97 word36_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_97 q_37_97 qb_37_97 bit_37_97 bitb_37_97 word37_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_97 q_38_97 qb_38_97 bit_38_97 bitb_38_97 word38_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_97 q_39_97 qb_39_97 bit_39_97 bitb_39_97 word39_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_97 q_40_97 qb_40_97 bit_40_97 bitb_40_97 word40_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_97 q_41_97 qb_41_97 bit_41_97 bitb_41_97 word41_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_97 q_42_97 qb_42_97 bit_42_97 bitb_42_97 word42_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_97 q_43_97 qb_43_97 bit_43_97 bitb_43_97 word43_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_97 q_44_97 qb_44_97 bit_44_97 bitb_44_97 word44_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_97 q_45_97 qb_45_97 bit_45_97 bitb_45_97 word45_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_97 q_46_97 qb_46_97 bit_46_97 bitb_46_97 word46_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_97 q_47_97 qb_47_97 bit_47_97 bitb_47_97 word47_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_97 q_48_97 qb_48_97 bit_48_97 bitb_48_97 word48_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_97 q_49_97 qb_49_97 bit_49_97 bitb_49_97 word49_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_97 q_50_97 qb_50_97 bit_50_97 bitb_50_97 word50_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_97 q_51_97 qb_51_97 bit_51_97 bitb_51_97 word51_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_97 q_52_97 qb_52_97 bit_52_97 bitb_52_97 word52_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_97 q_53_97 qb_53_97 bit_53_97 bitb_53_97 word53_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_97 q_54_97 qb_54_97 bit_54_97 bitb_54_97 word54_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_97 q_55_97 qb_55_97 bit_55_97 bitb_55_97 word55_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_97 q_56_97 qb_56_97 bit_56_97 bitb_56_97 word56_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_97 q_57_97 qb_57_97 bit_57_97 bitb_57_97 word57_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_97 q_58_97 qb_58_97 bit_58_97 bitb_58_97 word58_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_97 q_59_97 qb_59_97 bit_59_97 bitb_59_97 word59_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_97 q_60_97 qb_60_97 bit_60_97 bitb_60_97 word60_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_97 q_61_97 qb_61_97 bit_61_97 bitb_61_97 word61_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_97 q_62_97 qb_62_97 bit_62_97 bitb_62_97 word62_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_97 q_63_97 qb_63_97 bit_63_97 bitb_63_97 word63_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_97 q_64_97 qb_64_97 bit_64_97 bitb_64_97 word64_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_97 q_65_97 qb_65_97 bit_65_97 bitb_65_97 word65_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_97 q_66_97 qb_66_97 bit_66_97 bitb_66_97 word66_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_97 q_67_97 qb_67_97 bit_67_97 bitb_67_97 word67_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_97 q_68_97 qb_68_97 bit_68_97 bitb_68_97 word68_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_97 q_69_97 qb_69_97 bit_69_97 bitb_69_97 word69_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_97 q_70_97 qb_70_97 bit_70_97 bitb_70_97 word70_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_97 q_71_97 qb_71_97 bit_71_97 bitb_71_97 word71_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_97 q_72_97 qb_72_97 bit_72_97 bitb_72_97 word72_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_97 q_73_97 qb_73_97 bit_73_97 bitb_73_97 word73_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_97 q_74_97 qb_74_97 bit_74_97 bitb_74_97 word74_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_97 q_75_97 qb_75_97 bit_75_97 bitb_75_97 word75_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_97 q_76_97 qb_76_97 bit_76_97 bitb_76_97 word76_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_97 q_77_97 qb_77_97 bit_77_97 bitb_77_97 word77_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_97 q_78_97 qb_78_97 bit_78_97 bitb_78_97 word78_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_97 q_79_97 qb_79_97 bit_79_97 bitb_79_97 word79_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_97 q_80_97 qb_80_97 bit_80_97 bitb_80_97 word80_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_97 q_81_97 qb_81_97 bit_81_97 bitb_81_97 word81_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_97 q_82_97 qb_82_97 bit_82_97 bitb_82_97 word82_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_97 q_83_97 qb_83_97 bit_83_97 bitb_83_97 word83_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_97 q_84_97 qb_84_97 bit_84_97 bitb_84_97 word84_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_97 q_85_97 qb_85_97 bit_85_97 bitb_85_97 word85_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_97 q_86_97 qb_86_97 bit_86_97 bitb_86_97 word86_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_97 q_87_97 qb_87_97 bit_87_97 bitb_87_97 word87_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_97 q_88_97 qb_88_97 bit_88_97 bitb_88_97 word88_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_97 q_89_97 qb_89_97 bit_89_97 bitb_89_97 word89_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_97 q_90_97 qb_90_97 bit_90_97 bitb_90_97 word90_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_97 q_91_97 qb_91_97 bit_91_97 bitb_91_97 word91_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_97 q_92_97 qb_92_97 bit_92_97 bitb_92_97 word92_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_97 q_93_97 qb_93_97 bit_93_97 bitb_93_97 word93_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_97 q_94_97 qb_94_97 bit_94_97 bitb_94_97 word94_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_97 q_95_97 qb_95_97 bit_95_97 bitb_95_97 word95_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_97 q_96_97 qb_96_97 bit_96_97 bitb_96_97 word96_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_97 q_97_97 qb_97_97 bit_97_97 bitb_97_97 word97_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_97 q_98_97 qb_98_97 bit_98_97 bitb_98_97 word98_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_97 q_99_97 qb_99_97 bit_99_97 bitb_99_97 word99_97 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_98 q_0_98 qb_0_98 bit_0_98 bitb_0_98 word0_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_98 q_1_98 qb_1_98 bit_1_98 bitb_1_98 word1_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_98 q_2_98 qb_2_98 bit_2_98 bitb_2_98 word2_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_98 q_3_98 qb_3_98 bit_3_98 bitb_3_98 word3_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_98 q_4_98 qb_4_98 bit_4_98 bitb_4_98 word4_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_98 q_5_98 qb_5_98 bit_5_98 bitb_5_98 word5_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_98 q_6_98 qb_6_98 bit_6_98 bitb_6_98 word6_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_98 q_7_98 qb_7_98 bit_7_98 bitb_7_98 word7_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_98 q_8_98 qb_8_98 bit_8_98 bitb_8_98 word8_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_98 q_9_98 qb_9_98 bit_9_98 bitb_9_98 word9_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_98 q_10_98 qb_10_98 bit_10_98 bitb_10_98 word10_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_98 q_11_98 qb_11_98 bit_11_98 bitb_11_98 word11_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_98 q_12_98 qb_12_98 bit_12_98 bitb_12_98 word12_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_98 q_13_98 qb_13_98 bit_13_98 bitb_13_98 word13_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_98 q_14_98 qb_14_98 bit_14_98 bitb_14_98 word14_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_98 q_15_98 qb_15_98 bit_15_98 bitb_15_98 word15_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_98 q_16_98 qb_16_98 bit_16_98 bitb_16_98 word16_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_98 q_17_98 qb_17_98 bit_17_98 bitb_17_98 word17_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_98 q_18_98 qb_18_98 bit_18_98 bitb_18_98 word18_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_98 q_19_98 qb_19_98 bit_19_98 bitb_19_98 word19_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_98 q_20_98 qb_20_98 bit_20_98 bitb_20_98 word20_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_98 q_21_98 qb_21_98 bit_21_98 bitb_21_98 word21_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_98 q_22_98 qb_22_98 bit_22_98 bitb_22_98 word22_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_98 q_23_98 qb_23_98 bit_23_98 bitb_23_98 word23_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_98 q_24_98 qb_24_98 bit_24_98 bitb_24_98 word24_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_98 q_25_98 qb_25_98 bit_25_98 bitb_25_98 word25_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_98 q_26_98 qb_26_98 bit_26_98 bitb_26_98 word26_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_98 q_27_98 qb_27_98 bit_27_98 bitb_27_98 word27_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_98 q_28_98 qb_28_98 bit_28_98 bitb_28_98 word28_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_98 q_29_98 qb_29_98 bit_29_98 bitb_29_98 word29_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_98 q_30_98 qb_30_98 bit_30_98 bitb_30_98 word30_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_98 q_31_98 qb_31_98 bit_31_98 bitb_31_98 word31_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_98 q_32_98 qb_32_98 bit_32_98 bitb_32_98 word32_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_98 q_33_98 qb_33_98 bit_33_98 bitb_33_98 word33_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_98 q_34_98 qb_34_98 bit_34_98 bitb_34_98 word34_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_98 q_35_98 qb_35_98 bit_35_98 bitb_35_98 word35_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_98 q_36_98 qb_36_98 bit_36_98 bitb_36_98 word36_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_98 q_37_98 qb_37_98 bit_37_98 bitb_37_98 word37_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_98 q_38_98 qb_38_98 bit_38_98 bitb_38_98 word38_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_98 q_39_98 qb_39_98 bit_39_98 bitb_39_98 word39_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_98 q_40_98 qb_40_98 bit_40_98 bitb_40_98 word40_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_98 q_41_98 qb_41_98 bit_41_98 bitb_41_98 word41_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_98 q_42_98 qb_42_98 bit_42_98 bitb_42_98 word42_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_98 q_43_98 qb_43_98 bit_43_98 bitb_43_98 word43_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_98 q_44_98 qb_44_98 bit_44_98 bitb_44_98 word44_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_98 q_45_98 qb_45_98 bit_45_98 bitb_45_98 word45_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_98 q_46_98 qb_46_98 bit_46_98 bitb_46_98 word46_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_98 q_47_98 qb_47_98 bit_47_98 bitb_47_98 word47_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_98 q_48_98 qb_48_98 bit_48_98 bitb_48_98 word48_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_98 q_49_98 qb_49_98 bit_49_98 bitb_49_98 word49_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_98 q_50_98 qb_50_98 bit_50_98 bitb_50_98 word50_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_98 q_51_98 qb_51_98 bit_51_98 bitb_51_98 word51_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_98 q_52_98 qb_52_98 bit_52_98 bitb_52_98 word52_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_98 q_53_98 qb_53_98 bit_53_98 bitb_53_98 word53_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_98 q_54_98 qb_54_98 bit_54_98 bitb_54_98 word54_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_98 q_55_98 qb_55_98 bit_55_98 bitb_55_98 word55_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_98 q_56_98 qb_56_98 bit_56_98 bitb_56_98 word56_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_98 q_57_98 qb_57_98 bit_57_98 bitb_57_98 word57_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_98 q_58_98 qb_58_98 bit_58_98 bitb_58_98 word58_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_98 q_59_98 qb_59_98 bit_59_98 bitb_59_98 word59_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_98 q_60_98 qb_60_98 bit_60_98 bitb_60_98 word60_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_98 q_61_98 qb_61_98 bit_61_98 bitb_61_98 word61_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_98 q_62_98 qb_62_98 bit_62_98 bitb_62_98 word62_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_98 q_63_98 qb_63_98 bit_63_98 bitb_63_98 word63_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_98 q_64_98 qb_64_98 bit_64_98 bitb_64_98 word64_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_98 q_65_98 qb_65_98 bit_65_98 bitb_65_98 word65_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_98 q_66_98 qb_66_98 bit_66_98 bitb_66_98 word66_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_98 q_67_98 qb_67_98 bit_67_98 bitb_67_98 word67_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_98 q_68_98 qb_68_98 bit_68_98 bitb_68_98 word68_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_98 q_69_98 qb_69_98 bit_69_98 bitb_69_98 word69_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_98 q_70_98 qb_70_98 bit_70_98 bitb_70_98 word70_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_98 q_71_98 qb_71_98 bit_71_98 bitb_71_98 word71_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_98 q_72_98 qb_72_98 bit_72_98 bitb_72_98 word72_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_98 q_73_98 qb_73_98 bit_73_98 bitb_73_98 word73_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_98 q_74_98 qb_74_98 bit_74_98 bitb_74_98 word74_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_98 q_75_98 qb_75_98 bit_75_98 bitb_75_98 word75_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_98 q_76_98 qb_76_98 bit_76_98 bitb_76_98 word76_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_98 q_77_98 qb_77_98 bit_77_98 bitb_77_98 word77_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_98 q_78_98 qb_78_98 bit_78_98 bitb_78_98 word78_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_98 q_79_98 qb_79_98 bit_79_98 bitb_79_98 word79_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_98 q_80_98 qb_80_98 bit_80_98 bitb_80_98 word80_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_98 q_81_98 qb_81_98 bit_81_98 bitb_81_98 word81_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_98 q_82_98 qb_82_98 bit_82_98 bitb_82_98 word82_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_98 q_83_98 qb_83_98 bit_83_98 bitb_83_98 word83_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_98 q_84_98 qb_84_98 bit_84_98 bitb_84_98 word84_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_98 q_85_98 qb_85_98 bit_85_98 bitb_85_98 word85_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_98 q_86_98 qb_86_98 bit_86_98 bitb_86_98 word86_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_98 q_87_98 qb_87_98 bit_87_98 bitb_87_98 word87_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_98 q_88_98 qb_88_98 bit_88_98 bitb_88_98 word88_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_98 q_89_98 qb_89_98 bit_89_98 bitb_89_98 word89_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_98 q_90_98 qb_90_98 bit_90_98 bitb_90_98 word90_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_98 q_91_98 qb_91_98 bit_91_98 bitb_91_98 word91_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_98 q_92_98 qb_92_98 bit_92_98 bitb_92_98 word92_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_98 q_93_98 qb_93_98 bit_93_98 bitb_93_98 word93_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_98 q_94_98 qb_94_98 bit_94_98 bitb_94_98 word94_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_98 q_95_98 qb_95_98 bit_95_98 bitb_95_98 word95_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_98 q_96_98 qb_96_98 bit_96_98 bitb_96_98 word96_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_98 q_97_98 qb_97_98 bit_97_98 bitb_97_98 word97_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_98 q_98_98 qb_98_98 bit_98_98 bitb_98_98 word98_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_98 q_99_98 qb_99_98 bit_99_98 bitb_99_98 word99_98 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X0_99 q_0_99 qb_0_99 bit_0_99 bitb_0_99 word0_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X1_99 q_1_99 qb_1_99 bit_1_99 bitb_1_99 word1_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X2_99 q_2_99 qb_2_99 bit_2_99 bitb_2_99 word2_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X3_99 q_3_99 qb_3_99 bit_3_99 bitb_3_99 word3_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X4_99 q_4_99 qb_4_99 bit_4_99 bitb_4_99 word4_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X5_99 q_5_99 qb_5_99 bit_5_99 bitb_5_99 word5_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X6_99 q_6_99 qb_6_99 bit_6_99 bitb_6_99 word6_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X7_99 q_7_99 qb_7_99 bit_7_99 bitb_7_99 word7_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X8_99 q_8_99 qb_8_99 bit_8_99 bitb_8_99 word8_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X9_99 q_9_99 qb_9_99 bit_9_99 bitb_9_99 word9_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X10_99 q_10_99 qb_10_99 bit_10_99 bitb_10_99 word10_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X11_99 q_11_99 qb_11_99 bit_11_99 bitb_11_99 word11_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X12_99 q_12_99 qb_12_99 bit_12_99 bitb_12_99 word12_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X13_99 q_13_99 qb_13_99 bit_13_99 bitb_13_99 word13_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X14_99 q_14_99 qb_14_99 bit_14_99 bitb_14_99 word14_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X15_99 q_15_99 qb_15_99 bit_15_99 bitb_15_99 word15_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X16_99 q_16_99 qb_16_99 bit_16_99 bitb_16_99 word16_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X17_99 q_17_99 qb_17_99 bit_17_99 bitb_17_99 word17_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X18_99 q_18_99 qb_18_99 bit_18_99 bitb_18_99 word18_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X19_99 q_19_99 qb_19_99 bit_19_99 bitb_19_99 word19_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X20_99 q_20_99 qb_20_99 bit_20_99 bitb_20_99 word20_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X21_99 q_21_99 qb_21_99 bit_21_99 bitb_21_99 word21_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X22_99 q_22_99 qb_22_99 bit_22_99 bitb_22_99 word22_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X23_99 q_23_99 qb_23_99 bit_23_99 bitb_23_99 word23_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X24_99 q_24_99 qb_24_99 bit_24_99 bitb_24_99 word24_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X25_99 q_25_99 qb_25_99 bit_25_99 bitb_25_99 word25_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X26_99 q_26_99 qb_26_99 bit_26_99 bitb_26_99 word26_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X27_99 q_27_99 qb_27_99 bit_27_99 bitb_27_99 word27_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X28_99 q_28_99 qb_28_99 bit_28_99 bitb_28_99 word28_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X29_99 q_29_99 qb_29_99 bit_29_99 bitb_29_99 word29_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X30_99 q_30_99 qb_30_99 bit_30_99 bitb_30_99 word30_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X31_99 q_31_99 qb_31_99 bit_31_99 bitb_31_99 word31_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X32_99 q_32_99 qb_32_99 bit_32_99 bitb_32_99 word32_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X33_99 q_33_99 qb_33_99 bit_33_99 bitb_33_99 word33_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X34_99 q_34_99 qb_34_99 bit_34_99 bitb_34_99 word34_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X35_99 q_35_99 qb_35_99 bit_35_99 bitb_35_99 word35_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X36_99 q_36_99 qb_36_99 bit_36_99 bitb_36_99 word36_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X37_99 q_37_99 qb_37_99 bit_37_99 bitb_37_99 word37_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X38_99 q_38_99 qb_38_99 bit_38_99 bitb_38_99 word38_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X39_99 q_39_99 qb_39_99 bit_39_99 bitb_39_99 word39_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X40_99 q_40_99 qb_40_99 bit_40_99 bitb_40_99 word40_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X41_99 q_41_99 qb_41_99 bit_41_99 bitb_41_99 word41_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X42_99 q_42_99 qb_42_99 bit_42_99 bitb_42_99 word42_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X43_99 q_43_99 qb_43_99 bit_43_99 bitb_43_99 word43_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X44_99 q_44_99 qb_44_99 bit_44_99 bitb_44_99 word44_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X45_99 q_45_99 qb_45_99 bit_45_99 bitb_45_99 word45_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X46_99 q_46_99 qb_46_99 bit_46_99 bitb_46_99 word46_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X47_99 q_47_99 qb_47_99 bit_47_99 bitb_47_99 word47_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X48_99 q_48_99 qb_48_99 bit_48_99 bitb_48_99 word48_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X49_99 q_49_99 qb_49_99 bit_49_99 bitb_49_99 word49_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X50_99 q_50_99 qb_50_99 bit_50_99 bitb_50_99 word50_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X51_99 q_51_99 qb_51_99 bit_51_99 bitb_51_99 word51_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X52_99 q_52_99 qb_52_99 bit_52_99 bitb_52_99 word52_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X53_99 q_53_99 qb_53_99 bit_53_99 bitb_53_99 word53_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X54_99 q_54_99 qb_54_99 bit_54_99 bitb_54_99 word54_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X55_99 q_55_99 qb_55_99 bit_55_99 bitb_55_99 word55_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X56_99 q_56_99 qb_56_99 bit_56_99 bitb_56_99 word56_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X57_99 q_57_99 qb_57_99 bit_57_99 bitb_57_99 word57_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X58_99 q_58_99 qb_58_99 bit_58_99 bitb_58_99 word58_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X59_99 q_59_99 qb_59_99 bit_59_99 bitb_59_99 word59_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X60_99 q_60_99 qb_60_99 bit_60_99 bitb_60_99 word60_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X61_99 q_61_99 qb_61_99 bit_61_99 bitb_61_99 word61_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X62_99 q_62_99 qb_62_99 bit_62_99 bitb_62_99 word62_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X63_99 q_63_99 qb_63_99 bit_63_99 bitb_63_99 word63_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X64_99 q_64_99 qb_64_99 bit_64_99 bitb_64_99 word64_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X65_99 q_65_99 qb_65_99 bit_65_99 bitb_65_99 word65_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X66_99 q_66_99 qb_66_99 bit_66_99 bitb_66_99 word66_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X67_99 q_67_99 qb_67_99 bit_67_99 bitb_67_99 word67_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X68_99 q_68_99 qb_68_99 bit_68_99 bitb_68_99 word68_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X69_99 q_69_99 qb_69_99 bit_69_99 bitb_69_99 word69_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X70_99 q_70_99 qb_70_99 bit_70_99 bitb_70_99 word70_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X71_99 q_71_99 qb_71_99 bit_71_99 bitb_71_99 word71_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X72_99 q_72_99 qb_72_99 bit_72_99 bitb_72_99 word72_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X73_99 q_73_99 qb_73_99 bit_73_99 bitb_73_99 word73_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X74_99 q_74_99 qb_74_99 bit_74_99 bitb_74_99 word74_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X75_99 q_75_99 qb_75_99 bit_75_99 bitb_75_99 word75_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X76_99 q_76_99 qb_76_99 bit_76_99 bitb_76_99 word76_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X77_99 q_77_99 qb_77_99 bit_77_99 bitb_77_99 word77_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X78_99 q_78_99 qb_78_99 bit_78_99 bitb_78_99 word78_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X79_99 q_79_99 qb_79_99 bit_79_99 bitb_79_99 word79_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X80_99 q_80_99 qb_80_99 bit_80_99 bitb_80_99 word80_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X81_99 q_81_99 qb_81_99 bit_81_99 bitb_81_99 word81_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X82_99 q_82_99 qb_82_99 bit_82_99 bitb_82_99 word82_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X83_99 q_83_99 qb_83_99 bit_83_99 bitb_83_99 word83_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X84_99 q_84_99 qb_84_99 bit_84_99 bitb_84_99 word84_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X85_99 q_85_99 qb_85_99 bit_85_99 bitb_85_99 word85_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X86_99 q_86_99 qb_86_99 bit_86_99 bitb_86_99 word86_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X87_99 q_87_99 qb_87_99 bit_87_99 bitb_87_99 word87_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X88_99 q_88_99 qb_88_99 bit_88_99 bitb_88_99 word88_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X89_99 q_89_99 qb_89_99 bit_89_99 bitb_89_99 word89_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X90_99 q_90_99 qb_90_99 bit_90_99 bitb_90_99 word90_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X91_99 q_91_99 qb_91_99 bit_91_99 bitb_91_99 word91_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X92_99 q_92_99 qb_92_99 bit_92_99 bitb_92_99 word92_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X93_99 q_93_99 qb_93_99 bit_93_99 bitb_93_99 word93_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X94_99 q_94_99 qb_94_99 bit_94_99 bitb_94_99 word94_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X95_99 q_95_99 qb_95_99 bit_95_99 bitb_95_99 word95_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X96_99 q_96_99 qb_96_99 bit_96_99 bitb_96_99 word96_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X97_99 q_97_99 qb_97_99 bit_97_99 bitb_97_99 word97_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X98_99 q_98_99 qb_98_99 bit_98_99 bitb_98_99 word98_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
X99_99 q_99_99 qb_99_99 bit_99_99 bitb_99_99 word99_99 vdd gnd SRAM_cell W1=W1 L1=2 W3=4 L3=2 W5=W5 L5=2 
Xt0 bit_0_100 bitb_0_100 pc_0 vdd gnd column_pull_up 
Xbr0 bit_0_0 bitb_0_0 col_read_0 sa_vcs sa_out_0 vdd gnd read_driver 
Xbw0 bit_0_0 bitb_0_0 col_write_0 write_0 data_0 datab_0 vdd gnd write_driver
Xt1 bit_1_100 bitb_1_100 pc_1 vdd gnd column_pull_up 
Xbr1 bit_1_0 bitb_1_0 col_read_1 sa_vcs sa_out_1 vdd gnd read_driver 
Xbw1 bit_1_0 bitb_1_0 col_write_1 write_1 data_1 datab_1 vdd gnd write_driver
Xt2 bit_2_100 bitb_2_100 pc_2 vdd gnd column_pull_up 
Xbr2 bit_2_0 bitb_2_0 col_read_2 sa_vcs sa_out_2 vdd gnd read_driver 
Xbw2 bit_2_0 bitb_2_0 col_write_2 write_2 data_2 datab_2 vdd gnd write_driver
Xt3 bit_3_100 bitb_3_100 pc_3 vdd gnd column_pull_up 
Xbr3 bit_3_0 bitb_3_0 col_read_3 sa_vcs sa_out_3 vdd gnd read_driver 
Xbw3 bit_3_0 bitb_3_0 col_write_3 write_3 data_3 datab_3 vdd gnd write_driver
Xt4 bit_4_100 bitb_4_100 pc_4 vdd gnd column_pull_up 
Xbr4 bit_4_0 bitb_4_0 col_read_4 sa_vcs sa_out_4 vdd gnd read_driver 
Xbw4 bit_4_0 bitb_4_0 col_write_4 write_4 data_4 datab_4 vdd gnd write_driver
Xt5 bit_5_100 bitb_5_100 pc_5 vdd gnd column_pull_up 
Xbr5 bit_5_0 bitb_5_0 col_read_5 sa_vcs sa_out_5 vdd gnd read_driver 
Xbw5 bit_5_0 bitb_5_0 col_write_5 write_5 data_5 datab_5 vdd gnd write_driver
Xt6 bit_6_100 bitb_6_100 pc_6 vdd gnd column_pull_up 
Xbr6 bit_6_0 bitb_6_0 col_read_6 sa_vcs sa_out_6 vdd gnd read_driver 
Xbw6 bit_6_0 bitb_6_0 col_write_6 write_6 data_6 datab_6 vdd gnd write_driver
Xt7 bit_7_100 bitb_7_100 pc_7 vdd gnd column_pull_up 
Xbr7 bit_7_0 bitb_7_0 col_read_7 sa_vcs sa_out_7 vdd gnd read_driver 
Xbw7 bit_7_0 bitb_7_0 col_write_7 write_7 data_7 datab_7 vdd gnd write_driver
Xt8 bit_8_100 bitb_8_100 pc_8 vdd gnd column_pull_up 
Xbr8 bit_8_0 bitb_8_0 col_read_8 sa_vcs sa_out_8 vdd gnd read_driver 
Xbw8 bit_8_0 bitb_8_0 col_write_8 write_8 data_8 datab_8 vdd gnd write_driver
Xt9 bit_9_100 bitb_9_100 pc_9 vdd gnd column_pull_up 
Xbr9 bit_9_0 bitb_9_0 col_read_9 sa_vcs sa_out_9 vdd gnd read_driver 
Xbw9 bit_9_0 bitb_9_0 col_write_9 write_9 data_9 datab_9 vdd gnd write_driver
Xt10 bit_10_100 bitb_10_100 pc_10 vdd gnd column_pull_up 
Xbr10 bit_10_0 bitb_10_0 col_read_10 sa_vcs sa_out_10 vdd gnd read_driver 
Xbw10 bit_10_0 bitb_10_0 col_write_10 write_10 data_10 datab_10 vdd gnd write_driver
Xt11 bit_11_100 bitb_11_100 pc_11 vdd gnd column_pull_up 
Xbr11 bit_11_0 bitb_11_0 col_read_11 sa_vcs sa_out_11 vdd gnd read_driver 
Xbw11 bit_11_0 bitb_11_0 col_write_11 write_11 data_11 datab_11 vdd gnd write_driver
Xt12 bit_12_100 bitb_12_100 pc_12 vdd gnd column_pull_up 
Xbr12 bit_12_0 bitb_12_0 col_read_12 sa_vcs sa_out_12 vdd gnd read_driver 
Xbw12 bit_12_0 bitb_12_0 col_write_12 write_12 data_12 datab_12 vdd gnd write_driver
Xt13 bit_13_100 bitb_13_100 pc_13 vdd gnd column_pull_up 
Xbr13 bit_13_0 bitb_13_0 col_read_13 sa_vcs sa_out_13 vdd gnd read_driver 
Xbw13 bit_13_0 bitb_13_0 col_write_13 write_13 data_13 datab_13 vdd gnd write_driver
Xt14 bit_14_100 bitb_14_100 pc_14 vdd gnd column_pull_up 
Xbr14 bit_14_0 bitb_14_0 col_read_14 sa_vcs sa_out_14 vdd gnd read_driver 
Xbw14 bit_14_0 bitb_14_0 col_write_14 write_14 data_14 datab_14 vdd gnd write_driver
Xt15 bit_15_100 bitb_15_100 pc_15 vdd gnd column_pull_up 
Xbr15 bit_15_0 bitb_15_0 col_read_15 sa_vcs sa_out_15 vdd gnd read_driver 
Xbw15 bit_15_0 bitb_15_0 col_write_15 write_15 data_15 datab_15 vdd gnd write_driver
Xt16 bit_16_100 bitb_16_100 pc_16 vdd gnd column_pull_up 
Xbr16 bit_16_0 bitb_16_0 col_read_16 sa_vcs sa_out_16 vdd gnd read_driver 
Xbw16 bit_16_0 bitb_16_0 col_write_16 write_16 data_16 datab_16 vdd gnd write_driver
Xt17 bit_17_100 bitb_17_100 pc_17 vdd gnd column_pull_up 
Xbr17 bit_17_0 bitb_17_0 col_read_17 sa_vcs sa_out_17 vdd gnd read_driver 
Xbw17 bit_17_0 bitb_17_0 col_write_17 write_17 data_17 datab_17 vdd gnd write_driver
Xt18 bit_18_100 bitb_18_100 pc_18 vdd gnd column_pull_up 
Xbr18 bit_18_0 bitb_18_0 col_read_18 sa_vcs sa_out_18 vdd gnd read_driver 
Xbw18 bit_18_0 bitb_18_0 col_write_18 write_18 data_18 datab_18 vdd gnd write_driver
Xt19 bit_19_100 bitb_19_100 pc_19 vdd gnd column_pull_up 
Xbr19 bit_19_0 bitb_19_0 col_read_19 sa_vcs sa_out_19 vdd gnd read_driver 
Xbw19 bit_19_0 bitb_19_0 col_write_19 write_19 data_19 datab_19 vdd gnd write_driver
Xt20 bit_20_100 bitb_20_100 pc_20 vdd gnd column_pull_up 
Xbr20 bit_20_0 bitb_20_0 col_read_20 sa_vcs sa_out_20 vdd gnd read_driver 
Xbw20 bit_20_0 bitb_20_0 col_write_20 write_20 data_20 datab_20 vdd gnd write_driver
Xt21 bit_21_100 bitb_21_100 pc_21 vdd gnd column_pull_up 
Xbr21 bit_21_0 bitb_21_0 col_read_21 sa_vcs sa_out_21 vdd gnd read_driver 
Xbw21 bit_21_0 bitb_21_0 col_write_21 write_21 data_21 datab_21 vdd gnd write_driver
Xt22 bit_22_100 bitb_22_100 pc_22 vdd gnd column_pull_up 
Xbr22 bit_22_0 bitb_22_0 col_read_22 sa_vcs sa_out_22 vdd gnd read_driver 
Xbw22 bit_22_0 bitb_22_0 col_write_22 write_22 data_22 datab_22 vdd gnd write_driver
Xt23 bit_23_100 bitb_23_100 pc_23 vdd gnd column_pull_up 
Xbr23 bit_23_0 bitb_23_0 col_read_23 sa_vcs sa_out_23 vdd gnd read_driver 
Xbw23 bit_23_0 bitb_23_0 col_write_23 write_23 data_23 datab_23 vdd gnd write_driver
Xt24 bit_24_100 bitb_24_100 pc_24 vdd gnd column_pull_up 
Xbr24 bit_24_0 bitb_24_0 col_read_24 sa_vcs sa_out_24 vdd gnd read_driver 
Xbw24 bit_24_0 bitb_24_0 col_write_24 write_24 data_24 datab_24 vdd gnd write_driver
Xt25 bit_25_100 bitb_25_100 pc_25 vdd gnd column_pull_up 
Xbr25 bit_25_0 bitb_25_0 col_read_25 sa_vcs sa_out_25 vdd gnd read_driver 
Xbw25 bit_25_0 bitb_25_0 col_write_25 write_25 data_25 datab_25 vdd gnd write_driver
Xt26 bit_26_100 bitb_26_100 pc_26 vdd gnd column_pull_up 
Xbr26 bit_26_0 bitb_26_0 col_read_26 sa_vcs sa_out_26 vdd gnd read_driver 
Xbw26 bit_26_0 bitb_26_0 col_write_26 write_26 data_26 datab_26 vdd gnd write_driver
Xt27 bit_27_100 bitb_27_100 pc_27 vdd gnd column_pull_up 
Xbr27 bit_27_0 bitb_27_0 col_read_27 sa_vcs sa_out_27 vdd gnd read_driver 
Xbw27 bit_27_0 bitb_27_0 col_write_27 write_27 data_27 datab_27 vdd gnd write_driver
Xt28 bit_28_100 bitb_28_100 pc_28 vdd gnd column_pull_up 
Xbr28 bit_28_0 bitb_28_0 col_read_28 sa_vcs sa_out_28 vdd gnd read_driver 
Xbw28 bit_28_0 bitb_28_0 col_write_28 write_28 data_28 datab_28 vdd gnd write_driver
Xt29 bit_29_100 bitb_29_100 pc_29 vdd gnd column_pull_up 
Xbr29 bit_29_0 bitb_29_0 col_read_29 sa_vcs sa_out_29 vdd gnd read_driver 
Xbw29 bit_29_0 bitb_29_0 col_write_29 write_29 data_29 datab_29 vdd gnd write_driver
Xt30 bit_30_100 bitb_30_100 pc_30 vdd gnd column_pull_up 
Xbr30 bit_30_0 bitb_30_0 col_read_30 sa_vcs sa_out_30 vdd gnd read_driver 
Xbw30 bit_30_0 bitb_30_0 col_write_30 write_30 data_30 datab_30 vdd gnd write_driver
Xt31 bit_31_100 bitb_31_100 pc_31 vdd gnd column_pull_up 
Xbr31 bit_31_0 bitb_31_0 col_read_31 sa_vcs sa_out_31 vdd gnd read_driver 
Xbw31 bit_31_0 bitb_31_0 col_write_31 write_31 data_31 datab_31 vdd gnd write_driver
Xt32 bit_32_100 bitb_32_100 pc_32 vdd gnd column_pull_up 
Xbr32 bit_32_0 bitb_32_0 col_read_32 sa_vcs sa_out_32 vdd gnd read_driver 
Xbw32 bit_32_0 bitb_32_0 col_write_32 write_32 data_32 datab_32 vdd gnd write_driver
Xt33 bit_33_100 bitb_33_100 pc_33 vdd gnd column_pull_up 
Xbr33 bit_33_0 bitb_33_0 col_read_33 sa_vcs sa_out_33 vdd gnd read_driver 
Xbw33 bit_33_0 bitb_33_0 col_write_33 write_33 data_33 datab_33 vdd gnd write_driver
Xt34 bit_34_100 bitb_34_100 pc_34 vdd gnd column_pull_up 
Xbr34 bit_34_0 bitb_34_0 col_read_34 sa_vcs sa_out_34 vdd gnd read_driver 
Xbw34 bit_34_0 bitb_34_0 col_write_34 write_34 data_34 datab_34 vdd gnd write_driver
Xt35 bit_35_100 bitb_35_100 pc_35 vdd gnd column_pull_up 
Xbr35 bit_35_0 bitb_35_0 col_read_35 sa_vcs sa_out_35 vdd gnd read_driver 
Xbw35 bit_35_0 bitb_35_0 col_write_35 write_35 data_35 datab_35 vdd gnd write_driver
Xt36 bit_36_100 bitb_36_100 pc_36 vdd gnd column_pull_up 
Xbr36 bit_36_0 bitb_36_0 col_read_36 sa_vcs sa_out_36 vdd gnd read_driver 
Xbw36 bit_36_0 bitb_36_0 col_write_36 write_36 data_36 datab_36 vdd gnd write_driver
Xt37 bit_37_100 bitb_37_100 pc_37 vdd gnd column_pull_up 
Xbr37 bit_37_0 bitb_37_0 col_read_37 sa_vcs sa_out_37 vdd gnd read_driver 
Xbw37 bit_37_0 bitb_37_0 col_write_37 write_37 data_37 datab_37 vdd gnd write_driver
Xt38 bit_38_100 bitb_38_100 pc_38 vdd gnd column_pull_up 
Xbr38 bit_38_0 bitb_38_0 col_read_38 sa_vcs sa_out_38 vdd gnd read_driver 
Xbw38 bit_38_0 bitb_38_0 col_write_38 write_38 data_38 datab_38 vdd gnd write_driver
Xt39 bit_39_100 bitb_39_100 pc_39 vdd gnd column_pull_up 
Xbr39 bit_39_0 bitb_39_0 col_read_39 sa_vcs sa_out_39 vdd gnd read_driver 
Xbw39 bit_39_0 bitb_39_0 col_write_39 write_39 data_39 datab_39 vdd gnd write_driver
Xt40 bit_40_100 bitb_40_100 pc_40 vdd gnd column_pull_up 
Xbr40 bit_40_0 bitb_40_0 col_read_40 sa_vcs sa_out_40 vdd gnd read_driver 
Xbw40 bit_40_0 bitb_40_0 col_write_40 write_40 data_40 datab_40 vdd gnd write_driver
Xt41 bit_41_100 bitb_41_100 pc_41 vdd gnd column_pull_up 
Xbr41 bit_41_0 bitb_41_0 col_read_41 sa_vcs sa_out_41 vdd gnd read_driver 
Xbw41 bit_41_0 bitb_41_0 col_write_41 write_41 data_41 datab_41 vdd gnd write_driver
Xt42 bit_42_100 bitb_42_100 pc_42 vdd gnd column_pull_up 
Xbr42 bit_42_0 bitb_42_0 col_read_42 sa_vcs sa_out_42 vdd gnd read_driver 
Xbw42 bit_42_0 bitb_42_0 col_write_42 write_42 data_42 datab_42 vdd gnd write_driver
Xt43 bit_43_100 bitb_43_100 pc_43 vdd gnd column_pull_up 
Xbr43 bit_43_0 bitb_43_0 col_read_43 sa_vcs sa_out_43 vdd gnd read_driver 
Xbw43 bit_43_0 bitb_43_0 col_write_43 write_43 data_43 datab_43 vdd gnd write_driver
Xt44 bit_44_100 bitb_44_100 pc_44 vdd gnd column_pull_up 
Xbr44 bit_44_0 bitb_44_0 col_read_44 sa_vcs sa_out_44 vdd gnd read_driver 
Xbw44 bit_44_0 bitb_44_0 col_write_44 write_44 data_44 datab_44 vdd gnd write_driver
Xt45 bit_45_100 bitb_45_100 pc_45 vdd gnd column_pull_up 
Xbr45 bit_45_0 bitb_45_0 col_read_45 sa_vcs sa_out_45 vdd gnd read_driver 
Xbw45 bit_45_0 bitb_45_0 col_write_45 write_45 data_45 datab_45 vdd gnd write_driver
Xt46 bit_46_100 bitb_46_100 pc_46 vdd gnd column_pull_up 
Xbr46 bit_46_0 bitb_46_0 col_read_46 sa_vcs sa_out_46 vdd gnd read_driver 
Xbw46 bit_46_0 bitb_46_0 col_write_46 write_46 data_46 datab_46 vdd gnd write_driver
Xt47 bit_47_100 bitb_47_100 pc_47 vdd gnd column_pull_up 
Xbr47 bit_47_0 bitb_47_0 col_read_47 sa_vcs sa_out_47 vdd gnd read_driver 
Xbw47 bit_47_0 bitb_47_0 col_write_47 write_47 data_47 datab_47 vdd gnd write_driver
Xt48 bit_48_100 bitb_48_100 pc_48 vdd gnd column_pull_up 
Xbr48 bit_48_0 bitb_48_0 col_read_48 sa_vcs sa_out_48 vdd gnd read_driver 
Xbw48 bit_48_0 bitb_48_0 col_write_48 write_48 data_48 datab_48 vdd gnd write_driver
Xt49 bit_49_100 bitb_49_100 pc_49 vdd gnd column_pull_up 
Xbr49 bit_49_0 bitb_49_0 col_read_49 sa_vcs sa_out_49 vdd gnd read_driver 
Xbw49 bit_49_0 bitb_49_0 col_write_49 write_49 data_49 datab_49 vdd gnd write_driver
Xt50 bit_50_100 bitb_50_100 pc_50 vdd gnd column_pull_up 
Xbr50 bit_50_0 bitb_50_0 col_read_50 sa_vcs sa_out_50 vdd gnd read_driver 
Xbw50 bit_50_0 bitb_50_0 col_write_50 write_50 data_50 datab_50 vdd gnd write_driver
Xt51 bit_51_100 bitb_51_100 pc_51 vdd gnd column_pull_up 
Xbr51 bit_51_0 bitb_51_0 col_read_51 sa_vcs sa_out_51 vdd gnd read_driver 
Xbw51 bit_51_0 bitb_51_0 col_write_51 write_51 data_51 datab_51 vdd gnd write_driver
Xt52 bit_52_100 bitb_52_100 pc_52 vdd gnd column_pull_up 
Xbr52 bit_52_0 bitb_52_0 col_read_52 sa_vcs sa_out_52 vdd gnd read_driver 
Xbw52 bit_52_0 bitb_52_0 col_write_52 write_52 data_52 datab_52 vdd gnd write_driver
Xt53 bit_53_100 bitb_53_100 pc_53 vdd gnd column_pull_up 
Xbr53 bit_53_0 bitb_53_0 col_read_53 sa_vcs sa_out_53 vdd gnd read_driver 
Xbw53 bit_53_0 bitb_53_0 col_write_53 write_53 data_53 datab_53 vdd gnd write_driver
Xt54 bit_54_100 bitb_54_100 pc_54 vdd gnd column_pull_up 
Xbr54 bit_54_0 bitb_54_0 col_read_54 sa_vcs sa_out_54 vdd gnd read_driver 
Xbw54 bit_54_0 bitb_54_0 col_write_54 write_54 data_54 datab_54 vdd gnd write_driver
Xt55 bit_55_100 bitb_55_100 pc_55 vdd gnd column_pull_up 
Xbr55 bit_55_0 bitb_55_0 col_read_55 sa_vcs sa_out_55 vdd gnd read_driver 
Xbw55 bit_55_0 bitb_55_0 col_write_55 write_55 data_55 datab_55 vdd gnd write_driver
Xt56 bit_56_100 bitb_56_100 pc_56 vdd gnd column_pull_up 
Xbr56 bit_56_0 bitb_56_0 col_read_56 sa_vcs sa_out_56 vdd gnd read_driver 
Xbw56 bit_56_0 bitb_56_0 col_write_56 write_56 data_56 datab_56 vdd gnd write_driver
Xt57 bit_57_100 bitb_57_100 pc_57 vdd gnd column_pull_up 
Xbr57 bit_57_0 bitb_57_0 col_read_57 sa_vcs sa_out_57 vdd gnd read_driver 
Xbw57 bit_57_0 bitb_57_0 col_write_57 write_57 data_57 datab_57 vdd gnd write_driver
Xt58 bit_58_100 bitb_58_100 pc_58 vdd gnd column_pull_up 
Xbr58 bit_58_0 bitb_58_0 col_read_58 sa_vcs sa_out_58 vdd gnd read_driver 
Xbw58 bit_58_0 bitb_58_0 col_write_58 write_58 data_58 datab_58 vdd gnd write_driver
Xt59 bit_59_100 bitb_59_100 pc_59 vdd gnd column_pull_up 
Xbr59 bit_59_0 bitb_59_0 col_read_59 sa_vcs sa_out_59 vdd gnd read_driver 
Xbw59 bit_59_0 bitb_59_0 col_write_59 write_59 data_59 datab_59 vdd gnd write_driver
Xt60 bit_60_100 bitb_60_100 pc_60 vdd gnd column_pull_up 
Xbr60 bit_60_0 bitb_60_0 col_read_60 sa_vcs sa_out_60 vdd gnd read_driver 
Xbw60 bit_60_0 bitb_60_0 col_write_60 write_60 data_60 datab_60 vdd gnd write_driver
Xt61 bit_61_100 bitb_61_100 pc_61 vdd gnd column_pull_up 
Xbr61 bit_61_0 bitb_61_0 col_read_61 sa_vcs sa_out_61 vdd gnd read_driver 
Xbw61 bit_61_0 bitb_61_0 col_write_61 write_61 data_61 datab_61 vdd gnd write_driver
Xt62 bit_62_100 bitb_62_100 pc_62 vdd gnd column_pull_up 
Xbr62 bit_62_0 bitb_62_0 col_read_62 sa_vcs sa_out_62 vdd gnd read_driver 
Xbw62 bit_62_0 bitb_62_0 col_write_62 write_62 data_62 datab_62 vdd gnd write_driver
Xt63 bit_63_100 bitb_63_100 pc_63 vdd gnd column_pull_up 
Xbr63 bit_63_0 bitb_63_0 col_read_63 sa_vcs sa_out_63 vdd gnd read_driver 
Xbw63 bit_63_0 bitb_63_0 col_write_63 write_63 data_63 datab_63 vdd gnd write_driver
Xt64 bit_64_100 bitb_64_100 pc_64 vdd gnd column_pull_up 
Xbr64 bit_64_0 bitb_64_0 col_read_64 sa_vcs sa_out_64 vdd gnd read_driver 
Xbw64 bit_64_0 bitb_64_0 col_write_64 write_64 data_64 datab_64 vdd gnd write_driver
Xt65 bit_65_100 bitb_65_100 pc_65 vdd gnd column_pull_up 
Xbr65 bit_65_0 bitb_65_0 col_read_65 sa_vcs sa_out_65 vdd gnd read_driver 
Xbw65 bit_65_0 bitb_65_0 col_write_65 write_65 data_65 datab_65 vdd gnd write_driver
Xt66 bit_66_100 bitb_66_100 pc_66 vdd gnd column_pull_up 
Xbr66 bit_66_0 bitb_66_0 col_read_66 sa_vcs sa_out_66 vdd gnd read_driver 
Xbw66 bit_66_0 bitb_66_0 col_write_66 write_66 data_66 datab_66 vdd gnd write_driver
Xt67 bit_67_100 bitb_67_100 pc_67 vdd gnd column_pull_up 
Xbr67 bit_67_0 bitb_67_0 col_read_67 sa_vcs sa_out_67 vdd gnd read_driver 
Xbw67 bit_67_0 bitb_67_0 col_write_67 write_67 data_67 datab_67 vdd gnd write_driver
Xt68 bit_68_100 bitb_68_100 pc_68 vdd gnd column_pull_up 
Xbr68 bit_68_0 bitb_68_0 col_read_68 sa_vcs sa_out_68 vdd gnd read_driver 
Xbw68 bit_68_0 bitb_68_0 col_write_68 write_68 data_68 datab_68 vdd gnd write_driver
Xt69 bit_69_100 bitb_69_100 pc_69 vdd gnd column_pull_up 
Xbr69 bit_69_0 bitb_69_0 col_read_69 sa_vcs sa_out_69 vdd gnd read_driver 
Xbw69 bit_69_0 bitb_69_0 col_write_69 write_69 data_69 datab_69 vdd gnd write_driver
Xt70 bit_70_100 bitb_70_100 pc_70 vdd gnd column_pull_up 
Xbr70 bit_70_0 bitb_70_0 col_read_70 sa_vcs sa_out_70 vdd gnd read_driver 
Xbw70 bit_70_0 bitb_70_0 col_write_70 write_70 data_70 datab_70 vdd gnd write_driver
Xt71 bit_71_100 bitb_71_100 pc_71 vdd gnd column_pull_up 
Xbr71 bit_71_0 bitb_71_0 col_read_71 sa_vcs sa_out_71 vdd gnd read_driver 
Xbw71 bit_71_0 bitb_71_0 col_write_71 write_71 data_71 datab_71 vdd gnd write_driver
Xt72 bit_72_100 bitb_72_100 pc_72 vdd gnd column_pull_up 
Xbr72 bit_72_0 bitb_72_0 col_read_72 sa_vcs sa_out_72 vdd gnd read_driver 
Xbw72 bit_72_0 bitb_72_0 col_write_72 write_72 data_72 datab_72 vdd gnd write_driver
Xt73 bit_73_100 bitb_73_100 pc_73 vdd gnd column_pull_up 
Xbr73 bit_73_0 bitb_73_0 col_read_73 sa_vcs sa_out_73 vdd gnd read_driver 
Xbw73 bit_73_0 bitb_73_0 col_write_73 write_73 data_73 datab_73 vdd gnd write_driver
Xt74 bit_74_100 bitb_74_100 pc_74 vdd gnd column_pull_up 
Xbr74 bit_74_0 bitb_74_0 col_read_74 sa_vcs sa_out_74 vdd gnd read_driver 
Xbw74 bit_74_0 bitb_74_0 col_write_74 write_74 data_74 datab_74 vdd gnd write_driver
Xt75 bit_75_100 bitb_75_100 pc_75 vdd gnd column_pull_up 
Xbr75 bit_75_0 bitb_75_0 col_read_75 sa_vcs sa_out_75 vdd gnd read_driver 
Xbw75 bit_75_0 bitb_75_0 col_write_75 write_75 data_75 datab_75 vdd gnd write_driver
Xt76 bit_76_100 bitb_76_100 pc_76 vdd gnd column_pull_up 
Xbr76 bit_76_0 bitb_76_0 col_read_76 sa_vcs sa_out_76 vdd gnd read_driver 
Xbw76 bit_76_0 bitb_76_0 col_write_76 write_76 data_76 datab_76 vdd gnd write_driver
Xt77 bit_77_100 bitb_77_100 pc_77 vdd gnd column_pull_up 
Xbr77 bit_77_0 bitb_77_0 col_read_77 sa_vcs sa_out_77 vdd gnd read_driver 
Xbw77 bit_77_0 bitb_77_0 col_write_77 write_77 data_77 datab_77 vdd gnd write_driver
Xt78 bit_78_100 bitb_78_100 pc_78 vdd gnd column_pull_up 
Xbr78 bit_78_0 bitb_78_0 col_read_78 sa_vcs sa_out_78 vdd gnd read_driver 
Xbw78 bit_78_0 bitb_78_0 col_write_78 write_78 data_78 datab_78 vdd gnd write_driver
Xt79 bit_79_100 bitb_79_100 pc_79 vdd gnd column_pull_up 
Xbr79 bit_79_0 bitb_79_0 col_read_79 sa_vcs sa_out_79 vdd gnd read_driver 
Xbw79 bit_79_0 bitb_79_0 col_write_79 write_79 data_79 datab_79 vdd gnd write_driver
Xt80 bit_80_100 bitb_80_100 pc_80 vdd gnd column_pull_up 
Xbr80 bit_80_0 bitb_80_0 col_read_80 sa_vcs sa_out_80 vdd gnd read_driver 
Xbw80 bit_80_0 bitb_80_0 col_write_80 write_80 data_80 datab_80 vdd gnd write_driver
Xt81 bit_81_100 bitb_81_100 pc_81 vdd gnd column_pull_up 
Xbr81 bit_81_0 bitb_81_0 col_read_81 sa_vcs sa_out_81 vdd gnd read_driver 
Xbw81 bit_81_0 bitb_81_0 col_write_81 write_81 data_81 datab_81 vdd gnd write_driver
Xt82 bit_82_100 bitb_82_100 pc_82 vdd gnd column_pull_up 
Xbr82 bit_82_0 bitb_82_0 col_read_82 sa_vcs sa_out_82 vdd gnd read_driver 
Xbw82 bit_82_0 bitb_82_0 col_write_82 write_82 data_82 datab_82 vdd gnd write_driver
Xt83 bit_83_100 bitb_83_100 pc_83 vdd gnd column_pull_up 
Xbr83 bit_83_0 bitb_83_0 col_read_83 sa_vcs sa_out_83 vdd gnd read_driver 
Xbw83 bit_83_0 bitb_83_0 col_write_83 write_83 data_83 datab_83 vdd gnd write_driver
Xt84 bit_84_100 bitb_84_100 pc_84 vdd gnd column_pull_up 
Xbr84 bit_84_0 bitb_84_0 col_read_84 sa_vcs sa_out_84 vdd gnd read_driver 
Xbw84 bit_84_0 bitb_84_0 col_write_84 write_84 data_84 datab_84 vdd gnd write_driver
Xt85 bit_85_100 bitb_85_100 pc_85 vdd gnd column_pull_up 
Xbr85 bit_85_0 bitb_85_0 col_read_85 sa_vcs sa_out_85 vdd gnd read_driver 
Xbw85 bit_85_0 bitb_85_0 col_write_85 write_85 data_85 datab_85 vdd gnd write_driver
Xt86 bit_86_100 bitb_86_100 pc_86 vdd gnd column_pull_up 
Xbr86 bit_86_0 bitb_86_0 col_read_86 sa_vcs sa_out_86 vdd gnd read_driver 
Xbw86 bit_86_0 bitb_86_0 col_write_86 write_86 data_86 datab_86 vdd gnd write_driver
Xt87 bit_87_100 bitb_87_100 pc_87 vdd gnd column_pull_up 
Xbr87 bit_87_0 bitb_87_0 col_read_87 sa_vcs sa_out_87 vdd gnd read_driver 
Xbw87 bit_87_0 bitb_87_0 col_write_87 write_87 data_87 datab_87 vdd gnd write_driver
Xt88 bit_88_100 bitb_88_100 pc_88 vdd gnd column_pull_up 
Xbr88 bit_88_0 bitb_88_0 col_read_88 sa_vcs sa_out_88 vdd gnd read_driver 
Xbw88 bit_88_0 bitb_88_0 col_write_88 write_88 data_88 datab_88 vdd gnd write_driver
Xt89 bit_89_100 bitb_89_100 pc_89 vdd gnd column_pull_up 
Xbr89 bit_89_0 bitb_89_0 col_read_89 sa_vcs sa_out_89 vdd gnd read_driver 
Xbw89 bit_89_0 bitb_89_0 col_write_89 write_89 data_89 datab_89 vdd gnd write_driver
Xt90 bit_90_100 bitb_90_100 pc_90 vdd gnd column_pull_up 
Xbr90 bit_90_0 bitb_90_0 col_read_90 sa_vcs sa_out_90 vdd gnd read_driver 
Xbw90 bit_90_0 bitb_90_0 col_write_90 write_90 data_90 datab_90 vdd gnd write_driver
Xt91 bit_91_100 bitb_91_100 pc_91 vdd gnd column_pull_up 
Xbr91 bit_91_0 bitb_91_0 col_read_91 sa_vcs sa_out_91 vdd gnd read_driver 
Xbw91 bit_91_0 bitb_91_0 col_write_91 write_91 data_91 datab_91 vdd gnd write_driver
Xt92 bit_92_100 bitb_92_100 pc_92 vdd gnd column_pull_up 
Xbr92 bit_92_0 bitb_92_0 col_read_92 sa_vcs sa_out_92 vdd gnd read_driver 
Xbw92 bit_92_0 bitb_92_0 col_write_92 write_92 data_92 datab_92 vdd gnd write_driver
Xt93 bit_93_100 bitb_93_100 pc_93 vdd gnd column_pull_up 
Xbr93 bit_93_0 bitb_93_0 col_read_93 sa_vcs sa_out_93 vdd gnd read_driver 
Xbw93 bit_93_0 bitb_93_0 col_write_93 write_93 data_93 datab_93 vdd gnd write_driver
Xt94 bit_94_100 bitb_94_100 pc_94 vdd gnd column_pull_up 
Xbr94 bit_94_0 bitb_94_0 col_read_94 sa_vcs sa_out_94 vdd gnd read_driver 
Xbw94 bit_94_0 bitb_94_0 col_write_94 write_94 data_94 datab_94 vdd gnd write_driver
Xt95 bit_95_100 bitb_95_100 pc_95 vdd gnd column_pull_up 
Xbr95 bit_95_0 bitb_95_0 col_read_95 sa_vcs sa_out_95 vdd gnd read_driver 
Xbw95 bit_95_0 bitb_95_0 col_write_95 write_95 data_95 datab_95 vdd gnd write_driver
Xt96 bit_96_100 bitb_96_100 pc_96 vdd gnd column_pull_up 
Xbr96 bit_96_0 bitb_96_0 col_read_96 sa_vcs sa_out_96 vdd gnd read_driver 
Xbw96 bit_96_0 bitb_96_0 col_write_96 write_96 data_96 datab_96 vdd gnd write_driver
Xt97 bit_97_100 bitb_97_100 pc_97 vdd gnd column_pull_up 
Xbr97 bit_97_0 bitb_97_0 col_read_97 sa_vcs sa_out_97 vdd gnd read_driver 
Xbw97 bit_97_0 bitb_97_0 col_write_97 write_97 data_97 datab_97 vdd gnd write_driver
Xt98 bit_98_100 bitb_98_100 pc_98 vdd gnd column_pull_up 
Xbr98 bit_98_0 bitb_98_0 col_read_98 sa_vcs sa_out_98 vdd gnd read_driver 
Xbw98 bit_98_0 bitb_98_0 col_write_98 write_98 data_98 datab_98 vdd gnd write_driver
Xt99 bit_99_100 bitb_99_100 pc_99 vdd gnd column_pull_up 
Xbr99 bit_99_0 bitb_99_0 col_read_99 sa_vcs sa_out_99 vdd gnd read_driver 
Xbw99 bit_99_0 bitb_99_0 col_write_99 write_99 data_99 datab_99 vdd gnd write_driver
.options post probe
.tran 1n 70n uic
.probe I(X5_5.M3) I(X5_5.M4) V(bit_99_0) V(bitb_99_0) V(word_99) V(q_99_99) V(qb_99_99) V(sa_out_99) V(pc_99) V(col_read_99) V(col_write_99) V(write_99) V(data_99) V(datab_99)
.end
